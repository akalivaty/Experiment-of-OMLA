//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n202), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT64), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n235), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G13), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n249), .A2(new_n209), .A3(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n217), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n208), .A2(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n249), .A2(G1), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n254), .A2(new_n258), .B1(new_n260), .B2(new_n256), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G1), .A3(G13), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n266), .A2(new_n232), .B1(new_n267), .B2(new_n265), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n264), .B(KEYINPUT66), .ZN(new_n269));
  OR2_X1    g0069(.A1(G223), .A2(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(G226), .B2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  OAI22_X1  g0076(.A1(new_n272), .A2(new_n275), .B1(new_n276), .B2(new_n222), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n268), .B1(new_n269), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G200), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(G190), .B2(new_n278), .ZN(new_n281));
  INV_X1    g0081(.A(new_n252), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n276), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n209), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT7), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT7), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n284), .A2(new_n288), .A3(new_n209), .A4(new_n285), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(G68), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(G58), .B(G68), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n291), .A2(G20), .B1(G159), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT16), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n282), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT77), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n290), .A2(KEYINPUT16), .A3(new_n293), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n262), .B(new_n281), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT17), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n294), .A2(new_n295), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(new_n252), .A3(new_n298), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT77), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n308), .A2(KEYINPUT17), .A3(new_n262), .A4(new_n281), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n262), .B1(new_n299), .B2(new_n300), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT79), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n278), .A2(G169), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT78), .ZN(new_n314));
  INV_X1    g0114(.A(G179), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(new_n278), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n278), .A2(new_n314), .A3(new_n315), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT18), .A4(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT18), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n261), .B1(new_n306), .B2(new_n307), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n318), .B1(new_n313), .B2(new_n316), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n324), .B1(new_n308), .B2(new_n262), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n312), .B1(new_n327), .B2(KEYINPUT18), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n310), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n265), .A2(new_n267), .ZN(new_n330));
  INV_X1    g0130(.A(new_n266), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(G238), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT66), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n264), .B(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(G232), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT72), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n284), .A2(new_n285), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT72), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(G232), .A4(G1698), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(G226), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G97), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n334), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT73), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n332), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n343), .B1(new_n339), .B2(new_n336), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n348), .A2(KEYINPUT73), .A3(new_n334), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT13), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n345), .A2(new_n346), .ZN(new_n351));
  OAI21_X1  g0151(.A(KEYINPUT73), .B1(new_n348), .B2(new_n334), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT13), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .A4(new_n332), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n350), .A2(G190), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT75), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT74), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n350), .A2(new_n357), .A3(new_n354), .ZN(new_n358));
  OAI211_X1 g0158(.A(KEYINPUT74), .B(KEYINPUT13), .C1(new_n347), .C2(new_n349), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(G200), .A3(new_n359), .ZN(new_n360));
  AOI211_X1 g0160(.A(G68), .B(new_n260), .C1(KEYINPUT76), .C2(KEYINPUT12), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT76), .A2(KEYINPUT12), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n361), .B(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n253), .A2(G68), .A3(new_n257), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n292), .ZN(new_n366));
  INV_X1    g0166(.A(G50), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n366), .A2(new_n367), .B1(new_n209), .B2(G68), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n209), .A2(G33), .ZN(new_n369));
  INV_X1    g0169(.A(G77), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n252), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  XOR2_X1   g0172(.A(new_n372), .B(KEYINPUT11), .Z(new_n373));
  NOR2_X1   g0173(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n360), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n356), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n271), .B1(new_n284), .B2(new_n285), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(G223), .B1(new_n275), .B2(G77), .ZN(new_n378));
  INV_X1    g0178(.A(G222), .ZN(new_n379));
  AOI21_X1  g0179(.A(G1698), .B1(new_n284), .B2(new_n285), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n378), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n269), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n330), .B1(new_n331), .B2(G226), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G190), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n279), .B1(new_n383), .B2(new_n384), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n391));
  INV_X1    g0191(.A(G150), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(new_n366), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n255), .A2(new_n369), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n252), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n253), .A2(G50), .A3(new_n257), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n395), .B(new_n396), .C1(G50), .C2(new_n260), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT9), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n398), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT70), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT10), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n401), .A2(KEYINPUT10), .ZN(new_n404));
  OR3_X1    g0204(.A1(new_n390), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n404), .B1(new_n390), .B2(new_n403), .ZN(new_n406));
  INV_X1    g0206(.A(G169), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n385), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n408), .B(new_n397), .C1(G179), .C2(new_n385), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n405), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT68), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n255), .B1(new_n411), .B2(new_n366), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n411), .B2(new_n366), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT15), .B(G87), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n369), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(G20), .B2(G77), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n282), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n253), .A2(G77), .A3(new_n257), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT69), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n250), .B2(new_n370), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n260), .A2(KEYINPUT69), .A3(G77), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n330), .B1(new_n331), .B2(G244), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n337), .A2(G1698), .ZN(new_n425));
  INV_X1    g0225(.A(G107), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n425), .A2(new_n221), .B1(new_n426), .B2(new_n337), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT67), .B1(new_n381), .B2(new_n232), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT67), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n380), .A2(new_n429), .A3(G232), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n427), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n424), .B1(new_n431), .B2(new_n334), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n423), .B1(G200), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n386), .B2(new_n432), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n407), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n315), .B(new_n424), .C1(new_n431), .C2(new_n334), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n423), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT71), .B1(new_n410), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n410), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT71), .ZN(new_n441));
  INV_X1    g0241(.A(new_n438), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI211_X1 g0243(.A(new_n329), .B(new_n376), .C1(new_n439), .C2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n358), .A2(G169), .A3(new_n359), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT14), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT14), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n358), .A2(new_n447), .A3(G169), .A4(new_n359), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n350), .A2(G179), .A3(new_n354), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n374), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n444), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT6), .ZN(new_n455));
  AND2_X1   g0255(.A1(G97), .A2(G107), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n205), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n426), .A2(KEYINPUT6), .A3(G97), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n459), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n287), .A2(G107), .A3(new_n289), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n252), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT80), .B1(new_n260), .B2(G97), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT80), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n250), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n253), .B1(G1), .B2(new_n276), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n466), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT83), .B1(new_n463), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n282), .B1(new_n460), .B2(new_n461), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT83), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n473), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n380), .A2(KEYINPUT4), .A3(G244), .ZN(new_n476));
  OAI211_X1 g0276(.A(G244), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT4), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n377), .A2(G250), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n476), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n269), .ZN(new_n483));
  INV_X1    g0283(.A(G41), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n208), .B(G45), .C1(new_n484), .C2(KEYINPUT5), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT81), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n264), .A2(G274), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT82), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT5), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(G41), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n484), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n489), .A2(G41), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n264), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n486), .A2(new_n492), .B1(new_n496), .B2(G257), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n483), .A2(new_n497), .A3(G179), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n407), .B1(new_n483), .B2(new_n497), .ZN(new_n499));
  OAI22_X1  g0299(.A1(new_n472), .A2(new_n475), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(G244), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n501));
  OAI211_X1 g0301(.A(G238), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G116), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT84), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT84), .A4(new_n503), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n334), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G45), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G1), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(G250), .A3(new_n264), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n267), .B2(new_n511), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n315), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n407), .B1(new_n508), .B2(new_n513), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n337), .A2(new_n209), .A3(G68), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n209), .B1(new_n342), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(G87), .B2(new_n206), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n369), .B2(new_n466), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(new_n252), .B1(new_n250), .B2(new_n414), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n414), .B2(new_n469), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n515), .A2(new_n516), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n514), .A2(G190), .ZN(new_n526));
  OAI21_X1  g0326(.A(G200), .B1(new_n508), .B2(new_n513), .ZN(new_n527));
  INV_X1    g0327(.A(new_n469), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G87), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n529), .A2(new_n523), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n483), .A2(new_n497), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G200), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n473), .A2(new_n470), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n534), .C1(new_n386), .C2(new_n532), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n500), .A2(new_n525), .A3(new_n531), .A4(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n492), .A2(new_n486), .ZN(new_n538));
  OAI211_X1 g0338(.A(G264), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n540));
  INV_X1    g0340(.A(G303), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n337), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n269), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n496), .A2(G270), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n538), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n253), .B(G116), .C1(G1), .C2(new_n276), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n250), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(G20), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n252), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n481), .B(new_n209), .C1(G33), .C2(new_n466), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT20), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND4_X1   g0352(.A1(KEYINPUT20), .A2(new_n551), .A3(new_n252), .A4(new_n549), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n546), .B(new_n548), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n545), .A2(new_n554), .A3(G169), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT21), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n545), .A2(new_n554), .A3(KEYINPUT21), .A4(G169), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n538), .A2(new_n544), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n559), .A2(G179), .A3(new_n554), .A4(new_n543), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(G190), .A3(new_n543), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n554), .B1(new_n545), .B2(G200), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT24), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n209), .B(G87), .C1(new_n273), .C2(new_n274), .ZN(new_n566));
  XOR2_X1   g0366(.A(KEYINPUT85), .B(KEYINPUT22), .Z(new_n567));
  OR2_X1    g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT23), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n209), .B2(G107), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n426), .A2(KEYINPUT23), .A3(G20), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(G20), .B2(new_n503), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n565), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  AOI211_X1 g0377(.A(KEYINPUT24), .B(new_n575), .C1(new_n568), .C2(new_n569), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n252), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G250), .B(new_n271), .C1(new_n273), .C2(new_n274), .ZN(new_n580));
  OAI211_X1 g0380(.A(G257), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n581));
  INV_X1    g0381(.A(G294), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n580), .B(new_n581), .C1(new_n276), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n269), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n496), .A2(G264), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(G190), .A3(new_n538), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT25), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n260), .B2(G107), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n250), .A2(KEYINPUT25), .A3(new_n426), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n528), .A2(G107), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n538), .A2(new_n584), .A3(new_n585), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G200), .ZN(new_n593));
  AND4_X1   g0393(.A1(new_n579), .A2(new_n587), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n407), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n538), .A2(new_n584), .A3(new_n315), .A4(new_n585), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n579), .B2(new_n591), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AND4_X1   g0399(.A1(new_n454), .A2(new_n537), .A3(new_n564), .A4(new_n599), .ZN(G372));
  NAND2_X1  g0400(.A1(new_n525), .A2(new_n531), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT26), .B1(new_n601), .B2(new_n500), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n579), .A2(new_n591), .A3(new_n587), .A4(new_n593), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n598), .B2(new_n561), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n602), .B1(new_n536), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n498), .A2(new_n499), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n534), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(new_n525), .A3(new_n531), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n525), .B1(new_n608), .B2(KEYINPUT26), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n454), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g0411(.A(new_n611), .B(KEYINPUT86), .Z(new_n612));
  NAND2_X1  g0412(.A1(new_n303), .A2(new_n309), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n376), .A2(new_n437), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n452), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n311), .A2(KEYINPUT18), .A3(new_n320), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n325), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n406), .B(new_n405), .C1(new_n615), .C2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n409), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n612), .A2(new_n619), .ZN(G369));
  NAND2_X1  g0420(.A1(new_n259), .A2(new_n209), .ZN(new_n621));
  OR2_X1    g0421(.A1(new_n621), .A2(KEYINPUT27), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(KEYINPUT27), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(G213), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(G343), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n554), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n564), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(new_n627), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(G330), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n570), .A2(new_n576), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT24), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n570), .A2(new_n565), .A3(new_n576), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n282), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n591), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n626), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n599), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n595), .B(new_n596), .C1(new_n636), .C2(new_n637), .ZN(new_n640));
  INV_X1    g0440(.A(new_n626), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n632), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n629), .A2(new_n626), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n599), .ZN(new_n646));
  XOR2_X1   g0446(.A(new_n626), .B(KEYINPUT87), .Z(new_n647));
  OAI21_X1  g0447(.A(new_n646), .B1(new_n640), .B2(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n644), .A2(new_n648), .ZN(G399));
  INV_X1    g0449(.A(new_n212), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT88), .B1(new_n650), .B2(G41), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n650), .A2(KEYINPUT88), .A3(G41), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n205), .A2(new_n222), .A3(new_n547), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n654), .A2(new_n208), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n216), .B2(new_n654), .ZN(new_n657));
  XOR2_X1   g0457(.A(new_n657), .B(KEYINPUT28), .Z(new_n658));
  INV_X1    g0458(.A(new_n647), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n610), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT29), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n594), .B1(new_n629), .B2(new_n640), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n537), .A2(KEYINPUT90), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT90), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n604), .B2(new_n536), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  OR3_X1    g0467(.A1(new_n601), .A2(KEYINPUT26), .A3(new_n500), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n608), .A2(KEYINPUT26), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(new_n525), .ZN(new_n670));
  OAI211_X1 g0470(.A(KEYINPUT29), .B(new_n641), .C1(new_n667), .C2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n662), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT31), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n532), .A2(new_n315), .A3(new_n545), .A4(new_n592), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n514), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n559), .A2(KEYINPUT89), .A3(G179), .A4(new_n543), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT89), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n545), .B2(new_n315), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n532), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n514), .A3(new_n586), .ZN(new_n681));
  OR3_X1    g0481(.A1(new_n679), .A2(new_n681), .A3(KEYINPUT30), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT30), .B1(new_n679), .B2(new_n681), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n675), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n673), .B1(new_n684), .B2(new_n641), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n537), .A2(new_n564), .A3(new_n599), .A4(new_n659), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  INV_X1    g0487(.A(new_n675), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT31), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n685), .B(new_n686), .C1(new_n690), .C2(new_n659), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n672), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT91), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT91), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n658), .B1(new_n696), .B2(G1), .ZN(G364));
  XNOR2_X1  g0497(.A(new_n631), .B(KEYINPUT92), .ZN(new_n698));
  INV_X1    g0498(.A(new_n654), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n249), .A2(G20), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n208), .B1(new_n700), .B2(G45), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n698), .B(new_n702), .C1(G330), .C2(new_n630), .ZN(new_n703));
  INV_X1    g0503(.A(new_n702), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n315), .A2(new_n279), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n209), .A2(G190), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n315), .A2(G200), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n706), .ZN(new_n709));
  OAI22_X1  g0509(.A1(new_n707), .A2(new_n202), .B1(new_n709), .B2(new_n370), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n209), .A2(new_n386), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n279), .A2(G179), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n706), .A2(new_n712), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI22_X1  g0516(.A1(G87), .A2(new_n714), .B1(new_n716), .B2(G107), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n711), .A2(new_n705), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n717), .B(new_n337), .C1(new_n367), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n711), .A2(new_n708), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AOI211_X1 g0521(.A(new_n710), .B(new_n719), .C1(G58), .C2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G179), .A2(G200), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n706), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G159), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT32), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n209), .B1(new_n723), .B2(G190), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n466), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G311), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n275), .B1(new_n709), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G322), .ZN(new_n733));
  INV_X1    g0533(.A(G283), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n720), .A2(new_n733), .B1(new_n715), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n728), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n732), .B(new_n735), .C1(G294), .C2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n718), .ZN(new_n738));
  AOI22_X1  g0538(.A1(new_n738), .A2(G326), .B1(new_n725), .B2(G329), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n541), .B2(new_n713), .ZN(new_n740));
  XNOR2_X1  g0540(.A(KEYINPUT33), .B(G317), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT94), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n707), .B1(new_n741), .B2(KEYINPUT94), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n722), .A2(new_n730), .B1(new_n737), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n217), .B1(G20), .B2(new_n407), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n704), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n746), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT93), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n216), .A2(new_n509), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n650), .A2(new_n337), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(new_n244), .C2(new_n509), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n650), .A2(new_n275), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n757), .A2(G355), .B1(new_n547), .B2(new_n650), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n753), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n748), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n751), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n630), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n703), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(G396));
  NAND2_X1  g0564(.A1(new_n423), .A2(new_n626), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n434), .A2(new_n437), .A3(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n435), .A2(new_n436), .A3(new_n423), .A4(new_n626), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT96), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n660), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n766), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n659), .B(new_n771), .C1(new_n605), .C2(new_n609), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n704), .B1(new_n773), .B2(new_n692), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n692), .B2(new_n773), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n707), .A2(new_n734), .B1(new_n709), .B2(new_n547), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT95), .ZN(new_n777));
  AOI22_X1  g0577(.A1(G107), .A2(new_n714), .B1(new_n721), .B2(G294), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G87), .A2(new_n716), .B1(new_n725), .B2(G311), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n337), .B(new_n729), .C1(G303), .C2(new_n738), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n777), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n707), .A2(new_n392), .ZN(new_n782));
  INV_X1    g0582(.A(G143), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n720), .A2(new_n783), .B1(new_n709), .B2(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n782), .B(new_n785), .C1(G137), .C2(new_n738), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n337), .B1(new_n713), .B2(new_n367), .ZN(new_n788));
  INV_X1    g0588(.A(G132), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n715), .A2(new_n202), .B1(new_n724), .B2(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n788), .B(new_n790), .C1(G58), .C2(new_n736), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n781), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n746), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n746), .A2(new_n749), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n702), .B1(new_n370), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n795), .B(new_n797), .C1(new_n771), .C2(new_n750), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n775), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G384));
  NOR2_X1   g0600(.A1(new_n700), .A2(new_n208), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n305), .A2(new_n262), .ZN(new_n802));
  INV_X1    g0602(.A(new_n624), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT100), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n320), .A2(new_n802), .ZN(new_n806));
  AND3_X1   g0606(.A1(new_n805), .A2(new_n301), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT37), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n311), .B1(new_n320), .B2(new_n803), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n301), .A2(new_n808), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n807), .A2(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT101), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n616), .A2(KEYINPUT79), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n814), .A2(new_n321), .A3(new_n325), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n813), .B(new_n805), .C1(new_n815), .C2(new_n310), .ZN(new_n816));
  INV_X1    g0616(.A(new_n805), .ZN(new_n817));
  AOI21_X1  g0617(.A(KEYINPUT101), .B1(new_n329), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n812), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(KEYINPUT38), .B(new_n812), .C1(new_n816), .C2(new_n818), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n685), .B(new_n686), .C1(new_n690), .C2(new_n641), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n771), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n452), .A2(KEYINPUT99), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT99), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n450), .A2(new_n827), .A3(new_n451), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n451), .A2(new_n626), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n376), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n826), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n450), .A2(new_n830), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n825), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n823), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT40), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n311), .B(new_n803), .C1(new_n617), .C2(new_n613), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT102), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n301), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n323), .A2(KEYINPUT102), .A3(new_n281), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n809), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n843));
  OAI21_X1  g0643(.A(KEYINPUT104), .B1(new_n810), .B2(new_n811), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT104), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n809), .A2(new_n845), .A3(new_n808), .A4(new_n301), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT103), .B1(new_n842), .B2(KEYINPUT37), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n838), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n820), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n822), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n834), .A2(new_n851), .A3(KEYINPUT40), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT105), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT105), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n834), .A2(new_n851), .A3(new_n854), .A4(KEYINPUT40), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n837), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n454), .A2(new_n824), .ZN(new_n857));
  OAI21_X1  g0657(.A(G330), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(KEYINPUT106), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n858), .A2(KEYINPUT106), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n859), .B(new_n860), .C1(new_n857), .C2(new_n856), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT39), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n851), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n821), .A2(KEYINPUT39), .A3(new_n822), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n626), .B1(new_n826), .B2(new_n828), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n437), .A2(new_n626), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n772), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT98), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT98), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n772), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n871), .A2(new_n873), .B1(new_n832), .B2(new_n833), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n823), .A2(new_n874), .B1(new_n617), .B2(new_n624), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n867), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n444), .A2(new_n452), .A3(new_n662), .A4(new_n671), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n619), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n876), .B(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n801), .B1(new_n862), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n879), .B2(new_n862), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n459), .A2(KEYINPUT35), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n459), .A2(KEYINPUT35), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n882), .A2(G116), .A3(new_n218), .A4(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT36), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n370), .B(new_n215), .C1(G58), .C2(G68), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n202), .A2(G50), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT97), .Z(new_n888));
  OAI211_X1 g0688(.A(G1), .B(new_n249), .C1(new_n886), .C2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n881), .A2(new_n885), .A3(new_n889), .ZN(G367));
  AND2_X1   g0690(.A1(new_n239), .A2(new_n755), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n752), .B1(new_n212), .B2(new_n414), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n704), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n713), .A2(new_n547), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(KEYINPUT46), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT110), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n718), .A2(new_n731), .B1(new_n709), .B2(new_n734), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n337), .B(new_n897), .C1(G97), .C2(new_n716), .ZN(new_n898));
  XOR2_X1   g0698(.A(KEYINPUT111), .B(G317), .Z(new_n899));
  OAI22_X1  g0699(.A1(new_n899), .A2(new_n724), .B1(new_n707), .B2(new_n582), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(G303), .B2(new_n721), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n894), .A2(KEYINPUT46), .B1(G107), .B2(new_n736), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n896), .A2(new_n898), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n718), .A2(new_n783), .B1(new_n720), .B2(new_n392), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n728), .A2(new_n202), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT112), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n715), .A2(new_n370), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n201), .A2(new_n713), .B1(new_n707), .B2(new_n784), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n909), .B(new_n910), .C1(G137), .C2(new_n725), .ZN(new_n911));
  INV_X1    g0711(.A(new_n709), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n275), .B1(new_n912), .B2(G50), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n908), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n907), .A2(KEYINPUT112), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n903), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT47), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n893), .B1(new_n917), .B2(new_n746), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n530), .A2(new_n641), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n525), .A2(new_n531), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n525), .B2(new_n919), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n918), .B1(new_n921), .B2(new_n761), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n701), .B(KEYINPUT109), .Z(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n500), .B(new_n535), .C1(new_n659), .C2(new_n534), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT108), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n607), .B2(new_n647), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT45), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n927), .A2(new_n928), .A3(new_n648), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n928), .B1(new_n927), .B2(new_n648), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n927), .A2(new_n648), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT44), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n927), .A2(KEYINPUT44), .A3(new_n648), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n643), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n931), .A2(new_n936), .A3(new_n643), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n646), .B1(new_n642), .B2(new_n645), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(new_n631), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n698), .B2(new_n941), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n696), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n654), .B(KEYINPUT41), .Z(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n924), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n927), .A2(new_n646), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT42), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n500), .B1(new_n927), .B2(new_n640), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n659), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT107), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT43), .B1(new_n921), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n921), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(KEYINPUT43), .B2(new_n921), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n950), .A2(new_n952), .A3(new_n957), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n643), .B2(new_n927), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n643), .A2(new_n927), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n959), .A2(new_n963), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n922), .B1(new_n948), .B2(new_n965), .ZN(G387));
  NAND2_X1  g0766(.A1(new_n696), .A2(new_n943), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n695), .A2(new_n694), .A3(new_n944), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n967), .A2(new_n654), .A3(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n714), .A2(G294), .B1(new_n736), .B2(G283), .ZN(new_n970));
  INV_X1    g0770(.A(new_n707), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G322), .A2(new_n738), .B1(new_n971), .B2(G311), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n541), .B2(new_n709), .C1(new_n720), .C2(new_n899), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT48), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT114), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n974), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT49), .Z(new_n979));
  AOI21_X1  g0779(.A(new_n337), .B1(new_n725), .B2(G326), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n547), .B2(new_n715), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n728), .A2(new_n414), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G50), .B2(new_n721), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT113), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G68), .A2(new_n912), .B1(new_n725), .B2(G150), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n255), .B2(new_n707), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n275), .B1(new_n716), .B2(G97), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n370), .B2(new_n713), .C1(new_n784), .C2(new_n718), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n985), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n982), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n747), .ZN(new_n992));
  INV_X1    g0792(.A(new_n753), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n757), .A2(new_n655), .B1(new_n426), .B2(new_n650), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n235), .A2(new_n509), .ZN(new_n995));
  AOI211_X1 g0795(.A(G45), .B(new_n655), .C1(G68), .C2(G77), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n256), .A2(KEYINPUT50), .A3(new_n367), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT50), .B1(new_n256), .B2(new_n367), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n755), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n994), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n702), .B(new_n992), .C1(new_n993), .C2(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n642), .A2(new_n761), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1002), .A2(new_n1003), .B1(new_n943), .B2(new_n924), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n969), .A2(new_n1004), .ZN(G393));
  AND2_X1   g0805(.A1(new_n938), .A2(new_n939), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1006), .A2(new_n696), .A3(new_n943), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n967), .A2(new_n940), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n1008), .A3(new_n654), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n755), .A2(new_n247), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n752), .B1(new_n466), .B2(new_n212), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n707), .A2(new_n541), .B1(new_n709), .B2(new_n582), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G317), .A2(new_n738), .B1(new_n721), .B2(G311), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT52), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1012), .B(new_n1014), .C1(G116), .C2(new_n736), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G283), .A2(new_n714), .B1(new_n725), .B2(G322), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1016), .B(new_n275), .C1(new_n426), .C2(new_n715), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT115), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n718), .A2(new_n392), .B1(new_n720), .B2(new_n784), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT51), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n337), .B1(new_n728), .B2(new_n370), .C1(new_n222), .C2(new_n715), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n707), .A2(new_n367), .B1(new_n709), .B2(new_n255), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n713), .A2(new_n202), .B1(new_n724), .B2(new_n783), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1015), .A2(new_n1018), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n704), .B1(new_n1010), .B2(new_n1011), .C1(new_n1025), .C2(new_n747), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n927), .B2(new_n751), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n1006), .B2(new_n924), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1009), .A2(new_n1028), .ZN(G390));
  NAND2_X1  g0829(.A1(new_n871), .A2(new_n873), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n832), .A2(new_n833), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n866), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AND3_X1   g0834(.A1(new_n821), .A2(KEYINPUT39), .A3(new_n822), .ZN(new_n1035));
  AOI21_X1  g0835(.A(KEYINPUT39), .B1(new_n850), .B2(new_n822), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT116), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n641), .B(new_n771), .C1(new_n667), .C2(new_n670), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n869), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n450), .A2(new_n827), .A3(new_n451), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n827), .B1(new_n450), .B2(new_n451), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n829), .B1(new_n356), .B2(new_n375), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n833), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1040), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n851), .A2(new_n1033), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1031), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n691), .A2(G330), .A3(new_n771), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1037), .A2(new_n1038), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n834), .A2(G330), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n864), .A2(new_n865), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n1047), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n864), .A2(new_n865), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1047), .B1(new_n1057), .B2(new_n1034), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1038), .B1(new_n1058), .B2(new_n1051), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n444), .A2(G330), .A3(new_n452), .A4(new_n824), .ZN(new_n1060));
  AND3_X1   g0860(.A1(new_n619), .A2(new_n877), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1040), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n824), .A2(G330), .A3(new_n771), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1049), .A2(new_n1063), .ZN(new_n1064));
  AND3_X1   g0864(.A1(new_n1051), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n834), .A2(G330), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1066), .A2(new_n1067), .B1(new_n873), .B2(new_n871), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1061), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1056), .A2(new_n1059), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(KEYINPUT117), .B1(new_n1070), .B2(new_n699), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1037), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT116), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n619), .A2(new_n877), .A3(new_n1060), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1067), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1030), .B1(new_n1053), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1051), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1073), .A2(new_n1052), .A3(new_n1055), .A4(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT117), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n1080), .A3(new_n654), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1069), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1071), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1056), .A2(new_n1059), .A3(new_n923), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n796), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n714), .A2(G150), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT53), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n275), .B1(new_n971), .B2(G137), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n784), .B2(new_n728), .ZN(new_n1089));
  INV_X1    g0889(.A(G125), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n724), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(KEYINPUT54), .B(G143), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n367), .A2(new_n715), .B1(new_n709), .B2(new_n1092), .ZN(new_n1093));
  NOR4_X1   g0893(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(G128), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n718), .A2(new_n1095), .B1(new_n720), .B2(new_n789), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT118), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n715), .A2(new_n202), .B1(new_n724), .B2(new_n582), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT119), .Z(new_n1099));
  OAI221_X1 g0899(.A(new_n275), .B1(new_n728), .B2(new_n370), .C1(new_n222), .C2(new_n713), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n426), .A2(new_n707), .B1(new_n720), .B2(new_n547), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n718), .A2(new_n734), .B1(new_n709), .B2(new_n466), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1094), .A2(new_n1097), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n704), .B1(new_n256), .B2(new_n1085), .C1(new_n1104), .C2(new_n747), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT120), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n1057), .B2(new_n749), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1084), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1083), .A2(new_n1109), .ZN(G378));
  OAI22_X1  g0910(.A1(new_n718), .A2(new_n1090), .B1(new_n707), .B2(new_n789), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1092), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n714), .A2(new_n1112), .B1(new_n912), .B2(G137), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1095), .B2(new_n720), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1111), .B(new_n1114), .C1(G150), .C2(new_n736), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT59), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n716), .A2(G159), .ZN(new_n1119));
  AOI211_X1 g0919(.A(G33), .B(G41), .C1(new_n725), .C2(G124), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n905), .B1(G116), .B2(new_n738), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT122), .Z(new_n1123));
  NOR2_X1   g0923(.A1(new_n715), .A2(new_n201), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT121), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n720), .A2(new_n426), .B1(new_n709), .B2(new_n414), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n484), .B(new_n275), .C1(new_n713), .C2(new_n370), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n707), .A2(new_n466), .B1(new_n724), .B2(new_n734), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1123), .A2(new_n1125), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1131), .A2(KEYINPUT58), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n367), .B1(new_n273), .B2(G41), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(KEYINPUT58), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1121), .A2(new_n1132), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n746), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n702), .B1(new_n367), .B2(new_n796), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n397), .A2(new_n803), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n410), .B(new_n1138), .Z(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1139), .B(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1136), .B(new_n1137), .C1(new_n1142), .C2(new_n750), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n876), .A2(new_n1141), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n867), .A2(new_n875), .A3(new_n1142), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n856), .A2(new_n1145), .A3(G330), .A4(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n837), .A2(new_n853), .A3(G330), .A4(new_n855), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1146), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1142), .B1(new_n867), .B2(new_n875), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1144), .B1(new_n1152), .B2(new_n924), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1074), .B(KEYINPUT123), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1152), .B1(new_n1070), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n654), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1079), .A2(new_n1154), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(KEYINPUT57), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1153), .B1(new_n1158), .B2(new_n1160), .ZN(G375));
  NOR2_X1   g0961(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1074), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1163), .A2(new_n947), .A3(new_n1069), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1049), .A2(new_n749), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n704), .B1(G68), .B2(new_n1085), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G137), .A2(new_n721), .B1(new_n912), .B2(G150), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1125), .B(new_n1167), .C1(new_n784), .C2(new_n713), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n738), .A2(G132), .B1(new_n725), .B2(G128), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n275), .B1(new_n971), .B2(new_n1112), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(new_n367), .C2(new_n728), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n707), .A2(new_n547), .B1(new_n709), .B2(new_n426), .ZN(new_n1172));
  OR4_X1    g0972(.A1(new_n337), .A2(new_n1172), .A3(new_n909), .A4(new_n983), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n738), .A2(G294), .B1(new_n725), .B2(G303), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n466), .B2(new_n713), .C1(new_n734), .C2(new_n720), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1168), .A2(new_n1171), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1166), .B1(new_n1176), .B2(new_n746), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1165), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1162), .B2(new_n923), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1164), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT124), .ZN(G381));
  INV_X1    g0982(.A(new_n1153), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n699), .B1(new_n1159), .B2(KEYINPUT57), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1109), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n1071), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(G387), .A2(G390), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n969), .A2(new_n763), .A3(new_n1004), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(G384), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT125), .Z(new_n1194));
  OR4_X1    g0994(.A1(G381), .A2(new_n1190), .A3(new_n1191), .A4(new_n1194), .ZN(G407));
  OAI211_X1 g0995(.A(G407), .B(G213), .C1(G343), .C2(new_n1190), .ZN(G409));
  INV_X1    g0996(.A(KEYINPUT63), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1159), .A2(new_n947), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1083), .A2(new_n1109), .A3(new_n1153), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n625), .A2(G213), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n1186), .C2(new_n1189), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1076), .A2(new_n1074), .A3(KEYINPUT60), .A4(new_n1077), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n654), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1069), .A2(KEYINPUT60), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n1204), .B2(new_n1163), .ZN(new_n1205));
  OR3_X1    g1005(.A1(new_n1205), .A2(new_n799), .A3(new_n1179), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n799), .B1(new_n1205), .B2(new_n1179), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1197), .B1(new_n1201), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT126), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(G393), .A2(G396), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1192), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(G387), .A2(G390), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(G387), .A2(G390), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1191), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n625), .A2(G213), .A3(G2897), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1206), .A2(new_n1207), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(KEYINPUT61), .B(new_n1220), .C1(new_n1201), .C2(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(G375), .A2(G378), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1208), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1226), .A2(KEYINPUT63), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(KEYINPUT126), .B(new_n1197), .C1(new_n1201), .C2(new_n1208), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1211), .A2(new_n1225), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT62), .B1(new_n1201), .B2(new_n1208), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT61), .B1(new_n1201), .B2(new_n1224), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT62), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1220), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1231), .A2(new_n1237), .ZN(G405));
  NAND2_X1  g1038(.A1(new_n1227), .A2(new_n1190), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1208), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1227), .A2(new_n1190), .A3(new_n1228), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1220), .A2(KEYINPUT127), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1220), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT127), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1242), .A2(new_n1243), .A3(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1240), .A2(new_n1245), .A3(new_n1244), .A4(new_n1241), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(G402));
endmodule


