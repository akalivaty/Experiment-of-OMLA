//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OR2_X1    g0008(.A1(new_n208), .A2(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n209), .B(new_n210), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT64), .Z(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  NAND2_X1  g0024(.A1(new_n216), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT65), .Z(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G50), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n238), .B(new_n245), .ZN(G351));
  NAND2_X1  g0046(.A1(G33), .A2(G283), .ZN(new_n247));
  INV_X1    g0047(.A(G20), .ZN(new_n248));
  INV_X1    g0048(.A(G97), .ZN(new_n249));
  OAI211_X1 g0049(.A(new_n247), .B(new_n248), .C1(G33), .C2(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n211), .ZN(new_n252));
  INV_X1    g0052(.A(G116), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n250), .A2(KEYINPUT20), .A3(new_n252), .A4(new_n254), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT68), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n251), .A2(new_n261), .A3(new_n211), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(G33), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n263), .A2(G116), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n265), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n253), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n259), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT5), .B(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n264), .A2(G45), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n271), .A2(new_n273), .B1(new_n212), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n276), .B1(new_n212), .B2(new_n274), .ZN(new_n277));
  OR2_X1    g0077(.A1(KEYINPUT5), .A2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT5), .A2(G41), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n272), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n275), .A2(G270), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  OAI211_X1 g0083(.A(G264), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  OAI211_X1 g0085(.A(G257), .B(new_n285), .C1(new_n282), .C2(new_n283), .ZN(new_n286));
  OR2_X1    g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G303), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n284), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n281), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n270), .B1(G200), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(new_n293), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT21), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  AOI211_X1 g0098(.A(new_n297), .B(new_n298), .C1(new_n281), .C2(new_n292), .ZN(new_n299));
  AND3_X1   g0099(.A1(new_n281), .A2(G179), .A3(new_n292), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n270), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT83), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n298), .B1(new_n281), .B2(new_n292), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n270), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n304), .B2(new_n297), .ZN(new_n305));
  AOI211_X1 g0105(.A(KEYINPUT83), .B(KEYINPUT21), .C1(new_n303), .C2(new_n270), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n296), .B(new_n301), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT15), .B(G87), .Z(new_n309));
  INV_X1    g0109(.A(G33), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT69), .B1(new_n310), .B2(G20), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT69), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(new_n248), .A3(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n309), .A2(new_n314), .B1(G20), .B2(G77), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT8), .B(G58), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT70), .ZN(new_n317));
  NOR2_X1   g0117(.A1(G20), .A2(G33), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n315), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n251), .A2(new_n261), .A3(new_n211), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n261), .B1(new_n251), .B2(new_n211), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G77), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n320), .A2(new_n323), .B1(new_n324), .B2(new_n268), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n268), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n264), .A2(G20), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(G77), .A3(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n228), .B1(new_n287), .B2(new_n288), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n285), .ZN(new_n331));
  INV_X1    g0131(.A(G107), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT3), .B(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G1698), .ZN(new_n334));
  INV_X1    g0134(.A(G238), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n331), .B1(new_n332), .B2(new_n333), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n291), .ZN(new_n337));
  INV_X1    g0137(.A(G41), .ZN(new_n338));
  INV_X1    g0138(.A(G45), .ZN(new_n339));
  AOI21_X1  g0139(.A(G1), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(G274), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT66), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n343), .B1(new_n341), .B2(new_n344), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G244), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n337), .A2(new_n342), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G200), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n329), .B(new_n350), .C1(new_n295), .C2(new_n349), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n298), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n325), .A2(new_n328), .ZN(new_n353));
  INV_X1    g0153(.A(G179), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n337), .A2(new_n354), .A3(new_n348), .A4(new_n342), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT71), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n333), .A2(G222), .A3(new_n285), .ZN(new_n360));
  XOR2_X1   g0160(.A(KEYINPUT67), .B(G223), .Z(new_n361));
  OAI221_X1 g0161(.A(new_n360), .B1(new_n324), .B2(new_n333), .C1(new_n334), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n291), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n347), .A2(G226), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n342), .A3(new_n364), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n365), .A2(G179), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n326), .A2(G50), .A3(new_n327), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n311), .A2(new_n313), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(new_n316), .ZN(new_n369));
  OAI21_X1  g0169(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n370));
  INV_X1    g0170(.A(G150), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n319), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n323), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n268), .A2(new_n239), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n367), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n365), .A2(new_n298), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n366), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n365), .A2(G200), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT9), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT10), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n375), .A2(new_n380), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n363), .A2(G190), .A3(new_n364), .A4(new_n342), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n382), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n384), .A2(new_n379), .A3(new_n381), .A4(new_n385), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT10), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n378), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n314), .A2(G77), .B1(G20), .B2(new_n241), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT74), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n391), .A2(new_n392), .B1(G50), .B2(new_n318), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n392), .B2(new_n391), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(KEYINPUT11), .A3(new_n323), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n241), .B1(new_n264), .B2(G20), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT12), .B1(new_n265), .B2(G68), .ZN(new_n397));
  OR3_X1    g0197(.A1(new_n265), .A2(KEYINPUT12), .A3(G68), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n326), .A2(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n394), .A2(new_n323), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT11), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT14), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  OAI211_X1 g0206(.A(G226), .B(new_n285), .C1(new_n282), .C2(new_n283), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT72), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT72), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n333), .A2(new_n409), .A3(G226), .A4(new_n285), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT73), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n412), .A2(G33), .A3(G97), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G97), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT73), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n330), .A2(G1698), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n291), .ZN(new_n418));
  OAI21_X1  g0218(.A(G238), .B1(new_n345), .B2(new_n346), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n419), .A2(new_n342), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n406), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n341), .B1(new_n411), .B2(new_n416), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n342), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT13), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n405), .B(G169), .C1(new_n421), .C2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n418), .A2(new_n420), .A3(new_n406), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT13), .B1(new_n422), .B2(new_n423), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(G179), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n427), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n405), .B1(new_n430), .B2(G169), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n404), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(G200), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n426), .A2(G190), .A3(new_n427), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n400), .A2(new_n433), .A3(new_n403), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT16), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT7), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n333), .B2(G20), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n282), .A2(new_n283), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(KEYINPUT7), .A3(new_n248), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n241), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G58), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(new_n241), .ZN(new_n444));
  OAI21_X1  g0244(.A(G20), .B1(new_n444), .B2(new_n201), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n318), .A2(G159), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n437), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT7), .B1(new_n440), .B2(new_n248), .ZN(new_n449));
  NOR4_X1   g0249(.A1(new_n282), .A2(new_n283), .A3(new_n438), .A4(G20), .ZN(new_n450));
  OAI21_X1  g0250(.A(G68), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n447), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(KEYINPUT16), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n453), .A3(new_n323), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n316), .B1(new_n264), .B2(G20), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n326), .A2(new_n455), .B1(new_n268), .B2(new_n316), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n341), .A2(new_n344), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n342), .B1(new_n228), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(G226), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT75), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT75), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n333), .A2(new_n462), .A3(G226), .A4(G1698), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G87), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n333), .A2(G223), .A3(new_n285), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n461), .A2(new_n463), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n459), .B1(new_n466), .B2(new_n291), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n354), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(G169), .B2(new_n467), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT18), .B1(new_n457), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n467), .A2(G200), .ZN(new_n471));
  AOI211_X1 g0271(.A(G190), .B(new_n459), .C1(new_n466), .C2(new_n291), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n454), .B(new_n456), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT17), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n467), .A2(new_n295), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(G200), .B2(new_n467), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n457), .A2(KEYINPUT17), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n466), .A2(new_n291), .ZN(new_n479));
  INV_X1    g0279(.A(new_n459), .ZN(new_n480));
  AOI21_X1  g0280(.A(G169), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI211_X1 g0281(.A(G179), .B(new_n459), .C1(new_n466), .C2(new_n291), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n454), .A2(new_n456), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT18), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n470), .A2(new_n475), .A3(new_n478), .A4(new_n486), .ZN(new_n487));
  NOR4_X1   g0287(.A1(new_n359), .A2(new_n390), .A3(new_n436), .A4(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(G250), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n489));
  OAI211_X1 g0289(.A(G244), .B(new_n285), .C1(new_n282), .C2(new_n283), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n247), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n493));
  INV_X1    g0293(.A(G244), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n287), .B2(new_n288), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(new_n495), .B2(new_n285), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n291), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n275), .A2(G257), .B1(new_n277), .B2(new_n280), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(G190), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT80), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT80), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n497), .A2(new_n501), .A3(G190), .A4(new_n498), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  NOR2_X1   g0304(.A1(G97), .A2(G107), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT76), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n507));
  MUX2_X1   g0307(.A(new_n506), .B(G97), .S(KEYINPUT6), .Z(new_n508));
  XNOR2_X1  g0308(.A(G97), .B(G107), .ZN(new_n509));
  OAI211_X1 g0309(.A(G20), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n318), .A2(G77), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n332), .B1(new_n439), .B2(new_n441), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n323), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n265), .B(new_n266), .C1(new_n321), .C2(new_n322), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT77), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT77), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n263), .A2(new_n517), .A3(new_n265), .A4(new_n266), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n518), .A3(G97), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n268), .A2(new_n249), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n514), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n497), .A2(new_n498), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT79), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(G200), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n271), .A2(new_n273), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n526), .A2(G257), .A3(new_n341), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n280), .A2(new_n277), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n493), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n490), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n333), .A2(KEYINPUT4), .A3(G244), .A4(new_n285), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n531), .A2(new_n532), .A3(new_n247), .A4(new_n489), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n529), .B1(new_n291), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G200), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT79), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n503), .A2(new_n522), .A3(new_n525), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n523), .A2(new_n298), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n497), .A2(new_n354), .A3(new_n498), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n521), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n542));
  OAI211_X1 g0342(.A(G250), .B(new_n285), .C1(new_n282), .C2(new_n283), .ZN(new_n543));
  INV_X1    g0343(.A(G294), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n542), .B(new_n543), .C1(new_n310), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n291), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n275), .A2(G264), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n528), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n298), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n545), .A2(new_n291), .B1(G264), .B2(new_n275), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(new_n354), .A3(new_n528), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT25), .ZN(new_n553));
  AOI211_X1 g0353(.A(G107), .B(new_n265), .C1(KEYINPUT85), .C2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(KEYINPUT85), .ZN(new_n555));
  XOR2_X1   g0355(.A(new_n554), .B(new_n555), .Z(new_n556));
  OAI211_X1 g0356(.A(new_n248), .B(G87), .C1(new_n282), .C2(new_n283), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT22), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT22), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n333), .A2(new_n559), .A3(new_n248), .A4(G87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n310), .A2(new_n253), .A3(G20), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT84), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n248), .B2(G107), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT23), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT23), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n563), .B(new_n566), .C1(new_n248), .C2(G107), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n562), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT24), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n561), .A2(new_n571), .A3(new_n568), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n556), .B1(new_n573), .B2(new_n323), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n516), .A2(new_n518), .A3(G107), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n552), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT82), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n577), .B(new_n578), .C1(new_n368), .C2(new_n249), .ZN(new_n579));
  INV_X1    g0379(.A(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n505), .A2(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n415), .A2(new_n413), .A3(KEYINPUT19), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(G20), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n249), .B1(new_n311), .B2(new_n313), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT82), .B1(new_n584), .B2(KEYINPUT19), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n333), .A2(new_n248), .A3(G68), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n579), .A2(new_n583), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n323), .ZN(new_n588));
  INV_X1    g0388(.A(new_n309), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n268), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n516), .A2(new_n518), .A3(new_n309), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT81), .ZN(new_n593));
  OAI21_X1  g0393(.A(G250), .B1(new_n339), .B2(G1), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n291), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n341), .A2(KEYINPUT81), .A3(G250), .A4(new_n272), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n595), .A2(new_n596), .B1(new_n277), .B2(new_n273), .ZN(new_n597));
  OAI211_X1 g0397(.A(G244), .B(G1698), .C1(new_n282), .C2(new_n283), .ZN(new_n598));
  OAI211_X1 g0398(.A(G238), .B(new_n285), .C1(new_n282), .C2(new_n283), .ZN(new_n599));
  NAND2_X1  g0399(.A1(G33), .A2(G116), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n291), .ZN(new_n602));
  AOI21_X1  g0402(.A(G169), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n597), .A2(new_n602), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n603), .B1(new_n354), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n592), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n597), .A2(new_n602), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n535), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n597), .A2(new_n602), .A3(new_n295), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n587), .A2(new_n323), .B1(new_n268), .B2(new_n589), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n516), .A2(new_n518), .A3(G87), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n561), .A2(new_n571), .A3(new_n568), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n571), .B1(new_n561), .B2(new_n568), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n323), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n554), .B(new_n555), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n575), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n548), .A2(G200), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n295), .B2(new_n548), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n576), .A2(new_n614), .A3(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n308), .A2(new_n488), .A3(new_n541), .A4(new_n623), .ZN(G372));
  NAND2_X1  g0424(.A1(new_n386), .A2(new_n388), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n475), .A2(new_n478), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n435), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n432), .B2(new_n356), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n470), .A2(new_n486), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n625), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n631), .A2(new_n377), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n614), .A2(new_n622), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n541), .B(new_n633), .C1(new_n634), .C2(new_n576), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT26), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n614), .B2(new_n540), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n588), .A2(new_n590), .A3(new_n612), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n638), .A2(new_n610), .B1(new_n592), .B2(new_n605), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n521), .A2(new_n538), .A3(new_n539), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(KEYINPUT26), .A3(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n637), .A2(new_n641), .B1(new_n592), .B2(new_n605), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n488), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n632), .A2(new_n644), .ZN(G369));
  NAND3_X1  g0445(.A1(new_n264), .A2(new_n248), .A3(G13), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(G213), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G343), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n270), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n634), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT86), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n653), .B(KEYINPUT86), .C1(new_n307), .C2(new_n652), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G330), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n619), .A2(new_n551), .A3(new_n549), .ZN(new_n658));
  INV_X1    g0458(.A(new_n651), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n574), .B2(new_n575), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n660), .B2(new_n622), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n576), .A2(new_n659), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n657), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n663), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n634), .A2(new_n659), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n662), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n665), .A2(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n206), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n581), .A2(G116), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n214), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT29), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n643), .B2(new_n659), .ZN(new_n681));
  AOI211_X1 g0481(.A(KEYINPUT29), .B(new_n651), .C1(new_n635), .C2(new_n642), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n623), .A2(new_n308), .A3(new_n541), .A4(new_n659), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n300), .A2(new_n534), .A3(new_n550), .A4(new_n604), .ZN(new_n686));
  NOR2_X1   g0486(.A1(KEYINPUT87), .A2(KEYINPUT30), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n607), .A2(KEYINPUT88), .B1(new_n497), .B2(new_n498), .ZN(new_n689));
  AOI21_X1  g0489(.A(G179), .B1(new_n281), .B2(new_n292), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT88), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n597), .A2(new_n602), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n689), .A2(new_n548), .A3(new_n690), .A4(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n550), .A2(new_n602), .A3(new_n597), .ZN(new_n694));
  INV_X1    g0494(.A(new_n687), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n300), .A3(new_n534), .A4(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n688), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n697), .A2(KEYINPUT31), .A3(new_n651), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT31), .B1(new_n697), .B2(new_n651), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n684), .B1(new_n685), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n683), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n679), .B1(new_n702), .B2(G1), .ZN(G364));
  INV_X1    g0503(.A(G13), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G20), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n264), .B1(new_n705), .B2(G45), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n675), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT89), .Z(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n673), .A2(new_n440), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n710), .A2(G355), .B1(new_n253), .B2(new_n673), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n440), .A2(new_n206), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT90), .Z(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(G45), .B2(new_n214), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n245), .A2(new_n339), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G13), .A2(G33), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n211), .B1(G20), .B2(new_n298), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n709), .B1(new_n716), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n248), .A2(new_n354), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G190), .A2(G200), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n248), .A2(G179), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n295), .A3(G200), .ZN(new_n727));
  OAI221_X1 g0527(.A(new_n333), .B1(new_n725), .B2(new_n324), .C1(new_n332), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n724), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G159), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n726), .A2(G190), .A3(G200), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n731), .A2(KEYINPUT32), .B1(new_n733), .B2(G87), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n723), .A2(G200), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n295), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n734), .B1(KEYINPUT32), .B2(new_n731), .C1(new_n239), .C2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n723), .A2(G190), .A3(new_n535), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT91), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI211_X1 g0541(.A(new_n728), .B(new_n738), .C1(G58), .C2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n735), .A2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n248), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n744), .A2(new_n241), .B1(new_n249), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT92), .ZN(new_n748));
  INV_X1    g0548(.A(G303), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n732), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G283), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n746), .A2(new_n544), .B1(new_n727), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n750), .B(new_n752), .C1(G326), .C2(new_n736), .ZN(new_n753));
  INV_X1    g0553(.A(new_n739), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n754), .A2(G322), .B1(new_n730), .B2(G329), .ZN(new_n755));
  INV_X1    g0555(.A(G311), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n755), .B(new_n440), .C1(new_n756), .C2(new_n725), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT33), .B(G317), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n759), .A2(KEYINPUT93), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n744), .B1(KEYINPUT93), .B2(new_n759), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n742), .A2(new_n748), .B1(new_n753), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n720), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n722), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n656), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(new_n766), .B2(new_n719), .ZN(new_n767));
  INV_X1    g0567(.A(new_n657), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n707), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n656), .A2(G330), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n767), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(G396));
  INV_X1    g0573(.A(KEYINPUT95), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n356), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT95), .A4(new_n355), .ZN(new_n776));
  AND3_X1   g0576(.A1(new_n775), .A2(new_n351), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(KEYINPUT26), .B1(new_n639), .B2(new_n640), .ZN(new_n778));
  AND4_X1   g0578(.A1(KEYINPUT26), .A2(new_n640), .A3(new_n606), .A4(new_n613), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n606), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AND4_X1   g0580(.A1(G190), .A2(new_n546), .A3(new_n528), .A4(new_n547), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n535), .B1(new_n550), .B2(new_n528), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n574), .A2(new_n575), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n639), .A2(new_n537), .A3(new_n540), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n634), .A2(new_n576), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n659), .B(new_n777), .C1(new_n780), .C2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n651), .B1(new_n635), .B2(new_n642), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n353), .A2(new_n651), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n775), .A2(new_n351), .A3(new_n790), .A4(new_n776), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n356), .A2(new_n659), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n788), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n701), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT96), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n794), .A2(KEYINPUT97), .A3(new_n795), .ZN(new_n798));
  AOI21_X1  g0598(.A(KEYINPUT97), .B1(new_n794), .B2(new_n795), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n707), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n725), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n736), .A2(G137), .B1(new_n802), .B2(G159), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n371), .B2(new_n744), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G143), .B2(new_n741), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n807));
  INV_X1    g0607(.A(new_n746), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n808), .A2(G58), .B1(new_n733), .B2(G50), .ZN(new_n809));
  INV_X1    g0609(.A(new_n727), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G68), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n440), .B1(new_n730), .B2(G132), .ZN(new_n812));
  AND3_X1   g0612(.A1(new_n809), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n806), .A2(new_n807), .A3(new_n813), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n746), .A2(new_n249), .B1(new_n739), .B2(new_n544), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT94), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n440), .B1(new_n729), .B2(new_n756), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G116), .B2(new_n802), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n727), .A2(new_n580), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G303), .B2(new_n736), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n743), .A2(G283), .B1(new_n733), .B2(G107), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n816), .A2(new_n818), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n764), .B1(new_n814), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n720), .A2(new_n717), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n709), .B(new_n823), .C1(new_n324), .C2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n793), .B2(new_n718), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n801), .A2(new_n826), .ZN(G384));
  NOR2_X1   g0627(.A1(new_n705), .A2(new_n264), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n685), .A2(new_n700), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n488), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT101), .Z(new_n831));
  INV_X1    g0631(.A(new_n649), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n484), .B1(new_n483), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n833), .A2(KEYINPUT37), .A3(new_n473), .ZN(new_n834));
  AOI21_X1  g0634(.A(KEYINPUT37), .B1(new_n833), .B2(new_n473), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n484), .A2(new_n832), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n487), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n836), .A2(new_n839), .A3(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT98), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT98), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n836), .A2(new_n839), .A3(new_n842), .A4(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n836), .A2(new_n839), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n841), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n659), .B1(new_n400), .B2(new_n403), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n432), .A2(new_n435), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n848), .B1(new_n431), .B2(new_n429), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n829), .A2(new_n793), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT40), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n483), .A2(new_n484), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(new_n837), .A3(new_n473), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n837), .A3(KEYINPUT99), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT37), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT100), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n833), .B(new_n473), .C1(KEYINPUT99), .C2(new_n861), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n860), .B1(new_n859), .B2(new_n862), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n837), .B1(new_n629), .B2(new_n626), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n840), .B1(new_n866), .B2(KEYINPUT38), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n829), .A2(KEYINPUT40), .A3(new_n852), .A4(new_n793), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n854), .A2(new_n855), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n684), .B1(new_n831), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n870), .B2(new_n831), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT39), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n859), .A2(new_n862), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n874), .A2(KEYINPUT100), .B1(new_n487), .B2(new_n838), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT38), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n840), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n873), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n432), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n659), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n841), .A2(new_n846), .A3(KEYINPUT39), .A4(new_n843), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n852), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n775), .A2(new_n776), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n659), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n885), .B1(new_n788), .B2(new_n887), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n888), .A2(new_n847), .B1(new_n630), .B2(new_n649), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n488), .B1(new_n681), .B2(new_n682), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n632), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n890), .B(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n828), .B1(new_n872), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n872), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n213), .A2(new_n253), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT35), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n898), .B2(new_n897), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT36), .Z(new_n901));
  OAI21_X1  g0701(.A(G77), .B1(new_n443), .B2(new_n241), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n240), .B1(new_n214), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(G1), .A3(new_n704), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n895), .A2(new_n901), .A3(new_n904), .ZN(G367));
  NOR2_X1   g0705(.A1(new_n638), .A2(new_n659), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT102), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n907), .A2(new_n606), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n639), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n719), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n713), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n721), .B1(new_n206), .B2(new_n589), .C1(new_n911), .C2(new_n234), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n708), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n732), .A2(new_n253), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n914), .A2(KEYINPUT46), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n915), .A2(KEYINPUT106), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(KEYINPUT106), .ZN(new_n917));
  AOI22_X1  g0717(.A1(G294), .A2(new_n743), .B1(new_n736), .B2(G311), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n808), .A2(G107), .B1(new_n810), .B2(G97), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(KEYINPUT107), .B(G317), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n440), .B1(new_n729), .B2(new_n921), .C1(new_n751), .C2(new_n725), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n923), .B1(KEYINPUT46), .B2(new_n914), .C1(new_n749), .C2(new_n740), .ZN(new_n924));
  INV_X1    g0724(.A(G137), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n725), .A2(new_n239), .B1(new_n729), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(G150), .B2(new_n754), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n746), .A2(new_n241), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(G58), .B2(new_n733), .ZN(new_n929));
  AOI22_X1  g0729(.A1(G143), .A2(new_n736), .B1(new_n743), .B2(G159), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n727), .A2(new_n324), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n932), .A2(new_n440), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT108), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n920), .A2(new_n924), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT47), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n913), .B1(new_n936), .B2(new_n720), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n910), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n706), .B(KEYINPUT105), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT44), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n541), .B1(new_n522), .B2(new_n659), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n640), .A2(new_n651), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n941), .B1(new_n671), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n944), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n670), .A2(KEYINPUT44), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n671), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT45), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n670), .B2(new_n946), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n664), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n948), .A2(new_n665), .A3(new_n952), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n657), .B1(KEYINPUT104), .B2(new_n669), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n666), .A2(new_n668), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n657), .A2(KEYINPUT104), .A3(new_n669), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n960), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n962), .A2(new_n957), .B1(new_n666), .B2(new_n668), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n702), .B1(new_n956), .B2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n674), .B(KEYINPUT41), .Z(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n940), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n946), .A2(new_n669), .A3(KEYINPUT42), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n540), .B1(new_n942), .B2(new_n658), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n659), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT42), .B1(new_n946), .B2(new_n669), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n908), .A2(new_n909), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n976), .B1(new_n974), .B2(new_n977), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n665), .A2(new_n946), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(KEYINPUT103), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n981), .A2(KEYINPUT103), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n980), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n938), .B1(new_n969), .B2(new_n986), .ZN(G387));
  INV_X1    g0787(.A(new_n710), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n988), .A2(new_n676), .B1(G107), .B2(new_n206), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n317), .A2(G50), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT50), .ZN(new_n991));
  AOI21_X1  g0791(.A(G45), .B1(G68), .B2(G77), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(new_n676), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n911), .B1(new_n231), .B2(G45), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n989), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n721), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n708), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n725), .A2(new_n241), .B1(new_n729), .B2(new_n371), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n440), .B(new_n998), .C1(G50), .C2(new_n754), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n733), .A2(G77), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n589), .A2(new_n746), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n316), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1001), .B1(new_n1002), .B2(new_n743), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n736), .A2(G159), .B1(new_n810), .B2(G97), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n999), .A2(new_n1000), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n333), .B1(new_n730), .B2(G326), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n736), .A2(G322), .B1(new_n802), .B2(G303), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n756), .B2(new_n744), .C1(new_n740), .C2(new_n921), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT48), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n808), .A2(G283), .B1(new_n733), .B2(G294), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT49), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1006), .B1(new_n253), .B2(new_n727), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1005), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n997), .B1(new_n1017), .B2(new_n720), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n719), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(new_n666), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT110), .Z(new_n1021));
  NAND2_X1  g0821(.A1(new_n964), .A2(new_n702), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(new_n675), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n964), .A2(new_n702), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n964), .A2(new_n940), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT109), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(G393));
  NAND2_X1  g0829(.A1(new_n956), .A2(KEYINPUT111), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT111), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n954), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n940), .A3(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n721), .B1(new_n249), .B2(new_n206), .C1(new_n911), .C2(new_n238), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n708), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n736), .A2(G317), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n756), .B2(new_n739), .ZN(new_n1037));
  XOR2_X1   g0837(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n733), .A2(G283), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n727), .A2(new_n332), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n333), .B(new_n1043), .C1(G322), .C2(new_n730), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n808), .A2(G116), .B1(new_n802), .B2(G294), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n749), .B2(new_n744), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT113), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G150), .A2(new_n736), .B1(new_n754), .B2(G159), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT51), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n732), .A2(new_n241), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n746), .A2(new_n324), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(G50), .C2(new_n743), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n440), .B(new_n819), .C1(G143), .C2(new_n730), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(new_n317), .C2(new_n725), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1045), .A2(new_n1048), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1035), .B1(new_n1056), .B2(new_n720), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n944), .B2(new_n1019), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1023), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n674), .B1(new_n956), .B2(new_n1022), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1033), .B(new_n1058), .C1(new_n1059), .C2(new_n1060), .ZN(G390));
  NAND4_X1  g0861(.A1(new_n829), .A2(G330), .A3(new_n852), .A4(new_n793), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n881), .B1(new_n877), .B2(new_n878), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n788), .A2(new_n887), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT114), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT114), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n788), .A2(new_n1067), .A3(new_n887), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1064), .B1(new_n1069), .B2(new_n852), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n882), .B1(new_n1065), .B2(new_n852), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n879), .B2(new_n883), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1063), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n488), .A2(new_n701), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n891), .A2(new_n632), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n829), .A2(G330), .A3(new_n793), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n885), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1065), .B1(new_n1078), .B2(new_n1063), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1066), .A2(new_n1077), .A3(new_n1062), .A4(new_n1068), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1075), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AND3_X1   g0881(.A1(new_n788), .A2(new_n1067), .A3(new_n887), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1067), .B1(new_n788), .B2(new_n887), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n852), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n874), .A2(KEYINPUT100), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n839), .A3(new_n876), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n878), .B1(new_n1086), .B2(new_n845), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1087), .A2(new_n882), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n883), .B1(new_n1087), .B2(KEYINPUT39), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1065), .A2(new_n852), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n881), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1089), .A2(new_n1093), .A3(new_n1062), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1073), .A2(new_n1081), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(KEYINPUT115), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT115), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1073), .A2(new_n1094), .A3(new_n1081), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1073), .A2(new_n1094), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1081), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n675), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n744), .A2(new_n332), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1052), .B(new_n1104), .C1(G283), .C2(new_n736), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n733), .A2(G87), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n725), .A2(new_n249), .B1(new_n729), .B2(new_n544), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n333), .B(new_n1107), .C1(G116), .C2(new_n754), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n811), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(G128), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n737), .A2(new_n1110), .B1(new_n727), .B2(new_n239), .ZN(new_n1111));
  INV_X1    g0911(.A(G159), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n744), .A2(new_n925), .B1(new_n1112), .B2(new_n746), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n732), .A2(new_n371), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n440), .B1(new_n802), .B2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n754), .A2(G132), .B1(new_n730), .B2(G125), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1114), .A2(new_n1117), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n764), .B1(new_n1109), .B2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n709), .B(new_n1123), .C1(new_n316), .C2(new_n824), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1090), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(new_n718), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1073), .A2(new_n940), .A3(new_n1094), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(KEYINPUT116), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT116), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1073), .A2(new_n1094), .A3(new_n1129), .A4(new_n940), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1103), .A2(new_n1126), .A3(new_n1131), .ZN(G378));
  AOI211_X1 g0932(.A(G33), .B(G41), .C1(new_n730), .C2(G124), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n754), .A2(G128), .B1(new_n802), .B2(G137), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n732), .B2(new_n1118), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G150), .A2(new_n808), .B1(new_n736), .B2(G125), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT119), .Z(new_n1137));
  AOI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(G132), .C2(new_n743), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT59), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1133), .B1(new_n1112), .B2(new_n727), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1139), .B2(new_n1138), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n249), .A2(new_n744), .B1(new_n737), .B2(new_n253), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n727), .A2(new_n443), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1142), .A2(new_n928), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n802), .A2(new_n309), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n754), .A2(G107), .B1(new_n730), .B2(G283), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n440), .A2(new_n338), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n733), .B2(G77), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT118), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT58), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1147), .B(new_n239), .C1(G33), .C2(G41), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n720), .B1(new_n1141), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT120), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n375), .A2(new_n832), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT121), .Z(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  XOR2_X1   g0960(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n389), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n389), .A2(new_n1162), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1160), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1165), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n1159), .A3(new_n1163), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n717), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n824), .A2(new_n239), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1157), .A2(new_n707), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1169), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n870), .B2(G330), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT40), .B1(new_n847), .B2(new_n853), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1086), .A2(new_n845), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n868), .B1(new_n1177), .B2(new_n840), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1176), .A2(new_n1178), .A3(new_n684), .A4(new_n1169), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n890), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n854), .A2(new_n855), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n867), .A2(new_n869), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(G330), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n1169), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n884), .A2(new_n889), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n870), .A2(G330), .A3(new_n1174), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1180), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1173), .B1(new_n1188), .B2(new_n940), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1075), .B(KEYINPUT122), .Z(new_n1190));
  NAND2_X1  g0990(.A1(new_n1099), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT57), .B1(new_n1191), .B2(new_n1188), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1190), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT123), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1180), .A2(new_n1187), .A3(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(KEYINPUT123), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(KEYINPUT57), .A3(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n674), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1189), .B1(new_n1192), .B2(new_n1199), .ZN(G375));
  NAND2_X1  g1000(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1075), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n968), .A3(new_n1101), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n709), .B1(new_n241), .B2(new_n824), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G116), .A2(new_n743), .B1(new_n736), .B2(G294), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n249), .B2(new_n732), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G107), .A2(new_n802), .B1(new_n730), .B2(G303), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n440), .C1(new_n751), .C2(new_n739), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1207), .A2(new_n1209), .A3(new_n932), .A4(new_n1001), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n333), .B1(new_n729), .B2(new_n1110), .C1(new_n371), .C2(new_n725), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1143), .B1(G50), .B2(new_n808), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n1112), .B2(new_n732), .C1(new_n744), .C2(new_n1118), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1211), .B(new_n1213), .C1(G137), .C2(new_n741), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n736), .A2(G132), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT124), .Z(new_n1216));
  AOI21_X1  g1016(.A(new_n1210), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1205), .B1(new_n764), .B2(new_n1217), .C1(new_n852), .C2(new_n718), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1202), .B2(new_n939), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1204), .A2(new_n1220), .ZN(G381));
  INV_X1    g1021(.A(G390), .ZN(new_n1222));
  INV_X1    g1022(.A(G384), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1026), .A2(new_n772), .A3(new_n1028), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1224), .A2(G387), .A3(G381), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1131), .A2(new_n1126), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1228));
  INV_X1    g1028(.A(G375), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(new_n1228), .A3(new_n1229), .ZN(G407));
  NAND2_X1  g1030(.A1(new_n650), .A2(G213), .ZN(new_n1231));
  OR3_X1    g1031(.A1(G375), .A2(G378), .A3(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(G407), .A2(new_n1232), .A3(G213), .ZN(G409));
  NAND2_X1  g1033(.A1(new_n966), .A2(new_n968), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n939), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n986), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1235), .A2(new_n1236), .B1(new_n910), .B2(new_n937), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(G390), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1222), .A2(G387), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G393), .A2(G396), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1241), .A2(new_n1225), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT126), .B1(new_n1237), .B2(G390), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1240), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1241), .A2(new_n1225), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1245), .A2(new_n1238), .A3(new_n1239), .A4(KEYINPUT126), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G378), .B(new_n1189), .C1(new_n1192), .C2(new_n1199), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1188), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1194), .A2(new_n967), .A3(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1196), .A2(new_n940), .A3(new_n1197), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1172), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1228), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1248), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT60), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1203), .B1(new_n1255), .B2(new_n1081), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1202), .A2(KEYINPUT60), .A3(new_n1075), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n674), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1220), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1223), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(G384), .A3(new_n1220), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1254), .A2(new_n1231), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT125), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT125), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1254), .A2(new_n1266), .A3(new_n1231), .A4(new_n1263), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT62), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1254), .A2(new_n1231), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n650), .A2(G213), .A3(G2897), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1262), .B(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT61), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1264), .A2(KEYINPUT62), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1247), .B1(new_n1268), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1265), .A2(new_n1276), .A3(new_n1267), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1264), .A2(new_n1276), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .A4(new_n1272), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1275), .A2(new_n1280), .ZN(G405));
  OAI21_X1  g1081(.A(new_n1262), .B1(new_n1229), .B2(G378), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(G375), .A2(new_n1263), .A3(new_n1228), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1247), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT127), .B1(new_n1229), .B2(G378), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1279), .A2(new_n1283), .A3(new_n1282), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1286), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(G402));
endmodule


