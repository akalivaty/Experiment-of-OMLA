

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588;

  XNOR2_X1 U322 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n390) );
  XNOR2_X1 U323 ( .A(n339), .B(KEYINPUT65), .ZN(n551) );
  XOR2_X1 U324 ( .A(n391), .B(n390), .Z(n290) );
  XNOR2_X1 U325 ( .A(n332), .B(n365), .ZN(n333) );
  XNOR2_X1 U326 ( .A(n387), .B(KEYINPUT48), .ZN(n388) );
  XNOR2_X1 U327 ( .A(n334), .B(n333), .ZN(n336) );
  XNOR2_X1 U328 ( .A(n389), .B(n388), .ZN(n532) );
  XNOR2_X1 U329 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n433) );
  XNOR2_X1 U330 ( .A(n434), .B(n433), .ZN(n452) );
  INV_X1 U331 ( .A(G190GAT), .ZN(n453) );
  XOR2_X1 U332 ( .A(KEYINPUT28), .B(n464), .Z(n536) );
  XNOR2_X1 U333 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U334 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT94), .B(KEYINPUT90), .Z(n292) );
  XNOR2_X1 U336 ( .A(G190GAT), .B(G218GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n295) );
  XNOR2_X1 U338 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n293), .B(KEYINPUT91), .ZN(n294) );
  XOR2_X1 U340 ( .A(n295), .B(n294), .Z(n297) );
  NAND2_X1 U341 ( .A1(G226GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n308) );
  XOR2_X1 U343 ( .A(G64GAT), .B(G92GAT), .Z(n299) );
  XNOR2_X1 U344 ( .A(G176GAT), .B(G204GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n328) );
  XOR2_X1 U346 ( .A(G211GAT), .B(KEYINPUT82), .Z(n301) );
  XNOR2_X1 U347 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n425) );
  XOR2_X1 U349 ( .A(n328), .B(n425), .Z(n306) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G36GAT), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n302), .B(G8GAT), .ZN(n309) );
  XOR2_X1 U352 ( .A(G183GAT), .B(KEYINPUT17), .Z(n304) );
  XNOR2_X1 U353 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n304), .B(n303), .ZN(n439) );
  XNOR2_X1 U355 ( .A(n309), .B(n439), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n523) );
  XOR2_X1 U358 ( .A(n309), .B(KEYINPUT67), .Z(n311) );
  NAND2_X1 U359 ( .A1(G229GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U361 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n313) );
  XNOR2_X1 U362 ( .A(G113GAT), .B(G197GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U364 ( .A(n315), .B(n314), .Z(n317) );
  XOR2_X1 U365 ( .A(G141GAT), .B(G22GAT), .Z(n417) );
  XOR2_X1 U366 ( .A(G15GAT), .B(G1GAT), .Z(n355) );
  XNOR2_X1 U367 ( .A(n417), .B(n355), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U369 ( .A(KEYINPUT7), .B(G50GAT), .Z(n319) );
  XNOR2_X1 U370 ( .A(G43GAT), .B(G29GAT), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U372 ( .A(KEYINPUT8), .B(n320), .ZN(n376) );
  XNOR2_X1 U373 ( .A(n321), .B(n376), .ZN(n549) );
  XOR2_X1 U374 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n323) );
  NAND2_X1 U375 ( .A1(G230GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n325) );
  INV_X1 U377 ( .A(KEYINPUT32), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n330) );
  XOR2_X1 U379 ( .A(G78GAT), .B(G148GAT), .Z(n327) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n429) );
  XNOR2_X1 U382 ( .A(n429), .B(n328), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U384 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XNOR2_X1 U385 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n331), .B(KEYINPUT13), .ZN(n356) );
  XOR2_X1 U387 ( .A(n435), .B(n356), .Z(n332) );
  XOR2_X1 U388 ( .A(G99GAT), .B(G85GAT), .Z(n365) );
  INV_X1 U389 ( .A(n336), .ZN(n383) );
  INV_X1 U390 ( .A(KEYINPUT41), .ZN(n335) );
  NAND2_X1 U391 ( .A1(n383), .A2(n335), .ZN(n338) );
  NAND2_X1 U392 ( .A1(n336), .A2(KEYINPUT41), .ZN(n337) );
  NAND2_X1 U393 ( .A1(n338), .A2(n337), .ZN(n339) );
  NAND2_X1 U394 ( .A1(n549), .A2(n551), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n340), .B(KEYINPUT46), .ZN(n361) );
  XOR2_X1 U396 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n342) );
  XNOR2_X1 U397 ( .A(G64GAT), .B(KEYINPUT76), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n354) );
  XOR2_X1 U399 ( .A(G211GAT), .B(G127GAT), .Z(n344) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(G71GAT), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n344), .B(n343), .ZN(n352) );
  XOR2_X1 U402 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n346) );
  XNOR2_X1 U403 ( .A(KEYINPUT15), .B(KEYINPUT75), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U405 ( .A(G155GAT), .B(G78GAT), .Z(n348) );
  XNOR2_X1 U406 ( .A(G22GAT), .B(G8GAT), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U408 ( .A(n350), .B(n349), .Z(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n360) );
  XOR2_X1 U411 ( .A(n356), .B(n355), .Z(n358) );
  NAND2_X1 U412 ( .A1(G231GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n472) );
  NAND2_X1 U415 ( .A1(n361), .A2(n472), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n362), .B(KEYINPUT113), .ZN(n378) );
  XOR2_X1 U417 ( .A(KEYINPUT10), .B(KEYINPUT72), .Z(n364) );
  XNOR2_X1 U418 ( .A(KEYINPUT71), .B(KEYINPUT66), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n375) );
  XOR2_X1 U420 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n367) );
  XOR2_X1 U421 ( .A(G218GAT), .B(G162GAT), .Z(n416) );
  XNOR2_X1 U422 ( .A(n416), .B(n365), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U424 ( .A(G92GAT), .B(G106GAT), .Z(n369) );
  NAND2_X1 U425 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U427 ( .A(n371), .B(n370), .Z(n373) );
  XOR2_X1 U428 ( .A(G190GAT), .B(G134GAT), .Z(n436) );
  XNOR2_X1 U429 ( .A(G36GAT), .B(n436), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n473) );
  NAND2_X1 U433 ( .A1(n378), .A2(n473), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n379), .B(KEYINPUT47), .ZN(n386) );
  XNOR2_X1 U435 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n380), .B(n473), .ZN(n586) );
  NOR2_X1 U437 ( .A1(n586), .A2(n472), .ZN(n381) );
  XNOR2_X1 U438 ( .A(KEYINPUT45), .B(n381), .ZN(n382) );
  INV_X1 U439 ( .A(n549), .ZN(n574) );
  XOR2_X1 U440 ( .A(KEYINPUT68), .B(n574), .Z(n559) );
  INV_X1 U441 ( .A(n559), .ZN(n457) );
  NAND2_X1 U442 ( .A1(n382), .A2(n457), .ZN(n384) );
  NOR2_X1 U443 ( .A1(n384), .A2(n336), .ZN(n385) );
  NOR2_X1 U444 ( .A1(n386), .A2(n385), .ZN(n389) );
  XOR2_X1 U445 ( .A(KEYINPUT64), .B(KEYINPUT114), .Z(n387) );
  NAND2_X1 U446 ( .A1(n523), .A2(n532), .ZN(n391) );
  XOR2_X1 U447 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n393) );
  XNOR2_X1 U448 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n398) );
  XNOR2_X1 U450 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n394), .B(G127GAT), .ZN(n437) );
  XOR2_X1 U452 ( .A(n437), .B(G1GAT), .Z(n396) );
  NAND2_X1 U453 ( .A1(G225GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n413) );
  XOR2_X1 U456 ( .A(KEYINPUT6), .B(G148GAT), .Z(n400) );
  XNOR2_X1 U457 ( .A(G141GAT), .B(G120GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U459 ( .A(G57GAT), .B(KEYINPUT1), .Z(n402) );
  XNOR2_X1 U460 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U462 ( .A(n404), .B(n403), .Z(n411) );
  XOR2_X1 U463 ( .A(G85GAT), .B(G162GAT), .Z(n408) );
  XOR2_X1 U464 ( .A(G155GAT), .B(KEYINPUT83), .Z(n406) );
  XNOR2_X1 U465 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n428) );
  XNOR2_X1 U467 ( .A(G29GAT), .B(n428), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U469 ( .A(G134GAT), .B(n409), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n521) );
  INV_X1 U472 ( .A(n521), .ZN(n571) );
  XOR2_X1 U473 ( .A(KEYINPUT23), .B(KEYINPUT81), .Z(n415) );
  XNOR2_X1 U474 ( .A(KEYINPUT85), .B(G204GAT), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n421) );
  XOR2_X1 U476 ( .A(KEYINPUT24), .B(n416), .Z(n419) );
  XNOR2_X1 U477 ( .A(G50GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U478 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U479 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U480 ( .A1(G228GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U482 ( .A(n424), .B(KEYINPUT22), .Z(n427) );
  XNOR2_X1 U483 ( .A(n425), .B(KEYINPUT84), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U485 ( .A(n429), .B(n428), .Z(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n464) );
  AND2_X1 U487 ( .A1(n571), .A2(n464), .ZN(n432) );
  NAND2_X1 U488 ( .A1(n290), .A2(n432), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n443) );
  XOR2_X1 U491 ( .A(G15GAT), .B(n439), .Z(n441) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U494 ( .A(n443), .B(n442), .Z(n451) );
  XOR2_X1 U495 ( .A(KEYINPUT78), .B(KEYINPUT80), .Z(n445) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G99GAT), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U498 ( .A(G176GAT), .B(KEYINPUT20), .Z(n447) );
  XNOR2_X1 U499 ( .A(G169GAT), .B(KEYINPUT79), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n451), .B(n450), .ZN(n533) );
  NOR2_X1 U503 ( .A1(n452), .A2(n533), .ZN(n568) );
  INV_X1 U504 ( .A(n473), .ZN(n556) );
  NAND2_X1 U505 ( .A1(n568), .A2(n556), .ZN(n456) );
  XOR2_X1 U506 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n454) );
  NOR2_X1 U507 ( .A1(n457), .A2(n336), .ZN(n493) );
  INV_X1 U508 ( .A(n536), .ZN(n487) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(n523), .ZN(n466) );
  NAND2_X1 U510 ( .A1(n466), .A2(n521), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n458), .B(KEYINPUT95), .ZN(n531) );
  NAND2_X1 U512 ( .A1(n487), .A2(n531), .ZN(n459) );
  XOR2_X1 U513 ( .A(KEYINPUT96), .B(n459), .Z(n460) );
  NAND2_X1 U514 ( .A1(n533), .A2(n460), .ZN(n471) );
  INV_X1 U515 ( .A(n533), .ZN(n526) );
  NAND2_X1 U516 ( .A1(n526), .A2(n523), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n461), .A2(n464), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT97), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n463), .B(KEYINPUT25), .ZN(n468) );
  NOR2_X1 U520 ( .A1(n464), .A2(n526), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT26), .ZN(n572) );
  NAND2_X1 U522 ( .A1(n466), .A2(n572), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U524 ( .A1(n469), .A2(n571), .ZN(n470) );
  NAND2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n490) );
  INV_X1 U526 ( .A(n490), .ZN(n477) );
  XOR2_X1 U527 ( .A(KEYINPUT77), .B(KEYINPUT16), .Z(n475) );
  INV_X1 U528 ( .A(n472), .ZN(n582) );
  NAND2_X1 U529 ( .A1(n582), .A2(n473), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n477), .A2(n476), .ZN(n508) );
  NAND2_X1 U532 ( .A1(n493), .A2(n508), .ZN(n486) );
  NOR2_X1 U533 ( .A1(n571), .A2(n486), .ZN(n478) );
  XOR2_X1 U534 ( .A(G1GAT), .B(n478), .Z(n479) );
  XNOR2_X1 U535 ( .A(KEYINPUT34), .B(n479), .ZN(G1324GAT) );
  INV_X1 U536 ( .A(n523), .ZN(n480) );
  NOR2_X1 U537 ( .A1(n480), .A2(n486), .ZN(n481) );
  XOR2_X1 U538 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  NOR2_X1 U539 ( .A1(n486), .A2(n533), .ZN(n485) );
  XOR2_X1 U540 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n483) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT99), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NOR2_X1 U544 ( .A1(n487), .A2(n486), .ZN(n488) );
  XOR2_X1 U545 ( .A(KEYINPUT100), .B(n488), .Z(n489) );
  XNOR2_X1 U546 ( .A(G22GAT), .B(n489), .ZN(G1327GAT) );
  NOR2_X1 U547 ( .A1(n582), .A2(n586), .ZN(n491) );
  NAND2_X1 U548 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n492), .ZN(n518) );
  NAND2_X1 U550 ( .A1(n493), .A2(n518), .ZN(n494) );
  XOR2_X1 U551 ( .A(KEYINPUT38), .B(n494), .Z(n504) );
  NAND2_X1 U552 ( .A1(n504), .A2(n521), .ZN(n498) );
  XOR2_X1 U553 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n496) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n504), .A2(n523), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(KEYINPUT104), .ZN(n503) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n501) );
  NAND2_X1 U561 ( .A1(n504), .A2(n526), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n504), .A2(n536), .ZN(n505) );
  XNOR2_X1 U565 ( .A(n505), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  XOR2_X1 U567 ( .A(n551), .B(KEYINPUT107), .Z(n565) );
  NAND2_X1 U568 ( .A1(n574), .A2(n565), .ZN(n507) );
  XOR2_X1 U569 ( .A(KEYINPUT108), .B(n507), .Z(n519) );
  NAND2_X1 U570 ( .A1(n519), .A2(n508), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n509), .B(KEYINPUT109), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n521), .A2(n515), .ZN(n510) );
  XNOR2_X1 U573 ( .A(KEYINPUT42), .B(n510), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n523), .A2(n515), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n526), .A2(n515), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(KEYINPUT110), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U581 ( .A1(n515), .A2(n536), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(KEYINPUT111), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n528), .A2(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n522), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n528), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(KEYINPUT112), .ZN(n525) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(n525), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n526), .A2(n528), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n536), .A2(n528), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(KEYINPUT44), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n546) );
  NOR2_X1 U597 ( .A1(n533), .A2(n546), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(KEYINPUT115), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n543), .A2(n559), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U603 ( .A1(n543), .A2(n565), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NAND2_X1 U605 ( .A1(n543), .A2(n582), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U609 ( .A1(n543), .A2(n556), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  INV_X1 U611 ( .A(n572), .ZN(n547) );
  NOR2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U613 ( .A(KEYINPUT117), .B(n548), .Z(n557) );
  NAND2_X1 U614 ( .A1(n557), .A2(n549), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n550), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n553) );
  NAND2_X1 U617 ( .A1(n557), .A2(n551), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n557), .A2(n582), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n568), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n563) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(n564), .Z(n567) );
  NAND2_X1 U631 ( .A1(n565), .A2(n568), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  XOR2_X1 U633 ( .A(G183GAT), .B(KEYINPUT123), .Z(n570) );
  NAND2_X1 U634 ( .A1(n568), .A2(n582), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1350GAT) );
  AND2_X1 U636 ( .A1(n290), .A2(n571), .ZN(n573) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n585) );
  NOR2_X1 U638 ( .A1(n585), .A2(n574), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n580) );
  INV_X1 U644 ( .A(n585), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n583), .A2(n336), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

