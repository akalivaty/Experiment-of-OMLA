//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT66), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT67), .Z(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G319));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G2104), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n462), .A2(new_n464), .A3(G137), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n465), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  AND2_X1   g053(.A1(new_n464), .A2(new_n465), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n462), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n469), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT70), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n469), .B2(G112), .ZN(new_n484));
  INV_X1    g059(.A(G100), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(new_n469), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT71), .Z(new_n487));
  NOR2_X1   g062(.A1(new_n480), .A2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G136), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n483), .A2(new_n489), .ZN(G162));
  AND2_X1   g065(.A1(KEYINPUT4), .A2(G138), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n462), .A2(new_n464), .A3(new_n465), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(G102), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(G2105), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n462), .A2(new_n464), .A3(G126), .A4(new_n465), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n469), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n472), .A2(new_n465), .A3(G138), .A4(new_n469), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n494), .A2(new_n497), .A3(new_n500), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G651), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n503), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT72), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G88), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n516));
  INV_X1    g091(.A(G75), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(KEYINPUT73), .A2(G75), .A3(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n506), .A2(new_n507), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n519), .B(new_n520), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n503), .A2(new_n505), .A3(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n523), .A2(G651), .B1(G50), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n515), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n503), .A2(new_n505), .A3(G543), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n514), .A2(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XOR2_X1   g108(.A(new_n533), .B(KEYINPUT7), .Z(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n530), .B2(KEYINPUT74), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n531), .A2(new_n532), .A3(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n502), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n508), .A2(new_n509), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT72), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(G90), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n524), .A2(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n541), .A2(KEYINPUT75), .A3(new_n542), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n521), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n550), .A2(G651), .B1(G43), .B2(new_n524), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n539), .A2(G81), .A3(new_n540), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT76), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  OAI21_X1  g135(.A(KEYINPUT77), .B1(new_n510), .B2(new_n513), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n539), .A2(new_n562), .A3(new_n540), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(G91), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OR3_X1    g140(.A1(new_n529), .A2(KEYINPUT9), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT9), .B1(new_n529), .B2(new_n565), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n521), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n566), .A2(new_n567), .B1(new_n570), .B2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n564), .A2(new_n571), .ZN(G299));
  AND3_X1   g147(.A1(new_n541), .A2(KEYINPUT75), .A3(new_n542), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT75), .B1(new_n541), .B2(new_n542), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n573), .A2(new_n574), .B1(new_n502), .B2(new_n537), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  NAND2_X1  g151(.A1(new_n515), .A2(new_n525), .ZN(G303));
  NAND3_X1  g152(.A1(new_n561), .A2(G87), .A3(new_n563), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n512), .A2(G74), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(G49), .B2(new_n524), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G288));
  NAND3_X1  g156(.A1(new_n561), .A2(G86), .A3(new_n563), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n521), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G48), .B2(new_n524), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G305));
  NAND3_X1  g162(.A1(new_n539), .A2(G85), .A3(new_n540), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n524), .A2(G47), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n591), .A2(new_n592), .B1(new_n502), .B2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n561), .A2(G92), .A3(new_n563), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n561), .A2(KEYINPUT10), .A3(G92), .A4(new_n563), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n521), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(KEYINPUT79), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n502), .B1(new_n603), .B2(KEYINPUT79), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n604), .A2(new_n605), .B1(G54), .B2(new_n524), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n595), .B1(new_n607), .B2(G868), .ZN(G284));
  XOR2_X1   g183(.A(G284), .B(KEYINPUT80), .Z(G321));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(G299), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n610), .B2(G168), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(new_n610), .B2(G168), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NOR2_X1   g190(.A1(new_n553), .A2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n600), .A2(new_n606), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n617), .A2(G559), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT81), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n616), .B1(new_n619), .B2(G868), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n488), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n481), .A2(G123), .ZN(new_n623));
  NOR2_X1   g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(new_n469), .B2(G111), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n629));
  NOR3_X1   g204(.A1(new_n461), .A2(new_n463), .A3(G2105), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n633), .ZN(G156));
  INV_X1    g209(.A(KEYINPUT14), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT84), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n640), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(G14), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n645), .A2(new_n648), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  INV_X1    g233(.A(new_n656), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n655), .B1(new_n659), .B2(new_n653), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n660), .A2(KEYINPUT85), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(KEYINPUT85), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n653), .B(KEYINPUT17), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n661), .B(new_n662), .C1(new_n659), .C2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(new_n655), .A3(new_n659), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n658), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n627), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2100), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT86), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n672), .B(new_n673), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  MUX2_X1   g253(.A(new_n677), .B(new_n678), .S(new_n671), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1986), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(G229));
  MUX2_X1   g261(.A(G23), .B(G288), .S(G16), .Z(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT91), .B(KEYINPUT33), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G1976), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n688), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n687), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G1976), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G303), .B2(G16), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n695), .A2(G6), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G305), .B2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT32), .B(G1981), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n701), .A2(new_n703), .ZN(new_n705));
  NOR3_X1   g280(.A1(new_n699), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n691), .A2(new_n694), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT92), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT34), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n707), .B(KEYINPUT92), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT87), .B(G29), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(G25), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n488), .A2(G131), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT88), .Z(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(new_n469), .B2(G107), .ZN(new_n719));
  INV_X1    g294(.A(G95), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n469), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n481), .B2(G119), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(new_n714), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT89), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT90), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n725), .A2(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n695), .A2(G24), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n593), .A2(new_n502), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n588), .A2(new_n590), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(KEYINPUT78), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(new_n695), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1986), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n729), .A2(new_n730), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n711), .A2(new_n713), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(KEYINPUT36), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n711), .A2(new_n713), .A3(new_n742), .A4(new_n739), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT31), .B(G11), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(G28), .ZN(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n746), .B2(G28), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n745), .B1(new_n747), .B2(new_n749), .C1(new_n626), .C2(new_n714), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT99), .Z(new_n751));
  INV_X1    g326(.A(G1961), .ZN(new_n752));
  NOR2_X1   g327(.A1(G171), .A2(new_n695), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G5), .B2(new_n695), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(G168), .A2(G16), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT97), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G16), .B2(G21), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n755), .B1(new_n760), .B2(G1966), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n760), .A2(KEYINPUT100), .A3(G1966), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT100), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n758), .B(KEYINPUT98), .ZN(new_n764));
  INV_X1    g339(.A(G1966), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n761), .B1(new_n762), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n767), .A2(KEYINPUT101), .ZN(new_n768));
  NAND2_X1  g343(.A1(G162), .A2(new_n715), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n715), .A2(G35), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT29), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(KEYINPUT29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G2090), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n772), .A2(G2090), .A3(new_n773), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n714), .A2(G26), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT28), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n488), .A2(G140), .ZN(new_n780));
  OR2_X1    g355(.A1(G104), .A2(G2105), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n781), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n782));
  INV_X1    g357(.A(G128), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n479), .A2(new_n462), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n780), .B(new_n782), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n779), .B1(new_n787), .B2(new_n748), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT94), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2067), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n695), .A2(G4), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n607), .B2(new_n695), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT93), .B(G1348), .Z(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n776), .A2(new_n777), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n695), .A2(G19), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n554), .B2(new_n695), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(G1341), .Z(new_n798));
  INV_X1    g373(.A(G2084), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT24), .B(G34), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n714), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT96), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n477), .B2(new_n748), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n798), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n799), .B2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n748), .A2(G32), .ZN(new_n806));
  NAND3_X1  g381(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT26), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n469), .A2(G105), .A3(G2104), .ZN(new_n810));
  INV_X1    g385(.A(G129), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n809), .B(new_n810), .C1(new_n785), .C2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G141), .B2(new_n488), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n806), .B1(new_n813), .B2(new_n748), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT27), .B(G1996), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G2072), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n748), .A2(G33), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n488), .A2(G139), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT25), .Z(new_n821));
  AND2_X1   g396(.A1(new_n472), .A2(new_n465), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n822), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n819), .B(new_n821), .C1(new_n469), .C2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT95), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n818), .B1(new_n825), .B2(G29), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n816), .B1(new_n817), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n695), .A2(G20), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT23), .Z(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G299), .B2(G16), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1956), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n754), .A2(new_n752), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n805), .A2(new_n827), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n826), .A2(new_n817), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n792), .A2(new_n793), .ZN(new_n835));
  NAND2_X1  g410(.A1(G164), .A2(new_n715), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G27), .B2(new_n715), .ZN(new_n837));
  INV_X1    g412(.A(G2078), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n834), .A2(new_n835), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n795), .A2(new_n833), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n767), .B2(KEYINPUT101), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n768), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n744), .A2(new_n844), .ZN(G311));
  NAND2_X1  g420(.A1(new_n744), .A2(new_n844), .ZN(G150));
  OAI21_X1  g421(.A(G67), .B1(new_n506), .B2(new_n507), .ZN(new_n847));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n849), .A2(G651), .B1(new_n524), .B2(G55), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n539), .A2(G93), .A3(new_n540), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NOR2_X1   g429(.A1(new_n617), .A2(new_n614), .ZN(new_n855));
  AND4_X1   g430(.A1(new_n552), .A2(new_n551), .A3(new_n851), .A4(new_n850), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n552), .A2(new_n551), .B1(new_n850), .B2(new_n851), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n855), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT103), .ZN(new_n860));
  XNOR2_X1  g435(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  INV_X1    g438(.A(G860), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n862), .B2(KEYINPUT39), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n854), .B1(new_n863), .B2(new_n865), .ZN(G145));
  NAND2_X1  g441(.A1(new_n488), .A2(G142), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n481), .A2(G130), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n869), .A2(new_n469), .A3(G118), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n469), .B2(G118), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n867), .B(new_n868), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n723), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n631), .ZN(new_n875));
  INV_X1    g450(.A(new_n494), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n495), .A2(new_n496), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G2105), .ZN(new_n878));
  INV_X1    g453(.A(new_n500), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n786), .B(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n813), .ZN(new_n882));
  INV_X1    g457(.A(new_n825), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n821), .B1(new_n823), .B2(new_n469), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(G139), .B2(new_n488), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n886), .B2(new_n882), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n875), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n626), .B(G160), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G162), .ZN(new_n890));
  AOI21_X1  g465(.A(G37), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n890), .B2(new_n888), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n582), .A2(new_n586), .B1(new_n515), .B2(new_n525), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(G166), .A2(new_n582), .A3(new_n586), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT106), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(G305), .A2(G303), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT106), .B1(new_n900), .B2(new_n895), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n578), .A2(KEYINPUT105), .A3(new_n580), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT105), .B1(new_n578), .B2(new_n580), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n903), .A2(new_n736), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n906));
  NAND2_X1  g481(.A1(G288), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G290), .B1(new_n907), .B2(new_n902), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n899), .B(new_n901), .C1(new_n905), .C2(new_n908), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n900), .A2(KEYINPUT106), .A3(new_n895), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n736), .B1(new_n903), .B2(new_n904), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n907), .A2(G290), .A3(new_n902), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n894), .B1(new_n914), .B2(KEYINPUT42), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(KEYINPUT42), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n915), .B(new_n916), .Z(new_n917));
  AND2_X1   g492(.A1(new_n619), .A2(new_n858), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n619), .A2(new_n858), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G299), .B1(new_n600), .B2(new_n606), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n600), .A2(G299), .A3(new_n606), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(KEYINPUT41), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT41), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n600), .A2(G299), .A3(new_n606), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n921), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n920), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n922), .A2(new_n923), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n918), .B2(new_n919), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n929), .A2(new_n934), .A3(new_n931), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n917), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n935), .A2(new_n917), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n852), .A2(new_n610), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(G295));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n939), .ZN(G331));
  NAND2_X1  g516(.A1(new_n553), .A2(new_n852), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n551), .A2(new_n850), .A3(new_n552), .A4(new_n851), .ZN(new_n943));
  NAND3_X1  g518(.A1(G301), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NAND2_X1  g520(.A1(G171), .A2(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n944), .A2(new_n946), .A3(G168), .ZN(new_n947));
  AOI21_X1  g522(.A(G168), .B1(new_n944), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT41), .B1(new_n922), .B2(new_n923), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n926), .A2(new_n921), .A3(new_n925), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n858), .A2(G301), .ZN(new_n953));
  NOR2_X1   g528(.A1(G171), .A2(new_n945), .ZN(new_n954));
  OAI21_X1  g529(.A(G286), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n944), .A2(new_n946), .A3(G168), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n955), .A2(new_n956), .B1(new_n922), .B2(new_n923), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n952), .A2(new_n914), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G37), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n928), .B2(new_n949), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(new_n961), .B2(new_n914), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n962), .B2(KEYINPUT110), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n966), .B(new_n960), .C1(new_n961), .C2(new_n914), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n964), .B1(new_n962), .B2(new_n959), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n914), .B1(new_n952), .B2(new_n958), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT110), .B1(new_n972), .B2(G37), .ZN(new_n973));
  INV_X1    g548(.A(new_n959), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n973), .A2(new_n964), .A3(new_n974), .A4(new_n967), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT111), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n963), .A2(new_n977), .A3(new_n964), .A4(new_n967), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n962), .B2(new_n959), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT44), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT112), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n984), .B(new_n981), .C1(new_n976), .C2(new_n978), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n971), .B1(new_n983), .B2(new_n985), .ZN(G397));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(G164), .B2(G1384), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n470), .A2(G40), .A3(new_n476), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n813), .B(G1996), .ZN(new_n992));
  INV_X1    g567(.A(G2067), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n786), .B(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n995), .A2(new_n728), .A3(new_n718), .A4(new_n722), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n787), .A2(new_n993), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n991), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n991), .A2(G1986), .A3(G290), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(KEYINPUT48), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n723), .B(new_n728), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1000), .B1(new_n1002), .B2(new_n990), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(KEYINPUT48), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n998), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1996), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n990), .A2(KEYINPUT46), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n991), .B2(G1996), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n994), .A2(new_n813), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1007), .B(new_n1009), .C1(new_n1010), .C2(new_n991), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1005), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT127), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT126), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  INV_X1    g593(.A(G1384), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n880), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT117), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n497), .A2(new_n500), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1384), .B1(new_n1022), .B2(new_n876), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n1018), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1021), .A2(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n470), .A2(G40), .A3(new_n476), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(KEYINPUT116), .A3(new_n1027), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1026), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1956), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n987), .A2(G1384), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n989), .B1(new_n880), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT56), .B(G2072), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n988), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n1041));
  XNOR2_X1  g616(.A(G299), .B(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1031), .A2(new_n1027), .A3(new_n1020), .ZN(new_n1046));
  INV_X1    g621(.A(G1348), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1023), .A2(new_n993), .A3(new_n1027), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1045), .B1(new_n617), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1035), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1035), .A2(KEYINPUT118), .A3(new_n1039), .A4(new_n1042), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1052), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT120), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n988), .A2(new_n1037), .A3(new_n1006), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT58), .B(G1341), .Z(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n554), .ZN(new_n1068));
  NOR2_X1   g643(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1062), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n553), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1072), .A2(KEYINPUT121), .A3(new_n1069), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1061), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1068), .A2(new_n1062), .A3(new_n1070), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT121), .B1(new_n1072), .B2(new_n1069), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1075), .B(new_n1076), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1050), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n607), .B1(new_n1050), .B2(new_n1078), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1048), .A2(KEYINPUT60), .A3(new_n617), .A4(new_n1049), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1074), .A2(new_n1077), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1053), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1035), .A2(KEYINPUT122), .A3(new_n1039), .A4(new_n1042), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1085), .A2(new_n1045), .A3(KEYINPUT61), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1042), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1040), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT61), .B1(new_n1057), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1058), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1036), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1027), .B1(G164), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT45), .B1(new_n880), .B2(new_n1019), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n765), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1031), .A2(new_n1020), .A3(new_n799), .A4(new_n1027), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n1097), .A3(G168), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G8), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT51), .ZN(new_n1100));
  AOI21_X1  g675(.A(G168), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n1102));
  OAI211_X1 g677(.A(G8), .B(new_n1098), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1100), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1046), .A2(new_n752), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n988), .A2(new_n1037), .A3(new_n838), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1094), .A2(new_n1095), .A3(G2078), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n1114), .B2(KEYINPUT53), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(KEYINPUT124), .A3(new_n1110), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1112), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(G171), .A2(KEYINPUT125), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1108), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1114), .A2(KEYINPUT53), .B1(new_n752), .B2(new_n1046), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1116), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT124), .B1(new_n1111), .B2(new_n1110), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1121), .B(G301), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(G301), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1108), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n586), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT115), .B(G86), .Z(new_n1132));
  NOR3_X1   g707(.A1(new_n510), .A2(new_n513), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(G1981), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(G305), .B2(G1981), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT49), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(G8), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1138), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT49), .B(new_n1134), .C1(G305), .C2(G1981), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT114), .B(G1976), .Z(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT52), .B1(G288), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n578), .A2(G1976), .A3(new_n580), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n1139), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT52), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1141), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(G303), .A2(G8), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1149), .B(KEYINPUT55), .Z(new_n1150));
  NAND2_X1  g725(.A1(new_n988), .A2(new_n1037), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1151), .A2(KEYINPUT113), .A3(new_n698), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1031), .A2(new_n1020), .A3(new_n775), .A4(new_n1027), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT113), .B1(new_n1151), .B2(new_n698), .ZN(new_n1155));
  OAI211_X1 g730(.A(G8), .B(new_n1150), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1026), .A2(new_n1030), .A3(new_n775), .A4(new_n1032), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1151), .A2(new_n698), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1138), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1148), .B(new_n1156), .C1(new_n1150), .C2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1107), .A2(new_n1124), .A3(new_n1130), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1092), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1148), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1139), .ZN(new_n1166));
  NOR2_X1   g741(.A1(G305), .A2(G1981), .ZN(new_n1167));
  NOR2_X1   g742(.A1(G288), .A2(G1976), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1167), .B1(new_n1141), .B2(new_n1168), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n1165), .A2(new_n1156), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1172), .A2(G8), .A3(G168), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1171), .B1(new_n1160), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(G8), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1150), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1173), .A2(new_n1171), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1177), .A2(new_n1156), .A3(new_n1148), .A4(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1170), .B1(new_n1174), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(KEYINPUT123), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1100), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1184), .A2(KEYINPUT62), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1129), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1160), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1182), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1180), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1164), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(G290), .B(G1986), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n990), .B1(new_n1002), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1017), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  AOI22_X1  g769(.A1(new_n1055), .A2(new_n1056), .B1(new_n1040), .B2(new_n1089), .ZN(new_n1195));
  OAI211_X1 g770(.A(new_n1083), .B(new_n1087), .C1(new_n1195), .C2(KEYINPUT61), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1162), .B1(new_n1196), .B2(new_n1058), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1180), .A2(new_n1189), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1017), .B(new_n1193), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1016), .B1(new_n1194), .B2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g776(.A(new_n458), .B1(new_n650), .B2(new_n651), .ZN(new_n1203));
  NOR3_X1   g777(.A1(G229), .A2(G227), .A3(new_n1203), .ZN(new_n1204));
  NAND4_X1  g778(.A1(new_n1204), .A2(new_n892), .A3(new_n969), .A4(new_n968), .ZN(G225));
  INV_X1    g779(.A(G225), .ZN(G308));
endmodule


