

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737;

  INV_X1 U370 ( .A(G953), .ZN(n457) );
  XNOR2_X2 U371 ( .A(n409), .B(G469), .ZN(n535) );
  NOR2_X1 U372 ( .A1(n675), .A2(n734), .ZN(n596) );
  INV_X1 U373 ( .A(G125), .ZN(n425) );
  AND2_X1 U374 ( .A1(n387), .A2(n391), .ZN(n386) );
  NAND2_X1 U375 ( .A1(n572), .A2(n571), .ZN(n366) );
  XNOR2_X1 U376 ( .A(n596), .B(KEYINPUT81), .ZN(n603) );
  AND2_X1 U377 ( .A1(n595), .A2(n353), .ZN(n675) );
  NOR2_X1 U378 ( .A1(n429), .A2(n434), .ZN(n401) );
  NAND2_X1 U379 ( .A1(n433), .A2(n432), .ZN(n430) );
  NAND2_X1 U380 ( .A1(n435), .A2(n358), .ZN(n434) );
  AND2_X1 U381 ( .A1(n615), .A2(n582), .ZN(n583) );
  XNOR2_X1 U382 ( .A(n663), .B(n664), .ZN(n665) );
  XNOR2_X1 U383 ( .A(n427), .B(n426), .ZN(n623) );
  XNOR2_X1 U384 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U385 ( .A(n379), .B(n714), .ZN(n693) );
  XNOR2_X1 U386 ( .A(n378), .B(n377), .ZN(n714) );
  XNOR2_X1 U387 ( .A(n473), .B(n490), .ZN(n378) );
  XNOR2_X1 U388 ( .A(n381), .B(n380), .ZN(n379) );
  XNOR2_X1 U389 ( .A(n351), .B(n382), .ZN(n381) );
  XNOR2_X1 U390 ( .A(n472), .B(n471), .ZN(n490) );
  XOR2_X1 U391 ( .A(n474), .B(n475), .Z(n351) );
  XNOR2_X1 U392 ( .A(n462), .B(n464), .ZN(n380) );
  NAND2_X1 U393 ( .A1(n470), .A2(n469), .ZN(n472) );
  XNOR2_X1 U394 ( .A(n465), .B(n428), .ZN(n377) );
  XNOR2_X1 U395 ( .A(n425), .B(G146), .ZN(n463) );
  XNOR2_X1 U396 ( .A(n413), .B(G143), .ZN(n474) );
  XNOR2_X1 U397 ( .A(n452), .B(G122), .ZN(n465) );
  INV_X1 U398 ( .A(G128), .ZN(n413) );
  XOR2_X1 U399 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n475) );
  XNOR2_X1 U400 ( .A(G116), .B(G107), .ZN(n452) );
  XNOR2_X1 U401 ( .A(G119), .B(G113), .ZN(n471) );
  XNOR2_X1 U402 ( .A(G110), .B(G104), .ZN(n466) );
  BUF_X1 U403 ( .A(n597), .Z(n347) );
  INV_X1 U404 ( .A(n433), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n392), .B(n359), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n401), .B(n581), .ZN(n597) );
  XNOR2_X1 U407 ( .A(n479), .B(n478), .ZN(n541) );
  OR2_X2 U408 ( .A1(n651), .A2(KEYINPUT79), .ZN(n356) );
  XNOR2_X1 U409 ( .A(n392), .B(n359), .ZN(n717) );
  OR2_X1 U410 ( .A1(n626), .A2(n613), .ZN(n400) );
  NOR2_X1 U411 ( .A1(n623), .A2(n622), .ZN(n628) );
  OR2_X1 U412 ( .A1(n700), .A2(G902), .ZN(n409) );
  NOR2_X1 U413 ( .A1(n552), .A2(n680), .ZN(n422) );
  XNOR2_X1 U414 ( .A(n406), .B(n404), .ZN(n622) );
  XNOR2_X1 U415 ( .A(n405), .B(KEYINPUT95), .ZN(n404) );
  NAND2_X1 U416 ( .A1(n512), .A2(G221), .ZN(n406) );
  INV_X1 U417 ( .A(KEYINPUT21), .ZN(n405) );
  XNOR2_X1 U418 ( .A(n410), .B(KEYINPUT103), .ZN(n384) );
  XNOR2_X1 U419 ( .A(n412), .B(KEYINPUT98), .ZN(n411) );
  NAND2_X1 U420 ( .A1(n390), .A2(n669), .ZN(n385) );
  NOR2_X1 U421 ( .A1(n733), .A2(KEYINPUT44), .ZN(n388) );
  XNOR2_X1 U422 ( .A(n474), .B(n455), .ZN(n486) );
  INV_X1 U423 ( .A(G134), .ZN(n455) );
  XNOR2_X1 U424 ( .A(n486), .B(n373), .ZN(n414) );
  XNOR2_X1 U425 ( .A(n487), .B(n374), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n375), .B(G137), .ZN(n374) );
  INV_X1 U427 ( .A(KEYINPUT4), .ZN(n375) );
  XOR2_X1 U428 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n503) );
  XNOR2_X1 U429 ( .A(n463), .B(n424), .ZN(n722) );
  XNOR2_X1 U430 ( .A(KEYINPUT10), .B(G140), .ZN(n424) );
  XNOR2_X1 U431 ( .A(n454), .B(KEYINPUT100), .ZN(n438) );
  XOR2_X1 U432 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n454) );
  XOR2_X1 U433 ( .A(G140), .B(G107), .Z(n514) );
  XNOR2_X1 U434 ( .A(n414), .B(G146), .ZN(n519) );
  NAND2_X1 U435 ( .A1(n352), .A2(n367), .ZN(n569) );
  NAND2_X1 U436 ( .A1(n369), .A2(n368), .ZN(n367) );
  NAND2_X1 U437 ( .A1(n612), .A2(KEYINPUT39), .ZN(n370) );
  NOR2_X1 U438 ( .A1(n347), .A2(n619), .ZN(n601) );
  NOR2_X1 U439 ( .A1(n531), .A2(n497), .ZN(n524) );
  XNOR2_X1 U440 ( .A(n400), .B(KEYINPUT30), .ZN(n497) );
  XNOR2_X1 U441 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U442 ( .A1(n407), .A2(n536), .ZN(n545) );
  XNOR2_X1 U443 ( .A(n534), .B(n408), .ZN(n407) );
  XNOR2_X1 U444 ( .A(KEYINPUT111), .B(KEYINPUT28), .ZN(n408) );
  XNOR2_X1 U445 ( .A(n511), .B(n510), .ZN(n426) );
  OR2_X1 U446 ( .A1(n710), .A2(G902), .ZN(n427) );
  AND2_X2 U447 ( .A1(n415), .A2(n416), .ZN(n708) );
  XNOR2_X1 U448 ( .A(n695), .B(n694), .ZN(n697) );
  XNOR2_X1 U449 ( .A(n376), .B(G131), .ZN(n487) );
  INV_X1 U450 ( .A(KEYINPUT68), .ZN(n376) );
  NAND2_X1 U451 ( .A1(G237), .A2(G234), .ZN(n480) );
  OR2_X1 U452 ( .A1(G902), .A2(G237), .ZN(n495) );
  XNOR2_X1 U453 ( .A(n499), .B(n500), .ZN(n512) );
  XOR2_X1 U454 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n500) );
  NOR2_X1 U455 ( .A1(G953), .A2(G237), .ZN(n488) );
  XNOR2_X1 U456 ( .A(G113), .B(G143), .ZN(n441) );
  XNOR2_X1 U457 ( .A(n463), .B(n461), .ZN(n382) );
  XNOR2_X1 U458 ( .A(KEYINPUT4), .B(KEYINPUT86), .ZN(n461) );
  INV_X1 U459 ( .A(KEYINPUT79), .ZN(n364) );
  INV_X1 U460 ( .A(n528), .ZN(n369) );
  NAND2_X1 U461 ( .A1(n554), .A2(n555), .ZN(n562) );
  INV_X1 U462 ( .A(n622), .ZN(n582) );
  NOR2_X1 U463 ( .A1(n529), .A2(n539), .ZN(n615) );
  AND2_X1 U464 ( .A1(n627), .A2(n628), .ZN(n605) );
  INV_X1 U465 ( .A(KEYINPUT108), .ZN(n522) );
  NAND2_X1 U466 ( .A1(n386), .A2(n383), .ZN(n392) );
  NOR2_X1 U467 ( .A1(n385), .A2(n384), .ZN(n383) );
  INV_X1 U468 ( .A(KEYINPUT72), .ZN(n363) );
  XNOR2_X1 U469 ( .A(n562), .B(n393), .ZN(n556) );
  INV_X1 U470 ( .A(KEYINPUT113), .ZN(n393) );
  INV_X1 U471 ( .A(n623), .ZN(n594) );
  XNOR2_X1 U472 ( .A(n494), .B(n440), .ZN(n626) );
  NOR2_X1 U473 ( .A1(n663), .A2(G902), .ZN(n494) );
  XNOR2_X1 U474 ( .A(n521), .B(KEYINPUT96), .ZN(n607) );
  XNOR2_X1 U475 ( .A(n626), .B(KEYINPUT6), .ZN(n598) );
  INV_X1 U476 ( .A(n726), .ZN(n365) );
  INV_X1 U477 ( .A(KEYINPUT16), .ZN(n428) );
  XNOR2_X1 U478 ( .A(n507), .B(n506), .ZN(n509) );
  XNOR2_X1 U479 ( .A(n439), .B(n437), .ZN(n704) );
  XNOR2_X1 U480 ( .A(n456), .B(n453), .ZN(n439) );
  XNOR2_X1 U481 ( .A(n459), .B(n438), .ZN(n437) );
  XNOR2_X1 U482 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U483 ( .A(n519), .B(n520), .ZN(n700) );
  XNOR2_X1 U484 ( .A(KEYINPUT42), .B(n537), .ZN(n737) );
  XNOR2_X1 U485 ( .A(n372), .B(n360), .ZN(n732) );
  XNOR2_X1 U486 ( .A(n417), .B(KEYINPUT35), .ZN(n733) );
  INV_X1 U487 ( .A(n602), .ZN(n418) );
  XNOR2_X1 U488 ( .A(n590), .B(KEYINPUT76), .ZN(n591) );
  NOR2_X1 U489 ( .A1(n539), .A2(n540), .ZN(n681) );
  NOR2_X1 U490 ( .A1(n545), .A2(n580), .ZN(n682) );
  INV_X1 U491 ( .A(n434), .ZN(n431) );
  INV_X1 U492 ( .A(KEYINPUT56), .ZN(n402) );
  OR2_X1 U493 ( .A1(KEYINPUT2), .A2(n573), .ZN(n350) );
  AND2_X1 U494 ( .A1(n371), .A2(n370), .ZN(n352) );
  NOR2_X1 U495 ( .A1(n594), .A2(n604), .ZN(n353) );
  OR2_X1 U496 ( .A1(n681), .A2(n676), .ZN(n354) );
  XOR2_X1 U497 ( .A(n579), .B(KEYINPUT92), .Z(n355) );
  INV_X1 U498 ( .A(n613), .ZN(n436) );
  XOR2_X1 U499 ( .A(n492), .B(n491), .Z(n357) );
  OR2_X1 U500 ( .A1(n436), .A2(n543), .ZN(n358) );
  XNOR2_X1 U501 ( .A(n592), .B(n591), .ZN(n734) );
  XNOR2_X1 U502 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n359) );
  XNOR2_X1 U503 ( .A(n519), .B(n357), .ZN(n663) );
  XOR2_X1 U504 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n360) );
  XNOR2_X1 U505 ( .A(G902), .B(KEYINPUT15), .ZN(n498) );
  XOR2_X1 U506 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n361) );
  NAND2_X1 U507 ( .A1(n717), .A2(n362), .ZN(n609) );
  INV_X1 U508 ( .A(n366), .ZN(n362) );
  XNOR2_X1 U509 ( .A(n366), .B(n363), .ZN(n650) );
  XNOR2_X1 U510 ( .A(n366), .B(n364), .ZN(n573) );
  XNOR2_X1 U511 ( .A(n366), .B(n365), .ZN(n723) );
  NOR2_X1 U512 ( .A1(n612), .A2(KEYINPUT39), .ZN(n368) );
  NAND2_X1 U513 ( .A1(n528), .A2(KEYINPUT39), .ZN(n371) );
  NAND2_X1 U514 ( .A1(n569), .A2(n681), .ZN(n372) );
  NAND2_X1 U515 ( .A1(n389), .A2(n388), .ZN(n387) );
  INV_X1 U516 ( .A(n603), .ZN(n389) );
  NAND2_X1 U517 ( .A1(n733), .A2(KEYINPUT44), .ZN(n390) );
  NAND2_X1 U518 ( .A1(n603), .A2(KEYINPUT44), .ZN(n391) );
  NAND2_X1 U519 ( .A1(n422), .A2(n689), .ZN(n421) );
  NOR2_X1 U520 ( .A1(n349), .A2(KEYINPUT2), .ZN(n653) );
  NAND2_X1 U521 ( .A1(n647), .A2(n646), .ZN(n398) );
  NAND2_X1 U522 ( .A1(n394), .A2(n698), .ZN(n403) );
  XNOR2_X1 U523 ( .A(n696), .B(n697), .ZN(n394) );
  NAND2_X1 U524 ( .A1(n652), .A2(n651), .ZN(n415) );
  NAND2_X1 U525 ( .A1(n708), .A2(G210), .ZN(n696) );
  XNOR2_X1 U526 ( .A(n538), .B(KEYINPUT46), .ZN(n423) );
  NAND2_X1 U527 ( .A1(n693), .A2(n498), .ZN(n479) );
  NAND2_X1 U528 ( .A1(n396), .A2(n395), .ZN(n647) );
  INV_X1 U529 ( .A(n653), .ZN(n395) );
  NAND2_X1 U530 ( .A1(n356), .A2(n350), .ZN(n396) );
  XNOR2_X1 U531 ( .A(n397), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U532 ( .A1(n667), .A2(n698), .ZN(n397) );
  NOR2_X1 U533 ( .A1(n653), .A2(n498), .ZN(n416) );
  XNOR2_X1 U534 ( .A(n398), .B(KEYINPUT121), .ZN(n648) );
  NOR2_X1 U535 ( .A1(n553), .A2(n421), .ZN(n420) );
  NOR2_X1 U536 ( .A1(n528), .A2(n348), .ZN(n525) );
  NAND2_X1 U537 ( .A1(n523), .A2(n524), .ZN(n528) );
  NAND2_X1 U538 ( .A1(n541), .A2(n544), .ZN(n435) );
  NAND2_X1 U539 ( .A1(n423), .A2(n420), .ZN(n561) );
  XNOR2_X1 U540 ( .A(n399), .B(n361), .ZN(G75) );
  NAND2_X1 U541 ( .A1(n648), .A2(n457), .ZN(n399) );
  XNOR2_X1 U542 ( .A(n403), .B(n402), .ZN(G51) );
  XNOR2_X2 U543 ( .A(n535), .B(KEYINPUT1), .ZN(n627) );
  NAND2_X1 U544 ( .A1(n411), .A2(n354), .ZN(n410) );
  NAND2_X1 U545 ( .A1(n686), .A2(n671), .ZN(n412) );
  XNOR2_X1 U546 ( .A(n414), .B(n722), .ZN(n726) );
  NAND2_X1 U547 ( .A1(n535), .A2(n628), .ZN(n521) );
  NAND2_X1 U548 ( .A1(n419), .A2(n418), .ZN(n417) );
  XNOR2_X1 U549 ( .A(n601), .B(KEYINPUT34), .ZN(n419) );
  NAND2_X1 U550 ( .A1(n430), .A2(n355), .ZN(n429) );
  NAND2_X1 U551 ( .A1(n431), .A2(n430), .ZN(n580) );
  NAND2_X1 U552 ( .A1(n433), .A2(n436), .ZN(n557) );
  NOR2_X1 U553 ( .A1(n613), .A2(n544), .ZN(n432) );
  INV_X1 U554 ( .A(n541), .ZN(n433) );
  XNOR2_X1 U555 ( .A(n504), .B(n503), .ZN(n507) );
  INV_X1 U556 ( .A(n516), .ZN(n473) );
  XOR2_X1 U557 ( .A(n493), .B(KEYINPUT97), .Z(n440) );
  INV_X1 U558 ( .A(n692), .ZN(n570) );
  XNOR2_X1 U559 ( .A(n490), .B(n489), .ZN(n492) );
  NOR2_X1 U560 ( .A1(n735), .A2(n570), .ZN(n571) );
  XNOR2_X1 U561 ( .A(KEYINPUT83), .B(KEYINPUT33), .ZN(n599) );
  XNOR2_X1 U562 ( .A(n600), .B(n599), .ZN(n619) );
  INV_X1 U563 ( .A(n543), .ZN(n544) );
  XNOR2_X1 U564 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U565 ( .A(n658), .B(n657), .ZN(n660) );
  XNOR2_X1 U566 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U567 ( .A(KEYINPUT13), .B(G475), .ZN(n451) );
  XOR2_X1 U568 ( .A(KEYINPUT11), .B(G122), .Z(n442) );
  XNOR2_X1 U569 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U570 ( .A(n722), .B(n443), .ZN(n449) );
  XNOR2_X1 U571 ( .A(n487), .B(G104), .ZN(n447) );
  XOR2_X1 U572 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n445) );
  NAND2_X1 U573 ( .A1(G214), .A2(n488), .ZN(n444) );
  XNOR2_X1 U574 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U575 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U576 ( .A(n449), .B(n448), .ZN(n654) );
  NOR2_X1 U577 ( .A1(G902), .A2(n654), .ZN(n450) );
  XNOR2_X1 U578 ( .A(n451), .B(n450), .ZN(n529) );
  XNOR2_X1 U579 ( .A(n465), .B(KEYINPUT102), .ZN(n453) );
  XNOR2_X1 U580 ( .A(n486), .B(KEYINPUT7), .ZN(n456) );
  NAND2_X1 U581 ( .A1(G234), .A2(n457), .ZN(n458) );
  XOR2_X1 U582 ( .A(KEYINPUT8), .B(n458), .Z(n505) );
  NAND2_X1 U583 ( .A1(n505), .A2(G217), .ZN(n459) );
  NOR2_X1 U584 ( .A1(G902), .A2(n704), .ZN(n460) );
  XOR2_X1 U585 ( .A(G478), .B(n460), .Z(n539) );
  NAND2_X1 U586 ( .A1(n529), .A2(n539), .ZN(n602) );
  XOR2_X1 U587 ( .A(KEYINPUT87), .B(KEYINPUT75), .Z(n462) );
  NAND2_X1 U588 ( .A1(G224), .A2(n457), .ZN(n464) );
  XNOR2_X1 U589 ( .A(n466), .B(KEYINPUT85), .ZN(n516) );
  INV_X1 U590 ( .A(KEYINPUT3), .ZN(n467) );
  NAND2_X1 U591 ( .A1(G101), .A2(n467), .ZN(n470) );
  INV_X1 U592 ( .A(G101), .ZN(n468) );
  NAND2_X1 U593 ( .A1(n468), .A2(KEYINPUT3), .ZN(n469) );
  XOR2_X1 U594 ( .A(KEYINPUT88), .B(KEYINPUT77), .Z(n477) );
  NAND2_X1 U595 ( .A1(G210), .A2(n495), .ZN(n476) );
  XNOR2_X1 U596 ( .A(n480), .B(KEYINPUT90), .ZN(n481) );
  XNOR2_X1 U597 ( .A(KEYINPUT14), .B(n481), .ZN(n482) );
  NAND2_X1 U598 ( .A1(G952), .A2(n482), .ZN(n641) );
  NOR2_X1 U599 ( .A1(G953), .A2(n641), .ZN(n578) );
  NAND2_X1 U600 ( .A1(n482), .A2(G902), .ZN(n574) );
  NOR2_X1 U601 ( .A1(G900), .A2(n574), .ZN(n483) );
  NAND2_X1 U602 ( .A1(G953), .A2(n483), .ZN(n484) );
  XNOR2_X1 U603 ( .A(KEYINPUT105), .B(n484), .ZN(n485) );
  NOR2_X1 U604 ( .A1(n578), .A2(n485), .ZN(n531) );
  NAND2_X1 U605 ( .A1(G210), .A2(n488), .ZN(n489) );
  XNOR2_X1 U606 ( .A(G116), .B(KEYINPUT5), .ZN(n491) );
  XNOR2_X1 U607 ( .A(G472), .B(KEYINPUT70), .ZN(n493) );
  NAND2_X1 U608 ( .A1(n495), .A2(G214), .ZN(n496) );
  XNOR2_X1 U609 ( .A(n496), .B(KEYINPUT89), .ZN(n613) );
  NAND2_X1 U610 ( .A1(G234), .A2(n498), .ZN(n499) );
  NAND2_X1 U611 ( .A1(n512), .A2(G217), .ZN(n511) );
  XOR2_X1 U612 ( .A(G110), .B(G119), .Z(n502) );
  XNOR2_X1 U613 ( .A(G137), .B(G128), .ZN(n501) );
  XNOR2_X1 U614 ( .A(n502), .B(n501), .ZN(n504) );
  NAND2_X1 U615 ( .A1(G221), .A2(n505), .ZN(n506) );
  INV_X1 U616 ( .A(n722), .ZN(n508) );
  XNOR2_X1 U617 ( .A(n509), .B(n508), .ZN(n710) );
  XNOR2_X1 U618 ( .A(KEYINPUT94), .B(KEYINPUT25), .ZN(n510) );
  NAND2_X1 U619 ( .A1(G227), .A2(n457), .ZN(n513) );
  XNOR2_X1 U620 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U621 ( .A(n515), .B(KEYINPUT74), .Z(n518) );
  XNOR2_X1 U622 ( .A(n516), .B(G101), .ZN(n517) );
  XNOR2_X1 U623 ( .A(n518), .B(n517), .ZN(n520) );
  XNOR2_X1 U624 ( .A(n607), .B(n522), .ZN(n523) );
  XNOR2_X1 U625 ( .A(n525), .B(KEYINPUT109), .ZN(n526) );
  NOR2_X1 U626 ( .A1(n602), .A2(n526), .ZN(n680) );
  XNOR2_X1 U627 ( .A(KEYINPUT38), .B(KEYINPUT71), .ZN(n527) );
  XNOR2_X1 U628 ( .A(n348), .B(n527), .ZN(n612) );
  INV_X1 U629 ( .A(n529), .ZN(n540) );
  NOR2_X1 U630 ( .A1(n613), .A2(n612), .ZN(n610) );
  NAND2_X1 U631 ( .A1(n610), .A2(n615), .ZN(n530) );
  XOR2_X1 U632 ( .A(KEYINPUT41), .B(n530), .Z(n635) );
  INV_X1 U633 ( .A(n626), .ZN(n604) );
  NOR2_X1 U634 ( .A1(n622), .A2(n531), .ZN(n532) );
  XNOR2_X1 U635 ( .A(n532), .B(KEYINPUT69), .ZN(n533) );
  NOR2_X1 U636 ( .A1(n594), .A2(n533), .ZN(n555) );
  NAND2_X1 U637 ( .A1(n604), .A2(n555), .ZN(n534) );
  XNOR2_X1 U638 ( .A(n535), .B(KEYINPUT110), .ZN(n536) );
  NOR2_X1 U639 ( .A1(n635), .A2(n545), .ZN(n537) );
  NOR2_X1 U640 ( .A1(n732), .A2(n737), .ZN(n538) );
  NAND2_X1 U641 ( .A1(n540), .A2(n539), .ZN(n687) );
  INV_X1 U642 ( .A(n687), .ZN(n676) );
  XNOR2_X1 U643 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n542) );
  XNOR2_X1 U644 ( .A(n542), .B(KEYINPUT73), .ZN(n543) );
  NAND2_X1 U645 ( .A1(n354), .A2(n682), .ZN(n546) );
  XNOR2_X1 U646 ( .A(n546), .B(KEYINPUT47), .ZN(n547) );
  NAND2_X1 U647 ( .A1(n547), .A2(KEYINPUT78), .ZN(n550) );
  NAND2_X1 U648 ( .A1(n354), .A2(KEYINPUT47), .ZN(n548) );
  INV_X1 U649 ( .A(KEYINPUT78), .ZN(n551) );
  NAND2_X1 U650 ( .A1(n548), .A2(n551), .ZN(n549) );
  NAND2_X1 U651 ( .A1(n550), .A2(n549), .ZN(n553) );
  AND2_X1 U652 ( .A1(n551), .A2(n682), .ZN(n552) );
  AND2_X1 U653 ( .A1(n598), .A2(n681), .ZN(n554) );
  NOR2_X1 U654 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U655 ( .A(n558), .B(KEYINPUT36), .ZN(n559) );
  NAND2_X1 U656 ( .A1(n559), .A2(n627), .ZN(n689) );
  XOR2_X1 U657 ( .A(KEYINPUT48), .B(KEYINPUT80), .Z(n560) );
  XNOR2_X1 U658 ( .A(n561), .B(n560), .ZN(n572) );
  NOR2_X1 U659 ( .A1(n613), .A2(n562), .ZN(n563) );
  XNOR2_X1 U660 ( .A(KEYINPUT106), .B(n563), .ZN(n565) );
  INV_X1 U661 ( .A(n627), .ZN(n564) );
  NAND2_X1 U662 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U663 ( .A(KEYINPUT43), .B(n566), .ZN(n567) );
  NAND2_X1 U664 ( .A1(n567), .A2(n348), .ZN(n568) );
  XNOR2_X1 U665 ( .A(KEYINPUT107), .B(n568), .ZN(n735) );
  NAND2_X1 U666 ( .A1(n676), .A2(n569), .ZN(n692) );
  NOR2_X1 U667 ( .A1(G898), .A2(n457), .ZN(n713) );
  INV_X1 U668 ( .A(n574), .ZN(n575) );
  NAND2_X1 U669 ( .A1(n713), .A2(n575), .ZN(n576) );
  XNOR2_X1 U670 ( .A(KEYINPUT91), .B(n576), .ZN(n577) );
  NOR2_X1 U671 ( .A1(n578), .A2(n577), .ZN(n579) );
  INV_X1 U672 ( .A(KEYINPUT0), .ZN(n581) );
  INV_X1 U673 ( .A(n597), .ZN(n584) );
  NAND2_X1 U674 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U675 ( .A(n585), .B(KEYINPUT22), .ZN(n589) );
  NOR2_X1 U676 ( .A1(n589), .A2(n627), .ZN(n593) );
  NOR2_X1 U677 ( .A1(n623), .A2(n598), .ZN(n586) );
  NAND2_X1 U678 ( .A1(n593), .A2(n586), .ZN(n669) );
  NOR2_X1 U679 ( .A1(n598), .A2(n594), .ZN(n587) );
  NAND2_X1 U680 ( .A1(n627), .A2(n587), .ZN(n588) );
  OR2_X1 U681 ( .A1(n589), .A2(n588), .ZN(n592) );
  XNOR2_X1 U682 ( .A(KEYINPUT32), .B(KEYINPUT65), .ZN(n590) );
  XNOR2_X1 U683 ( .A(n593), .B(KEYINPUT104), .ZN(n595) );
  NAND2_X1 U684 ( .A1(n598), .A2(n605), .ZN(n600) );
  NAND2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n621) );
  NOR2_X1 U686 ( .A1(n621), .A2(n347), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n606), .B(KEYINPUT31), .ZN(n686) );
  NOR2_X1 U688 ( .A1(n347), .A2(n607), .ZN(n608) );
  NAND2_X1 U689 ( .A1(n626), .A2(n608), .ZN(n671) );
  NAND2_X1 U690 ( .A1(n609), .A2(KEYINPUT2), .ZN(n651) );
  AND2_X1 U691 ( .A1(n354), .A2(n610), .ZN(n611) );
  XNOR2_X1 U692 ( .A(n611), .B(KEYINPUT119), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n618), .B(KEYINPUT120), .ZN(n620) );
  INV_X1 U697 ( .A(n619), .ZN(n643) );
  NAND2_X1 U698 ( .A1(n620), .A2(n643), .ZN(n638) );
  INV_X1 U699 ( .A(n621), .ZN(n633) );
  AND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n624), .B(KEYINPUT49), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n631) );
  NOR2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U704 ( .A(n629), .B(KEYINPUT50), .ZN(n630) );
  NOR2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U707 ( .A(KEYINPUT51), .B(n634), .ZN(n636) );
  INV_X1 U708 ( .A(n635), .ZN(n642) );
  NAND2_X1 U709 ( .A1(n636), .A2(n642), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U711 ( .A(KEYINPUT52), .B(n639), .Z(n640) );
  NOR2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n645) );
  AND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n646) );
  INV_X1 U715 ( .A(KEYINPUT2), .ZN(n649) );
  NAND2_X1 U716 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U717 ( .A1(n708), .A2(G475), .ZN(n658) );
  INV_X1 U718 ( .A(n654), .ZN(n656) );
  XOR2_X1 U719 ( .A(KEYINPUT66), .B(KEYINPUT59), .Z(n655) );
  NOR2_X1 U720 ( .A1(n457), .A2(G952), .ZN(n659) );
  XNOR2_X1 U721 ( .A(n659), .B(KEYINPUT84), .ZN(n712) );
  INV_X1 U722 ( .A(n712), .ZN(n698) );
  NAND2_X1 U723 ( .A1(n660), .A2(n698), .ZN(n662) );
  XNOR2_X1 U724 ( .A(KEYINPUT60), .B(KEYINPUT123), .ZN(n661) );
  XNOR2_X1 U725 ( .A(n662), .B(n661), .ZN(G60) );
  NAND2_X1 U726 ( .A1(n708), .A2(G472), .ZN(n666) );
  XOR2_X1 U727 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n664) );
  XOR2_X1 U728 ( .A(G101), .B(KEYINPUT115), .Z(n668) );
  XNOR2_X1 U729 ( .A(n669), .B(n668), .ZN(G3) );
  INV_X1 U730 ( .A(n681), .ZN(n684) );
  NOR2_X1 U731 ( .A1(n684), .A2(n671), .ZN(n670) );
  XOR2_X1 U732 ( .A(G104), .B(n670), .Z(G6) );
  NOR2_X1 U733 ( .A1(n687), .A2(n671), .ZN(n673) );
  XNOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n672) );
  XNOR2_X1 U735 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U736 ( .A(G107), .B(n674), .ZN(G9) );
  XOR2_X1 U737 ( .A(n675), .B(G110), .Z(G12) );
  XOR2_X1 U738 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n678) );
  NAND2_X1 U739 ( .A1(n682), .A2(n676), .ZN(n677) );
  XNOR2_X1 U740 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U741 ( .A(G128), .B(n679), .ZN(G30) );
  XOR2_X1 U742 ( .A(G143), .B(n680), .Z(G45) );
  NAND2_X1 U743 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U744 ( .A(n683), .B(G146), .ZN(G48) );
  NOR2_X1 U745 ( .A1(n684), .A2(n686), .ZN(n685) );
  XOR2_X1 U746 ( .A(G113), .B(n685), .Z(G15) );
  NOR2_X1 U747 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U748 ( .A(G116), .B(n688), .Z(G18) );
  XNOR2_X1 U749 ( .A(KEYINPUT117), .B(KEYINPUT37), .ZN(n690) );
  XNOR2_X1 U750 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U751 ( .A(G125), .B(n691), .ZN(G27) );
  XNOR2_X1 U752 ( .A(G134), .B(n692), .ZN(G36) );
  XOR2_X1 U753 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n695) );
  XNOR2_X1 U754 ( .A(n693), .B(KEYINPUT82), .ZN(n694) );
  NAND2_X1 U755 ( .A1(n708), .A2(G469), .ZN(n702) );
  XOR2_X1 U756 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n699) );
  NOR2_X1 U757 ( .A1(n712), .A2(n703), .ZN(G54) );
  XNOR2_X1 U758 ( .A(n704), .B(KEYINPUT124), .ZN(n706) );
  NAND2_X1 U759 ( .A1(G478), .A2(n708), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n707), .A2(n712), .ZN(G63) );
  NAND2_X1 U762 ( .A1(G217), .A2(n708), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n712), .A2(n711), .ZN(G66) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n721) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n715) );
  XNOR2_X1 U767 ( .A(KEYINPUT61), .B(n715), .ZN(n716) );
  NAND2_X1 U768 ( .A1(n716), .A2(G898), .ZN(n719) );
  NAND2_X1 U769 ( .A1(n349), .A2(n457), .ZN(n718) );
  NAND2_X1 U770 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U771 ( .A(n721), .B(n720), .ZN(G69) );
  XNOR2_X1 U772 ( .A(n723), .B(KEYINPUT125), .ZN(n724) );
  NAND2_X1 U773 ( .A1(n724), .A2(n457), .ZN(n725) );
  XNOR2_X1 U774 ( .A(n725), .B(KEYINPUT126), .ZN(n731) );
  XNOR2_X1 U775 ( .A(G227), .B(n726), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n727), .A2(G900), .ZN(n728) );
  XOR2_X1 U777 ( .A(KEYINPUT127), .B(n728), .Z(n729) );
  NAND2_X1 U778 ( .A1(G953), .A2(n729), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n731), .A2(n730), .ZN(G72) );
  XOR2_X1 U780 ( .A(n732), .B(G131), .Z(G33) );
  XOR2_X1 U781 ( .A(n733), .B(G122), .Z(G24) );
  XOR2_X1 U782 ( .A(G119), .B(n734), .Z(G21) );
  XOR2_X1 U783 ( .A(G140), .B(n735), .Z(n736) );
  XNOR2_X1 U784 ( .A(KEYINPUT118), .B(n736), .ZN(G42) );
  XOR2_X1 U785 ( .A(G137), .B(n737), .Z(G39) );
endmodule

