//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G68), .B2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n206), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n230), .A2(new_n204), .A3(new_n231), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n226), .A2(new_n229), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT64), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n213), .A2(G97), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n209), .A2(G107), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(new_n231), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G238), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n253), .A2(new_n209), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT65), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n253), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(KEYINPUT65), .A3(new_n265), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n268), .A2(new_n271), .B1(new_n223), .B2(G1698), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G226), .A2(G1698), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n263), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n259), .B(new_n262), .C1(new_n275), .C2(new_n255), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G169), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n277), .A2(G179), .A3(new_n278), .ZN(new_n282));
  INV_X1    g0082(.A(G169), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(new_n277), .B2(new_n278), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT14), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n281), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n231), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n291), .A2(new_n217), .B1(new_n204), .B2(G68), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n204), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n219), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n289), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT11), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n298), .A2(new_n204), .A3(G1), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n300), .A2(KEYINPUT12), .A3(G68), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT12), .ZN(new_n302));
  INV_X1    g0102(.A(G68), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n289), .B1(new_n203), .B2(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n301), .A2(new_n304), .B1(new_n306), .B2(new_n303), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n297), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n287), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n268), .A2(new_n271), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G238), .A2(G1698), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n311), .B(new_n312), .C1(new_n223), .C2(G1698), .ZN(new_n313));
  INV_X1    g0113(.A(new_n255), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n313), .B(new_n314), .C1(G107), .C2(new_n311), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(new_n262), .C1(new_n220), .C2(new_n257), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n283), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n305), .A2(G77), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT68), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n300), .A2(G77), .ZN(new_n320));
  INV_X1    g0120(.A(new_n289), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT8), .B(G58), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n323), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n324));
  XOR2_X1   g0124(.A(KEYINPUT15), .B(G87), .Z(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(new_n204), .A3(G33), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n321), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n319), .A2(new_n320), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n317), .B(new_n329), .C1(G179), .C2(new_n316), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n310), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n279), .A2(G200), .ZN(new_n332));
  INV_X1    g0132(.A(G190), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n279), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(new_n309), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n331), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n222), .A2(new_n303), .ZN(new_n337));
  NOR2_X1   g0137(.A1(G58), .A2(G68), .ZN(new_n338));
  OAI21_X1  g0138(.A(G20), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n290), .A2(G159), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n269), .A2(KEYINPUT69), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT69), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n345));
  AOI21_X1  g0145(.A(G33), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT70), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT70), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT69), .B(KEYINPUT3), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n349), .B(new_n350), .C1(new_n351), .C2(G33), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n268), .A2(new_n204), .A3(new_n271), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n348), .A2(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n342), .B1(new_n355), .B2(new_n303), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n343), .A2(new_n345), .A3(G33), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(new_n204), .A3(new_n270), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n303), .B1(new_n360), .B2(KEYINPUT7), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n267), .B1(new_n351), .B2(G33), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(new_n354), .A3(new_n204), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n341), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n321), .B1(new_n364), .B2(KEYINPUT16), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n323), .A2(new_n299), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n306), .B2(new_n323), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT71), .ZN(new_n370));
  NOR2_X1   g0170(.A1(G223), .A2(G1698), .ZN(new_n371));
  INV_X1    g0171(.A(G1698), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(G226), .ZN(new_n373));
  AOI211_X1 g0173(.A(new_n371), .B(new_n373), .C1(new_n359), .C2(new_n270), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n253), .A2(new_n207), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n370), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n359), .A2(new_n270), .ZN(new_n377));
  INV_X1    g0177(.A(new_n371), .ZN(new_n378));
  INV_X1    g0178(.A(new_n373), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n375), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(KEYINPUT71), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n376), .A2(new_n314), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n261), .B1(new_n258), .B2(G232), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(G190), .A3(new_n384), .ZN(new_n385));
  AND3_X1   g0185(.A1(new_n366), .A2(new_n369), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(KEYINPUT73), .A2(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n384), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G200), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT73), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT17), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n386), .A2(new_n387), .A3(new_n389), .A4(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n368), .B1(new_n358), .B2(new_n365), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n394), .A2(new_n389), .A3(new_n387), .A4(new_n385), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(new_n390), .A3(new_n391), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n394), .ZN(new_n398));
  INV_X1    g0198(.A(G179), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n383), .A2(new_n399), .A3(new_n384), .ZN(new_n400));
  AOI21_X1  g0200(.A(G169), .B1(new_n383), .B2(new_n384), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT72), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT72), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n388), .A2(new_n283), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n383), .A2(new_n399), .A3(new_n384), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n398), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT72), .B1(new_n400), .B2(new_n401), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n404), .A2(new_n403), .A3(new_n405), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n394), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT18), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n397), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n372), .A2(G222), .ZN(new_n415));
  XOR2_X1   g0215(.A(KEYINPUT66), .B(G223), .Z(new_n416));
  OAI211_X1 g0216(.A(new_n311), .B(new_n415), .C1(new_n372), .C2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(new_n314), .C1(G77), .C2(new_n311), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(new_n262), .C1(new_n218), .C2(new_n257), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n419), .A2(new_n283), .ZN(new_n420));
  INV_X1    g0220(.A(G150), .ZN(new_n421));
  NOR3_X1   g0221(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n421), .A2(new_n291), .B1(new_n422), .B2(new_n204), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n322), .A2(new_n293), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n289), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n300), .A2(new_n217), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n305), .B2(new_n217), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n427), .A2(KEYINPUT67), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(KEYINPUT67), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n419), .B2(G179), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n420), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n414), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n419), .A2(new_n333), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT9), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n419), .A2(G200), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n430), .A2(new_n437), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n436), .A2(new_n438), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT10), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n316), .A2(G200), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(new_n328), .C1(new_n333), .C2(new_n316), .ZN(new_n444));
  AND4_X1   g0244(.A1(new_n336), .A2(new_n435), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G45), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G1), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n255), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(new_n214), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n377), .A2(G257), .A3(G1698), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT86), .ZN(new_n455));
  AOI21_X1  g0255(.A(G1698), .B1(new_n359), .B2(new_n270), .ZN(new_n456));
  XOR2_X1   g0256(.A(KEYINPUT87), .B(G294), .Z(new_n457));
  AOI22_X1  g0257(.A1(new_n456), .A2(G250), .B1(G33), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT86), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n377), .A2(new_n459), .A3(G257), .A4(G1698), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n455), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n453), .B1(new_n461), .B2(new_n314), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n448), .B(G274), .C1(new_n450), .C2(new_n449), .ZN(new_n463));
  AOI21_X1  g0263(.A(G169), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n462), .A2(new_n463), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(new_n399), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT23), .B1(new_n204), .B2(G107), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT23), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(new_n213), .A3(G20), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n471), .B(KEYINPUT82), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n377), .A2(KEYINPUT22), .A3(new_n204), .A4(G87), .ZN(new_n473));
  AOI211_X1 g0273(.A(G20), .B(new_n207), .C1(new_n268), .C2(new_n271), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n472), .B(new_n473), .C1(new_n474), .C2(KEYINPUT22), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT83), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n311), .A2(new_n204), .A3(G87), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT83), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(new_n472), .A4(new_n473), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n476), .A2(KEYINPUT24), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT24), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n475), .A2(KEYINPUT83), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n289), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT25), .B1(new_n299), .B2(new_n213), .ZN(new_n486));
  XOR2_X1   g0286(.A(new_n486), .B(KEYINPUT85), .Z(new_n487));
  NAND3_X1  g0287(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n213), .ZN(new_n488));
  XOR2_X1   g0288(.A(new_n488), .B(KEYINPUT84), .Z(new_n489));
  INV_X1    g0289(.A(KEYINPUT74), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n253), .A2(G1), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n299), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n491), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n289), .B1(new_n493), .B2(KEYINPUT74), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n487), .A2(new_n489), .B1(G107), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n485), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n466), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n462), .A2(new_n333), .A3(new_n463), .ZN(new_n499));
  AOI21_X1  g0299(.A(G200), .B1(new_n462), .B2(new_n463), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n485), .B(new_n496), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT88), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT88), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n498), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n448), .A2(new_n260), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n255), .B(new_n507), .C1(G250), .C2(new_n448), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT77), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n377), .A2(G244), .A3(G1698), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT78), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n456), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n377), .A2(KEYINPUT78), .A3(G244), .A4(G1698), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n509), .B1(new_n515), .B2(new_n314), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G190), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n516), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n377), .A2(new_n204), .A3(G68), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n293), .A2(new_n209), .ZN(new_n523));
  AOI21_X1  g0323(.A(G20), .B1(new_n263), .B2(KEYINPUT19), .ZN(new_n524));
  XNOR2_X1  g0324(.A(KEYINPUT79), .B(G87), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n525), .A2(G97), .A3(G107), .ZN(new_n526));
  OAI221_X1 g0326(.A(new_n522), .B1(KEYINPUT19), .B2(new_n523), .C1(new_n524), .C2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n325), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n527), .A2(new_n289), .B1(new_n299), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n495), .A2(G87), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n516), .A2(KEYINPUT81), .A3(G190), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n519), .A2(new_n521), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n495), .A2(new_n325), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n534), .B(KEYINPUT80), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(new_n529), .B1(new_n516), .B2(new_n399), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(G169), .B2(new_n516), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n208), .B1(new_n268), .B2(new_n271), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT4), .ZN(new_n540));
  OAI21_X1  g0340(.A(G1698), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G283), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n362), .B2(new_n220), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n311), .A2(KEYINPUT4), .A3(G244), .A4(new_n372), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n314), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n463), .B1(new_n452), .B2(new_n210), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT75), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT75), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n549), .B(new_n463), .C1(new_n452), .C2(new_n210), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n546), .A2(KEYINPUT76), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT76), .B1(new_n546), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g0354(.A(G190), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n290), .A2(G77), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT6), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n209), .A2(new_n213), .ZN(new_n558));
  NOR2_X1   g0358(.A1(G97), .A2(G107), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n557), .B2(new_n246), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G20), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n556), .B(new_n562), .C1(new_n355), .C2(new_n213), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n563), .A2(new_n289), .B1(G97), .B2(new_n495), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n299), .A2(new_n209), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n551), .B1(new_n545), .B2(new_n314), .ZN(new_n567));
  INV_X1    g0367(.A(G200), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n546), .A2(new_n552), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT76), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n567), .A2(KEYINPUT76), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n283), .A3(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n564), .A2(new_n565), .B1(new_n567), .B2(new_n399), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n555), .A2(new_n570), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT21), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n492), .A2(G116), .A3(new_n494), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n542), .B(new_n204), .C1(G33), .C2(new_n209), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n580), .B(new_n289), .C1(new_n204), .C2(G116), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT20), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  OAI221_X1 g0384(.A(new_n579), .B1(G116), .B2(new_n300), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G169), .ZN(new_n586));
  INV_X1    g0386(.A(new_n463), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n451), .A2(new_n255), .A3(G270), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n214), .A2(G1698), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n210), .A2(new_n372), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n377), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(G303), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n311), .ZN(new_n593));
  AOI211_X1 g0393(.A(new_n587), .B(new_n588), .C1(new_n593), .C2(new_n314), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n578), .B1(new_n586), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n588), .B1(new_n593), .B2(new_n314), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n463), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n597), .A2(KEYINPUT21), .A3(G169), .A4(new_n585), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(G179), .A3(new_n585), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n594), .A2(G190), .ZN(new_n601));
  INV_X1    g0401(.A(new_n585), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(new_n602), .C1(new_n568), .C2(new_n594), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n538), .A2(new_n577), .A3(new_n600), .A4(new_n603), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n446), .A2(new_n506), .A3(new_n604), .ZN(G372));
  NAND2_X1  g0405(.A1(new_n498), .A2(new_n600), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n521), .A2(new_n531), .A3(new_n517), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n606), .A2(new_n577), .A3(new_n501), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n575), .A2(new_n576), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT26), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(new_n537), .A4(new_n607), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n533), .A2(new_n537), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT26), .B1(new_n613), .B2(new_n609), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n608), .A2(new_n537), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n445), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n332), .B(new_n308), .C1(new_n333), .C2(new_n279), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n395), .B(new_n392), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n331), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n409), .A2(new_n413), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g0421(.A(new_n442), .B(KEYINPUT89), .Z(new_n622));
  AOI21_X1  g0422(.A(new_n432), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n616), .A2(new_n623), .ZN(G369));
  NOR2_X1   g0424(.A1(new_n298), .A2(G20), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n203), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n627), .A2(G213), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G343), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n630), .B(KEYINPUT90), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n485), .B2(new_n496), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n506), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n631), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n466), .A2(new_n497), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n600), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n631), .A2(new_n602), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n600), .A2(new_n603), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n639), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G330), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n503), .A2(new_n505), .A3(new_n638), .A4(new_n631), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n466), .A2(new_n497), .A3(new_n631), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n644), .A2(new_n647), .ZN(G399));
  INV_X1    g0448(.A(new_n227), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(G41), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G116), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n526), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n651), .A2(G1), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n230), .B2(new_n651), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT28), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT91), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n537), .A2(new_n607), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT26), .B1(new_n659), .B2(new_n609), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n538), .A2(new_n610), .A3(new_n611), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n608), .A2(new_n537), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n662), .A2(KEYINPUT29), .A3(new_n631), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT29), .B1(new_n615), .B2(new_n631), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G330), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n516), .A2(new_n594), .A3(G179), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n667), .B(new_n462), .C1(new_n553), .C2(new_n554), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT30), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n573), .A2(new_n574), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(KEYINPUT30), .A3(new_n462), .A4(new_n667), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n465), .A2(new_n567), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n399), .A3(new_n597), .A4(new_n520), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n670), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n634), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT31), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT31), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n678), .A3(new_n634), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n570), .A2(new_n555), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n609), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n682), .A2(new_n641), .A3(new_n613), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n503), .A3(new_n505), .A4(new_n631), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n666), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n658), .B1(new_n665), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n675), .A2(new_n678), .A3(new_n634), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n678), .B1(new_n675), .B2(new_n634), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n498), .A2(new_n501), .A3(new_n504), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n504), .B1(new_n498), .B2(new_n501), .ZN(new_n691));
  NOR4_X1   g0491(.A1(new_n604), .A2(new_n690), .A3(new_n691), .A4(new_n634), .ZN(new_n692));
  OAI21_X1  g0492(.A(G330), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n693), .B(KEYINPUT91), .C1(new_n663), .C2(new_n664), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n657), .B1(new_n695), .B2(G1), .ZN(G364));
  NAND2_X1  g0496(.A1(new_n625), .A2(G45), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n651), .A2(G1), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n649), .A2(new_n652), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n311), .A2(new_n227), .ZN(new_n701));
  XOR2_X1   g0501(.A(G355), .B(KEYINPUT92), .Z(new_n702));
  NOR2_X1   g0502(.A1(new_n649), .A2(new_n377), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(G45), .B2(new_n230), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n245), .A2(new_n447), .ZN(new_n705));
  OAI221_X1 g0505(.A(new_n700), .B1(new_n701), .B2(new_n702), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(G13), .A2(G33), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G20), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n231), .B1(G20), .B2(new_n283), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n204), .A2(new_n399), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n714), .A2(new_n568), .A3(G190), .ZN(new_n715));
  INV_X1    g0515(.A(G317), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT33), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n716), .A2(KEYINPUT33), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G179), .A2(G200), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n721), .A2(new_n204), .A3(G190), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n722), .A2(KEYINPUT93), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(KEYINPUT93), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n719), .B1(new_n725), .B2(G329), .ZN(new_n726));
  INV_X1    g0526(.A(G283), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n568), .A2(G179), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(G20), .A3(new_n333), .ZN(new_n729));
  INV_X1    g0529(.A(G322), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n714), .A2(new_n333), .A3(G200), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI221_X1 g0532(.A(new_n726), .B1(new_n727), .B2(new_n729), .C1(new_n730), .C2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(G20), .B1(new_n721), .B2(new_n333), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT95), .ZN(new_n735));
  OR2_X1    g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n457), .ZN(new_n740));
  INV_X1    g0540(.A(G326), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n713), .A2(G190), .A3(G200), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT96), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n739), .A2(new_n740), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n733), .A2(new_n311), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n728), .A2(G20), .A3(G190), .ZN(new_n746));
  INV_X1    g0546(.A(G311), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n714), .A2(G190), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n745), .B1(new_n592), .B2(new_n746), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n746), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n715), .A2(G68), .B1(new_n525), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n213), .B2(new_n729), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n725), .A2(G159), .ZN(new_n754));
  XOR2_X1   g0554(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n755));
  OAI21_X1  g0555(.A(new_n311), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n753), .B(new_n756), .C1(G77), .C2(new_n748), .ZN(new_n757));
  INV_X1    g0557(.A(new_n742), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G50), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n754), .A2(new_n755), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n738), .A2(G97), .B1(G58), .B2(new_n731), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n757), .A2(new_n759), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n750), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n710), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n699), .B(new_n712), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT97), .ZN(new_n766));
  INV_X1    g0566(.A(new_n709), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n642), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n643), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n699), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(G330), .B2(new_n642), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(G396));
  NOR2_X1   g0573(.A1(new_n685), .A2(KEYINPUT100), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n615), .A2(new_n631), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n330), .A2(new_n634), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n444), .B1(new_n328), .B2(new_n631), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(new_n777), .B2(new_n330), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n615), .A2(new_n631), .A3(new_n778), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n774), .A2(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(KEYINPUT100), .A2(new_n685), .B1(new_n780), .B2(new_n781), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n783), .B(new_n698), .C1(new_n784), .C2(new_n774), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n779), .A2(new_n707), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n710), .A2(new_n707), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n219), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G143), .A2(new_n731), .B1(new_n748), .B2(G159), .ZN(new_n789));
  INV_X1    g0589(.A(G137), .ZN(new_n790));
  INV_X1    g0590(.A(new_n715), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(new_n790), .B2(new_n742), .C1(new_n421), .C2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT34), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G132), .ZN(new_n795));
  INV_X1    g0595(.A(new_n725), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n739), .A2(new_n222), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n377), .B1(new_n792), .B2(new_n793), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n729), .A2(new_n303), .B1(new_n746), .B2(new_n217), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT99), .Z(new_n801));
  NOR4_X1   g0601(.A1(new_n797), .A2(new_n798), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n731), .A2(G294), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n749), .A2(new_n652), .B1(new_n791), .B2(new_n727), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT98), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n803), .B1(new_n209), .B2(new_n739), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n796), .A2(new_n747), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n746), .A2(new_n213), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n268), .A2(new_n271), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n811), .B1(new_n207), .B2(new_n729), .C1(new_n592), .C2(new_n742), .ZN(new_n812));
  NOR4_X1   g0612(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n710), .B1(new_n802), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n786), .A2(new_n699), .A3(new_n788), .A4(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n785), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G384));
  NAND3_X1  g0617(.A1(new_n287), .A2(new_n309), .A3(new_n631), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n284), .B(KEYINPUT14), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n308), .B1(new_n819), .B2(new_n282), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n335), .A2(new_n332), .B1(new_n309), .B2(new_n634), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n818), .B(new_n778), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(KEYINPUT40), .B(new_n822), .C1(new_n680), .C2(new_n684), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT105), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT38), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n394), .A2(new_n389), .A3(new_n385), .ZN(new_n826));
  INV_X1    g0626(.A(new_n629), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n394), .A2(new_n827), .ZN(new_n828));
  NOR4_X1   g0628(.A1(new_n412), .A2(new_n826), .A3(KEYINPUT37), .A4(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n826), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n361), .A2(new_n363), .ZN(new_n831));
  OR2_X1    g0631(.A1(KEYINPUT103), .A2(KEYINPUT16), .ZN(new_n832));
  AND3_X1   g0632(.A1(new_n831), .A2(new_n342), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n831), .B2(new_n342), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n833), .A2(new_n834), .A3(new_n321), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT104), .B1(new_n835), .B2(new_n368), .ZN(new_n836));
  INV_X1    g0636(.A(new_n834), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n364), .A2(new_n832), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n837), .A2(new_n289), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT104), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(new_n840), .A3(new_n369), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n836), .A2(new_n629), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n402), .A2(new_n406), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n836), .A2(new_n841), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n830), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n829), .B1(KEYINPUT37), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n842), .B1(new_n620), .B2(new_n618), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n824), .B(new_n825), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n825), .B1(new_n846), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n407), .A2(new_n408), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n412), .A2(KEYINPUT18), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n618), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n842), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n845), .A2(KEYINPUT37), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n412), .A2(new_n828), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(new_n830), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n854), .A2(new_n859), .A3(KEYINPUT38), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n849), .A2(KEYINPUT105), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n823), .A2(new_n848), .A3(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n852), .A2(new_n853), .B1(new_n855), .B2(new_n858), .ZN(new_n863));
  INV_X1    g0663(.A(new_n828), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n857), .B1(new_n856), .B2(new_n830), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n414), .A2(new_n864), .B1(new_n865), .B2(new_n829), .ZN(new_n866));
  XOR2_X1   g0666(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n867));
  AOI22_X1  g0667(.A1(KEYINPUT38), .A2(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n822), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n689), .B2(new_n692), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT40), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n862), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n680), .A2(new_n684), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n445), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n872), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(G330), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(KEYINPUT107), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n665), .A2(new_n445), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n623), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n876), .A2(KEYINPUT107), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT39), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n861), .B2(new_n848), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n866), .A2(new_n867), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT39), .B1(new_n887), .B2(new_n860), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n886), .A2(new_n818), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n861), .A2(new_n848), .ZN(new_n890));
  INV_X1    g0690(.A(new_n776), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n781), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n617), .B1(new_n308), .B2(new_n631), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n310), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n818), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n890), .A2(new_n897), .B1(new_n620), .B2(new_n629), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n889), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n881), .B1(new_n878), .B2(new_n882), .ZN(new_n901));
  OR3_X1    g0701(.A1(new_n884), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n900), .B1(new_n884), .B2(new_n901), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n902), .B(new_n903), .C1(new_n203), .C2(new_n625), .ZN(new_n904));
  OAI211_X1 g0704(.A(G20), .B(new_n252), .C1(new_n561), .C2(KEYINPUT35), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n652), .B(new_n905), .C1(KEYINPUT35), .C2(new_n561), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT36), .Z(new_n907));
  NOR3_X1   g0707(.A1(new_n337), .A2(new_n230), .A3(new_n219), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT101), .Z(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(G50), .B2(new_n303), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(G1), .A3(new_n298), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT102), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n904), .A2(new_n913), .ZN(G367));
  NAND2_X1  g0714(.A1(new_n566), .A2(new_n634), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n577), .A2(new_n915), .B1(new_n610), .B2(new_n634), .ZN(new_n916));
  OR3_X1    g0716(.A1(new_n645), .A2(KEYINPUT42), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n681), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n609), .B1(new_n918), .B2(new_n498), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n631), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT42), .B1(new_n645), .B2(new_n916), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n531), .A2(new_n631), .ZN(new_n923));
  MUX2_X1   g0723(.A(new_n659), .B(new_n537), .S(new_n923), .Z(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT108), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n922), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n922), .A2(KEYINPUT43), .A3(new_n925), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n915), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n682), .A2(new_n931), .B1(new_n609), .B2(new_n631), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n644), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n930), .B(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n650), .B(KEYINPUT41), .Z(new_n935));
  INV_X1    g0735(.A(KEYINPUT44), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT109), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n647), .B2(new_n916), .ZN(new_n938));
  AOI211_X1 g0738(.A(KEYINPUT109), .B(new_n932), .C1(new_n645), .C2(new_n646), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n638), .A2(new_n631), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n690), .A2(new_n691), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n646), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n916), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT109), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n647), .A2(new_n937), .A3(new_n916), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(KEYINPUT44), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n645), .A2(new_n646), .A3(new_n932), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT45), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n940), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n644), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n635), .B(new_n941), .C1(new_n506), .C2(new_n632), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n953), .A2(new_n643), .A3(new_n645), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n643), .B1(new_n953), .B2(new_n645), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n644), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n940), .A2(new_n958), .A3(new_n950), .A4(new_n947), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n952), .A2(new_n695), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n935), .B1(new_n960), .B2(new_n695), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n697), .A2(G1), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n934), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n711), .ZN(new_n964));
  INV_X1    g0764(.A(new_n703), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n241), .A2(new_n965), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n964), .B(new_n966), .C1(new_n649), .C2(new_n325), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n725), .A2(G317), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n457), .A2(new_n715), .B1(new_n748), .B2(G283), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n362), .A3(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n746), .A2(new_n652), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT46), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n732), .A2(new_n592), .B1(new_n209), .B2(new_n729), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n974), .B1(new_n213), .B2(new_n739), .C1(new_n747), .C2(new_n743), .ZN(new_n975));
  INV_X1    g0775(.A(G159), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n311), .B1(new_n749), .B2(new_n217), .C1(new_n976), .C2(new_n791), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n738), .A2(G68), .ZN(new_n978));
  INV_X1    g0778(.A(G143), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n743), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n731), .A2(G150), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n751), .A2(G58), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n729), .A2(new_n219), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n790), .B2(new_n796), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n975), .B1(new_n977), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT110), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n967), .B1(new_n989), .B2(new_n710), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n990), .B(new_n699), .C1(new_n767), .C2(new_n925), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT111), .Z(new_n992));
  NAND2_X1  g0792(.A1(new_n963), .A2(new_n992), .ZN(G387));
  INV_X1    g0793(.A(new_n694), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n662), .A2(KEYINPUT29), .A3(new_n631), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n615), .A2(new_n631), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n995), .B1(new_n996), .B2(KEYINPUT29), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT91), .B1(new_n997), .B2(new_n693), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n957), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n686), .A2(new_n694), .A3(new_n956), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n650), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n637), .A2(new_n709), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n703), .B1(new_n237), .B2(new_n447), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n654), .B2(new_n701), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n322), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(G45), .ZN(new_n1006));
  OAI21_X1  g0806(.A(KEYINPUT50), .B1(new_n322), .B2(G50), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n303), .C2(new_n219), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1004), .B1(new_n653), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n649), .A2(new_n213), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n964), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G50), .A2(new_n731), .B1(new_n748), .B2(G68), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n729), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n362), .B1(G97), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1012), .B(new_n1014), .C1(new_n322), .C2(new_n791), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n739), .A2(new_n528), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(G150), .C2(new_n725), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n751), .A2(G77), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n976), .C2(new_n742), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT113), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G311), .A2(new_n715), .B1(new_n731), .B2(G317), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n592), .B2(new_n749), .C1(new_n743), .C2(new_n730), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT48), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n727), .B2(new_n739), .C1(new_n740), .C2(new_n746), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT49), .Z(new_n1025));
  OAI221_X1 g0825(.A(new_n362), .B1(new_n652), .B2(new_n729), .C1(new_n796), .C2(new_n741), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT114), .Z(new_n1027));
  OAI21_X1  g0827(.A(new_n1020), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1011), .B1(new_n1028), .B2(new_n710), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1002), .A2(new_n1029), .A3(new_n699), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n962), .B1(new_n954), .B2(new_n955), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT112), .Z(new_n1032));
  NAND3_X1  g0832(.A1(new_n1001), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT115), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1030), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n651), .B1(new_n695), .B2(new_n957), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(new_n1000), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT115), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n1032), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1034), .A2(new_n1039), .ZN(G393));
  NAND3_X1  g0840(.A1(new_n952), .A2(KEYINPUT116), .A3(new_n959), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT116), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n951), .A2(new_n1042), .A3(new_n644), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n999), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1044), .A2(new_n650), .A3(new_n960), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n711), .B1(new_n209), .B2(new_n227), .C1(new_n965), .C2(new_n250), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n932), .B2(new_n767), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n796), .A2(new_n730), .B1(new_n213), .B2(new_n729), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n311), .B(new_n1048), .C1(G283), .C2(new_n751), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n738), .A2(G116), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n748), .A2(G294), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n731), .A2(G311), .B1(new_n758), .B2(G317), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT52), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G303), .B2(new_n715), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n796), .A2(new_n979), .B1(new_n303), .B2(new_n746), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT117), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n362), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n1057), .B2(new_n1056), .C1(new_n207), .C2(new_n729), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT118), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n739), .A2(new_n219), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n217), .B2(new_n791), .C1(new_n322), .C2(new_n749), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n731), .A2(G159), .B1(new_n758), .B2(G150), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT51), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1055), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n698), .B(new_n1047), .C1(new_n1066), .C2(new_n710), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n962), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1045), .A2(new_n1069), .ZN(G390));
  INV_X1    g0870(.A(new_n868), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n818), .B(KEYINPUT119), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n662), .A2(new_n631), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n777), .A2(new_n330), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n776), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1071), .B(new_n1072), .C1(new_n1075), .C2(new_n895), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n888), .B1(new_n890), .B2(KEYINPUT39), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n818), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n892), .B2(new_n896), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1076), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n685), .A2(new_n778), .A3(new_n896), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1076), .B(new_n1081), .C1(new_n1077), .C2(new_n1079), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n962), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n707), .B1(new_n886), .B2(new_n888), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n787), .A2(new_n322), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n746), .A2(new_n207), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1088), .B(new_n1061), .C1(G294), .C2(new_n725), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n811), .B1(new_n303), .B2(new_n729), .C1(new_n732), .C2(new_n652), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G97), .B2(new_n748), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1089), .B(new_n1091), .C1(new_n213), .C2(new_n791), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G283), .B2(new_n758), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n731), .A2(G132), .B1(new_n758), .B2(G128), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT120), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(G125), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1096), .B1(new_n796), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G159), .B2(new_n738), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n751), .A2(G150), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT53), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1094), .A2(new_n1095), .B1(KEYINPUT53), .B2(new_n1100), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT54), .B(G143), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n790), .A2(new_n791), .B1(new_n749), .B2(new_n1103), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1102), .A2(new_n811), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1099), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G50), .B2(new_n1013), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n710), .B1(new_n1093), .B2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1086), .A2(new_n699), .A3(new_n1087), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1085), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n445), .A2(G330), .A3(new_n873), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1111), .A2(new_n879), .A3(new_n623), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n896), .B1(new_n685), .B2(new_n778), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n892), .B1(new_n1082), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1113), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n1075), .A3(new_n1081), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1112), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1083), .A2(new_n1084), .A3(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(new_n650), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1112), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1110), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(G378));
  NAND2_X1  g0926(.A1(new_n622), .A2(new_n433), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n430), .A2(new_n629), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1127), .B(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1131), .A2(new_n708), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n731), .A2(G107), .B1(new_n758), .B2(G116), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1013), .A2(G58), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1133), .A2(new_n254), .A3(new_n1018), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n377), .B1(new_n725), .B2(G283), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1136), .B(new_n978), .C1(new_n528), .C2(new_n749), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(G97), .C2(new_n715), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT58), .Z(new_n1139));
  AOI21_X1  g0939(.A(G41), .B1(new_n351), .B2(G33), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n742), .A2(new_n1097), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G132), .A2(new_n715), .B1(new_n748), .B2(G137), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT121), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n731), .A2(G128), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n746), .C2(new_n1103), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1141), .B(new_n1145), .C1(G150), .C2(new_n738), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT59), .ZN(new_n1147));
  AOI21_X1  g0947(.A(G33), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(G41), .B1(new_n725), .B2(G124), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(new_n976), .C2(new_n729), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1139), .B1(G50), .B2(new_n1140), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1152), .A2(new_n710), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n787), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(G50), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1132), .A2(new_n698), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n872), .A2(G330), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n898), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n666), .B1(new_n862), .B2(new_n871), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n889), .B2(new_n898), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1160), .A2(new_n1131), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1131), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1156), .B1(new_n1165), .B2(new_n962), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1160), .A2(new_n1131), .A3(new_n1162), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1131), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n889), .A2(new_n1161), .A3(new_n898), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1167), .A2(KEYINPUT57), .A3(new_n1168), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n650), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT57), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1166), .B1(new_n1174), .B2(new_n1175), .ZN(G375));
  NAND2_X1  g0976(.A1(new_n731), .A2(G137), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n795), .B2(new_n742), .C1(new_n791), .C2(new_n1103), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT122), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1134), .B1(new_n749), .B2(new_n421), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n362), .B(new_n1180), .C1(G159), .C2(new_n751), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(new_n217), .C2(new_n739), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G128), .B2(new_n725), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n751), .A2(G97), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1016), .B1(G116), .B2(new_n715), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n749), .A2(new_n213), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n984), .B(new_n1186), .C1(G294), .C2(new_n758), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n311), .B1(new_n731), .B2(G283), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1185), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G303), .B2(new_n725), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1183), .B1(new_n1184), .B2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT123), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(new_n764), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n896), .A2(new_n708), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1154), .A2(G68), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n698), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1121), .B2(new_n962), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1114), .A2(new_n1116), .A3(new_n1112), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(new_n935), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1197), .B1(new_n1200), .B2(new_n1117), .ZN(G381));
  OR2_X1    g1001(.A1(G375), .A2(G378), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1034), .A2(new_n1039), .A3(new_n772), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n963), .A2(new_n992), .A3(new_n1069), .A4(new_n1045), .ZN(new_n1204));
  OR3_X1    g1004(.A1(new_n1204), .A2(G384), .A3(G381), .ZN(new_n1205));
  OR3_X1    g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(G407));
  OAI211_X1 g1006(.A(G407), .B(G213), .C1(G343), .C2(new_n1202), .ZN(G409));
  NAND2_X1  g1007(.A1(G375), .A2(G378), .ZN(new_n1208));
  INV_X1    g1008(.A(G343), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(G213), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1166), .B(new_n1125), .C1(new_n935), .C2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n816), .A2(KEYINPUT124), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n816), .A2(KEYINPUT124), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT60), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1198), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1114), .A2(new_n1116), .A3(new_n1112), .A4(KEYINPUT60), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1216), .A2(new_n1123), .A3(new_n650), .A4(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1213), .B(new_n1214), .C1(new_n1197), .C2(new_n1218), .ZN(new_n1219));
  AND4_X1   g1019(.A1(KEYINPUT124), .A2(new_n1218), .A3(new_n816), .A4(new_n1197), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1208), .A2(new_n1210), .A3(new_n1212), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT62), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1208), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1209), .A2(G213), .A3(G2897), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT125), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1210), .A2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1226), .B1(new_n1221), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1226), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n1227), .B2(new_n1210), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1225), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT61), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G375), .A2(G378), .B1(G213), .B2(new_n1209), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT62), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n1212), .A4(new_n1222), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1224), .A2(new_n1233), .A3(new_n1234), .A4(new_n1237), .ZN(new_n1238));
  AND4_X1   g1038(.A1(new_n963), .A2(new_n992), .A3(new_n1069), .A4(new_n1045), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n963), .A2(new_n992), .B1(new_n1045), .B2(new_n1069), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT126), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1038), .B1(new_n1037), .B2(new_n1032), .ZN(new_n1242));
  AND4_X1   g1042(.A1(new_n1038), .A2(new_n1001), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1243));
  OAI21_X1  g1043(.A(G396), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1203), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT126), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(G390), .A2(new_n1247), .A3(new_n963), .A4(new_n992), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1241), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1245), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT127), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(G390), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1204), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(KEYINPUT127), .A3(new_n1245), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1249), .A2(new_n1252), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1238), .A2(new_n1257), .ZN(new_n1258));
  AOI221_X4 g1058(.A(new_n1251), .B1(new_n1244), .B2(new_n1203), .C1(new_n1253), .C2(new_n1204), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT127), .B1(new_n1254), .B2(new_n1245), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1249), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1235), .A2(KEYINPUT63), .A3(new_n1212), .A4(new_n1222), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1225), .B2(new_n1232), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1223), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1262), .B(new_n1263), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1258), .A2(new_n1267), .ZN(G405));
  XNOR2_X1  g1068(.A(G375), .B(G378), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(new_n1261), .A3(new_n1249), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(G375), .B(new_n1125), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1256), .A2(new_n1271), .ZN(new_n1272));
  AND3_X1   g1072(.A1(new_n1270), .A2(new_n1221), .A3(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1221), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(G402));
endmodule


