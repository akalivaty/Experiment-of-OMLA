

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782;

  NOR2_X1 U368 ( .A1(n549), .A2(n548), .ZN(n565) );
  INV_X1 U369 ( .A(n660), .ZN(n684) );
  NOR2_X1 U370 ( .A1(n666), .A2(G902), .ZN(n405) );
  XNOR2_X1 U371 ( .A(KEYINPUT79), .B(G110), .ZN(n483) );
  NOR2_X1 U372 ( .A1(G953), .A2(G237), .ZN(n515) );
  NAND2_X1 U373 ( .A1(n344), .A2(n637), .ZN(n639) );
  NOR2_X1 U374 ( .A1(n635), .A2(n634), .ZN(n344) );
  NAND2_X2 U375 ( .A1(n561), .A2(n509), .ZN(n510) );
  XNOR2_X1 U376 ( .A(n472), .B(n471), .ZN(n567) );
  XNOR2_X2 U377 ( .A(n762), .B(n395), .ZN(n394) );
  XNOR2_X1 U378 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n770) );
  NOR2_X1 U379 ( .A1(n355), .A2(n616), .ZN(n345) );
  NOR2_X2 U380 ( .A1(n349), .A2(n347), .ZN(n432) );
  XNOR2_X2 U381 ( .A(G137), .B(KEYINPUT96), .ZN(n388) );
  INV_X2 U382 ( .A(G143), .ZN(n377) );
  NOR2_X2 U383 ( .A1(n632), .A2(n631), .ZN(n635) );
  XNOR2_X2 U384 ( .A(n390), .B(n563), .ZN(n781) );
  NAND2_X2 U385 ( .A1(n698), .A2(n562), .ZN(n390) );
  XNOR2_X2 U386 ( .A(n447), .B(n368), .ZN(n617) );
  OR2_X2 U387 ( .A1(n584), .A2(n423), .ZN(n419) );
  XNOR2_X2 U388 ( .A(n613), .B(n573), .ZN(n584) );
  AND2_X2 U389 ( .A1(n438), .A2(n446), .ZN(n356) );
  NOR2_X2 U390 ( .A1(n684), .A2(n686), .ZN(n719) );
  INV_X1 U391 ( .A(G143), .ZN(n473) );
  INV_X1 U392 ( .A(KEYINPUT109), .ZN(n361) );
  NOR2_X1 U393 ( .A1(n735), .A2(G953), .ZN(n736) );
  NAND2_X1 U394 ( .A1(n444), .A2(n581), .ZN(n640) );
  XNOR2_X1 U395 ( .A(n595), .B(n415), .ZN(n397) );
  NAND2_X1 U396 ( .A1(n781), .A2(KEYINPUT46), .ZN(n351) );
  INV_X1 U397 ( .A(n781), .ZN(n352) );
  NAND2_X1 U398 ( .A1(n350), .A2(n690), .ZN(n349) );
  NOR2_X1 U399 ( .A1(n782), .A2(KEYINPUT46), .ZN(n353) );
  NOR2_X1 U400 ( .A1(n418), .A2(n416), .ZN(n585) );
  XNOR2_X1 U401 ( .A(n381), .B(KEYINPUT39), .ZN(n576) );
  NAND2_X1 U402 ( .A1(n417), .A2(n420), .ZN(n416) );
  AND2_X1 U403 ( .A1(n425), .A2(n424), .ZN(n392) );
  AND2_X1 U404 ( .A1(n564), .A2(n715), .ZN(n358) );
  XNOR2_X1 U405 ( .A(n413), .B(KEYINPUT19), .ZN(n590) );
  NAND2_X1 U406 ( .A1(n443), .A2(n583), .ZN(n612) );
  NOR2_X1 U407 ( .A1(n746), .A2(G902), .ZN(n489) );
  XNOR2_X1 U408 ( .A(n400), .B(n399), .ZN(n398) );
  XNOR2_X1 U409 ( .A(n478), .B(n346), .ZN(n666) );
  XNOR2_X1 U410 ( .A(n383), .B(KEYINPUT25), .ZN(n382) );
  XNOR2_X1 U411 ( .A(n770), .B(G101), .ZN(n481) );
  XNOR2_X1 U412 ( .A(n476), .B(KEYINPUT3), .ZN(n442) );
  XNOR2_X1 U413 ( .A(n389), .B(n460), .ZN(n503) );
  XNOR2_X1 U414 ( .A(G902), .B(KEYINPUT91), .ZN(n389) );
  XNOR2_X1 U415 ( .A(G104), .B(G107), .ZN(n482) );
  XNOR2_X1 U416 ( .A(KEYINPUT5), .B(KEYINPUT78), .ZN(n475) );
  XNOR2_X1 U417 ( .A(n398), .B(n346), .ZN(n746) );
  XNOR2_X2 U418 ( .A(n771), .B(G146), .ZN(n346) );
  NAND2_X1 U419 ( .A1(n348), .A2(n351), .ZN(n347) );
  NAND2_X1 U420 ( .A1(n353), .A2(n352), .ZN(n348) );
  NAND2_X1 U421 ( .A1(n782), .A2(KEYINPUT46), .ZN(n350) );
  XNOR2_X2 U422 ( .A(n380), .B(n566), .ZN(n782) );
  XNOR2_X2 U423 ( .A(n384), .B(n382), .ZN(n470) );
  BUF_X1 U424 ( .A(n446), .Z(n354) );
  INV_X1 U425 ( .A(n610), .ZN(n355) );
  AND2_X2 U426 ( .A1(n665), .A2(n414), .ZN(n607) );
  XNOR2_X1 U427 ( .A(n475), .B(n388), .ZN(n387) );
  BUF_X1 U428 ( .A(n624), .Z(n357) );
  NAND2_X1 U429 ( .A1(n564), .A2(n715), .ZN(n359) );
  NAND2_X1 U430 ( .A1(n564), .A2(n715), .ZN(n718) );
  AND2_X2 U431 ( .A1(n491), .A2(n490), .ZN(n561) );
  AND2_X1 U432 ( .A1(n392), .A2(n391), .ZN(n360) );
  XNOR2_X2 U433 ( .A(n484), .B(n483), .ZN(n761) );
  XNOR2_X1 U434 ( .A(n361), .B(n464), .ZN(n466) );
  XNOR2_X2 U435 ( .A(n606), .B(n605), .ZN(n414) );
  NOR2_X1 U436 ( .A1(n590), .A2(n589), .ZN(n447) );
  BUF_X1 U437 ( .A(n539), .Z(n679) );
  NOR2_X2 U438 ( .A1(n738), .A2(n633), .ZN(n364) );
  BUF_X1 U439 ( .A(n438), .Z(n362) );
  INV_X1 U440 ( .A(n443), .ZN(n363) );
  XNOR2_X2 U441 ( .A(n364), .B(n507), .ZN(n407) );
  OR2_X1 U442 ( .A1(n738), .A2(n375), .ZN(n374) );
  NAND2_X1 U443 ( .A1(n507), .A2(n376), .ZN(n375) );
  XNOR2_X1 U444 ( .A(G119), .B(G116), .ZN(n441) );
  INV_X1 U445 ( .A(KEYINPUT47), .ZN(n428) );
  NOR2_X1 U446 ( .A1(n683), .A2(n452), .ZN(n451) );
  INV_X1 U447 ( .A(G902), .ZN(n505) );
  XNOR2_X1 U448 ( .A(n403), .B(KEYINPUT20), .ZN(n467) );
  XNOR2_X1 U449 ( .A(n517), .B(n485), .ZN(n772) );
  XNOR2_X1 U450 ( .A(n519), .B(n473), .ZN(n520) );
  XNOR2_X1 U451 ( .A(G113), .B(G122), .ZN(n511) );
  XOR2_X1 U452 ( .A(KEYINPUT98), .B(G140), .Z(n512) );
  NOR2_X2 U453 ( .A1(n371), .A2(n370), .ZN(n413) );
  XNOR2_X1 U454 ( .A(n386), .B(n481), .ZN(n477) );
  XNOR2_X1 U455 ( .A(n387), .B(n365), .ZN(n386) );
  XNOR2_X1 U456 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n494) );
  XNOR2_X1 U457 ( .A(G122), .B(KEYINPUT74), .ZN(n493) );
  XNOR2_X1 U458 ( .A(KEYINPUT101), .B(KEYINPUT103), .ZN(n528) );
  XNOR2_X1 U459 ( .A(G116), .B(G107), .ZN(n526) );
  INV_X1 U460 ( .A(G134), .ZN(n474) );
  INV_X1 U461 ( .A(KEYINPUT65), .ZN(n638) );
  NAND2_X1 U462 ( .A1(n392), .A2(n391), .ZN(n698) );
  XNOR2_X1 U463 ( .A(n367), .B(n440), .ZN(n559) );
  INV_X1 U464 ( .A(G478), .ZN(n440) );
  XNOR2_X1 U465 ( .A(n486), .B(n401), .ZN(n400) );
  NOR2_X1 U466 ( .A1(n686), .A2(n428), .ZN(n427) );
  INV_X1 U467 ( .A(G237), .ZN(n504) );
  INV_X1 U468 ( .A(KEYINPUT15), .ZN(n460) );
  NAND2_X1 U469 ( .A1(n584), .A2(n421), .ZN(n417) );
  NOR2_X1 U470 ( .A1(n612), .A2(KEYINPUT108), .ZN(n421) );
  NAND2_X1 U471 ( .A1(n612), .A2(KEYINPUT108), .ZN(n420) );
  AND2_X1 U472 ( .A1(n373), .A2(n715), .ZN(n372) );
  NAND2_X1 U473 ( .A1(n437), .A2(n633), .ZN(n373) );
  INV_X1 U474 ( .A(G472), .ZN(n404) );
  XNOR2_X1 U475 ( .A(G128), .B(G119), .ZN(n448) );
  XNOR2_X1 U476 ( .A(KEYINPUT30), .B(KEYINPUT110), .ZN(n544) );
  NAND2_X1 U477 ( .A1(n467), .A2(G217), .ZN(n383) );
  NAND2_X1 U478 ( .A1(n467), .A2(G221), .ZN(n468) );
  XNOR2_X1 U479 ( .A(n439), .B(KEYINPUT105), .ZN(n717) );
  XNOR2_X1 U480 ( .A(n411), .B(n522), .ZN(n647) );
  XNOR2_X1 U481 ( .A(n521), .B(n523), .ZN(n411) );
  XNOR2_X1 U482 ( .A(n502), .B(n396), .ZN(n393) );
  BUF_X1 U483 ( .A(n722), .Z(n729) );
  XNOR2_X1 U484 ( .A(n666), .B(KEYINPUT62), .ZN(n667) );
  XNOR2_X1 U485 ( .A(n379), .B(n378), .ZN(n751) );
  XNOR2_X1 U486 ( .A(n534), .B(n530), .ZN(n378) );
  XNOR2_X1 U487 ( .A(n533), .B(n531), .ZN(n379) );
  INV_X1 U488 ( .A(G140), .ZN(n663) );
  NAND2_X1 U489 ( .A1(n578), .A2(n436), .ZN(n572) );
  INV_X1 U490 ( .A(KEYINPUT35), .ZN(n415) );
  AND2_X1 U491 ( .A1(n593), .A2(n436), .ZN(n550) );
  XNOR2_X1 U492 ( .A(n746), .B(n745), .ZN(n747) );
  INV_X1 U493 ( .A(n621), .ZN(n422) );
  AND2_X1 U494 ( .A1(n515), .A2(G210), .ZN(n365) );
  AND2_X1 U495 ( .A1(n429), .A2(n538), .ZN(n366) );
  INV_X1 U496 ( .A(n612), .ZN(n705) );
  NOR2_X1 U497 ( .A1(n751), .A2(G902), .ZN(n367) );
  XOR2_X1 U498 ( .A(n591), .B(KEYINPUT0), .Z(n368) );
  INV_X1 U499 ( .A(n715), .ZN(n435) );
  INV_X1 U500 ( .A(KEYINPUT108), .ZN(n423) );
  XOR2_X1 U501 ( .A(n647), .B(n646), .Z(n369) );
  INV_X1 U502 ( .A(KEYINPUT84), .ZN(n452) );
  AND2_X1 U503 ( .A1(n738), .A2(n437), .ZN(n370) );
  NAND2_X1 U504 ( .A1(n374), .A2(n372), .ZN(n371) );
  INV_X1 U505 ( .A(n633), .ZN(n376) );
  XNOR2_X2 U506 ( .A(n394), .B(n393), .ZN(n738) );
  XNOR2_X2 U507 ( .A(G131), .B(KEYINPUT69), .ZN(n519) );
  NAND2_X1 U508 ( .A1(n576), .A2(n684), .ZN(n380) );
  NAND2_X1 U509 ( .A1(n565), .A2(n564), .ZN(n381) );
  NAND2_X1 U510 ( .A1(n654), .A2(n505), .ZN(n384) );
  XNOR2_X1 U511 ( .A(n385), .B(n772), .ZN(n654) );
  XNOR2_X1 U512 ( .A(n456), .B(n457), .ZN(n385) );
  NAND2_X1 U513 ( .A1(n503), .A2(G234), .ZN(n403) );
  NAND2_X1 U514 ( .A1(n358), .A2(n426), .ZN(n391) );
  XNOR2_X2 U515 ( .A(n496), .B(n495), .ZN(n762) );
  XNOR2_X2 U516 ( .A(n442), .B(n441), .ZN(n496) );
  XNOR2_X1 U517 ( .A(n761), .B(n481), .ZN(n395) );
  XNOR2_X1 U518 ( .A(n492), .B(KEYINPUT73), .ZN(n396) );
  NAND2_X1 U519 ( .A1(n607), .A2(n397), .ZN(n410) );
  XNOR2_X1 U520 ( .A(n397), .B(G122), .ZN(G24) );
  XNOR2_X1 U521 ( .A(n481), .B(KEYINPUT73), .ZN(n399) );
  INV_X1 U522 ( .A(n761), .ZN(n401) );
  XNOR2_X2 U523 ( .A(n534), .B(n519), .ZN(n771) );
  NAND2_X1 U524 ( .A1(n402), .A2(n551), .ZN(n552) );
  NAND2_X1 U525 ( .A1(n402), .A2(n451), .ZN(n553) );
  NAND2_X1 U526 ( .A1(n543), .A2(n542), .ZN(n402) );
  XNOR2_X2 U527 ( .A(n405), .B(n404), .ZN(n703) );
  BUF_X1 U528 ( .A(n654), .Z(n406) );
  NAND2_X1 U529 ( .A1(n419), .A2(n422), .ZN(n418) );
  XNOR2_X1 U530 ( .A(n434), .B(n558), .ZN(n433) );
  NAND2_X1 U531 ( .A1(n430), .A2(n366), .ZN(n543) );
  NAND2_X1 U532 ( .A1(n539), .A2(KEYINPUT47), .ZN(n430) );
  XNOR2_X2 U533 ( .A(n510), .B(KEYINPUT82), .ZN(n539) );
  XNOR2_X2 U534 ( .A(n407), .B(KEYINPUT38), .ZN(n564) );
  BUF_X1 U535 ( .A(n703), .Z(n408) );
  NOR2_X2 U536 ( .A1(n617), .A2(n596), .ZN(n409) );
  XNOR2_X2 U537 ( .A(n409), .B(KEYINPUT22), .ZN(n624) );
  XNOR2_X1 U538 ( .A(n410), .B(n608), .ZN(n627) );
  NAND2_X1 U539 ( .A1(n703), .A2(n715), .ZN(n545) );
  XNOR2_X1 U540 ( .A(n412), .B(n514), .ZN(n518) );
  XNOR2_X1 U541 ( .A(n516), .B(n513), .ZN(n412) );
  XNOR2_X2 U542 ( .A(n602), .B(n601), .ZN(n665) );
  XNOR2_X1 U543 ( .A(n414), .B(G110), .ZN(G12) );
  NAND2_X1 U544 ( .A1(n584), .A2(n705), .ZN(n609) );
  NAND2_X1 U545 ( .A1(n717), .A2(KEYINPUT41), .ZN(n424) );
  NAND2_X1 U546 ( .A1(n718), .A2(KEYINPUT41), .ZN(n425) );
  NOR2_X1 U547 ( .A1(n717), .A2(KEYINPUT41), .ZN(n426) );
  NAND2_X1 U548 ( .A1(n660), .A2(n427), .ZN(n429) );
  NAND2_X1 U549 ( .A1(n431), .A2(n557), .ZN(n434) );
  NAND2_X1 U550 ( .A1(n554), .A2(n553), .ZN(n431) );
  NAND2_X1 U551 ( .A1(n432), .A2(n433), .ZN(n445) );
  XNOR2_X2 U552 ( .A(n377), .B(G128), .ZN(n498) );
  XNOR2_X2 U553 ( .A(n498), .B(n474), .ZN(n534) );
  INV_X1 U554 ( .A(n407), .ZN(n436) );
  INV_X1 U555 ( .A(n507), .ZN(n437) );
  NAND2_X1 U556 ( .A1(n438), .A2(n446), .ZN(n632) );
  XNOR2_X1 U557 ( .A(n362), .B(n776), .ZN(n774) );
  XNOR2_X2 U558 ( .A(n640), .B(n582), .ZN(n438) );
  NOR2_X1 U559 ( .A1(n559), .A2(n560), .ZN(n439) );
  NAND2_X1 U560 ( .A1(n546), .A2(n443), .ZN(n547) );
  INV_X1 U561 ( .A(n470), .ZN(n443) );
  NAND2_X1 U562 ( .A1(n614), .A2(n363), .ZN(n603) );
  XNOR2_X1 U563 ( .A(n363), .B(KEYINPUT106), .ZN(n700) );
  XNOR2_X1 U564 ( .A(n445), .B(n575), .ZN(n444) );
  NAND2_X1 U565 ( .A1(n446), .A2(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U566 ( .A1(n354), .A2(n765), .ZN(n755) );
  XNOR2_X2 U567 ( .A(n628), .B(KEYINPUT45), .ZN(n446) );
  XNOR2_X1 U568 ( .A(n449), .B(n448), .ZN(n456) );
  XNOR2_X1 U569 ( .A(n455), .B(n450), .ZN(n449) );
  XNOR2_X2 U570 ( .A(G110), .B(KEYINPUT24), .ZN(n450) );
  XNOR2_X1 U571 ( .A(n748), .B(n747), .ZN(n749) );
  BUF_X1 U572 ( .A(n744), .Z(n750) );
  XNOR2_X2 U573 ( .A(G146), .B(G125), .ZN(n497) );
  AND2_X1 U574 ( .A1(G227), .A2(n765), .ZN(n453) );
  INV_X1 U575 ( .A(KEYINPUT76), .ZN(n558) );
  XNOR2_X1 U576 ( .A(n520), .B(G104), .ZN(n521) );
  XNOR2_X1 U577 ( .A(n485), .B(n453), .ZN(n486) );
  INV_X2 U578 ( .A(G953), .ZN(n765) );
  XNOR2_X1 U579 ( .A(n560), .B(KEYINPUT100), .ZN(n537) );
  XNOR2_X1 U580 ( .A(n545), .B(n544), .ZN(n549) );
  INV_X1 U581 ( .A(n754), .ZN(n650) );
  INV_X1 U582 ( .A(KEYINPUT123), .ZN(n658) );
  NAND2_X1 U583 ( .A1(G234), .A2(n765), .ZN(n454) );
  XOR2_X1 U584 ( .A(KEYINPUT8), .B(n454), .Z(n532) );
  NAND2_X1 U585 ( .A1(n532), .A2(G221), .ZN(n457) );
  XNOR2_X2 U586 ( .A(KEYINPUT95), .B(KEYINPUT23), .ZN(n455) );
  INV_X1 U587 ( .A(KEYINPUT68), .ZN(n458) );
  XNOR2_X1 U588 ( .A(n458), .B(KEYINPUT10), .ZN(n459) );
  XNOR2_X1 U589 ( .A(n497), .B(n459), .ZN(n517) );
  XNOR2_X1 U590 ( .A(n663), .B(G137), .ZN(n485) );
  NAND2_X1 U591 ( .A1(G234), .A2(G237), .ZN(n461) );
  XNOR2_X1 U592 ( .A(n461), .B(KEYINPUT14), .ZN(n465) );
  NAND2_X1 U593 ( .A1(G902), .A2(n465), .ZN(n462) );
  XOR2_X1 U594 ( .A(KEYINPUT94), .B(n462), .Z(n463) );
  NAND2_X1 U595 ( .A1(G953), .A2(n463), .ZN(n586) );
  NOR2_X1 U596 ( .A1(G900), .A2(n586), .ZN(n464) );
  NAND2_X1 U597 ( .A1(G952), .A2(n465), .ZN(n728) );
  NOR2_X1 U598 ( .A1(n728), .A2(G953), .ZN(n587) );
  NOR2_X1 U599 ( .A1(n466), .A2(n587), .ZN(n469) );
  XNOR2_X1 U600 ( .A(n468), .B(KEYINPUT21), .ZN(n699) );
  NOR2_X1 U601 ( .A1(n469), .A2(n699), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n470), .A2(n546), .ZN(n472) );
  INV_X1 U603 ( .A(KEYINPUT70), .ZN(n471) );
  XNOR2_X2 U604 ( .A(G113), .B(KEYINPUT72), .ZN(n476) );
  XNOR2_X1 U605 ( .A(n477), .B(n496), .ZN(n478) );
  NAND2_X1 U606 ( .A1(n567), .A2(n703), .ZN(n480) );
  INV_X1 U607 ( .A(KEYINPUT28), .ZN(n479) );
  XNOR2_X1 U608 ( .A(n480), .B(n479), .ZN(n491) );
  INV_X1 U609 ( .A(n482), .ZN(n484) );
  INV_X1 U610 ( .A(KEYINPUT71), .ZN(n487) );
  XNOR2_X1 U611 ( .A(n487), .B(G469), .ZN(n488) );
  XNOR2_X2 U612 ( .A(n489), .B(n488), .ZN(n613) );
  INV_X1 U613 ( .A(n613), .ZN(n490) );
  XOR2_X1 U614 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n492) );
  XNOR2_X1 U615 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U616 ( .A(n498), .B(n497), .ZN(n501) );
  NAND2_X1 U617 ( .A1(G224), .A2(n765), .ZN(n499) );
  XNOR2_X1 U618 ( .A(n499), .B(KEYINPUT92), .ZN(n500) );
  XNOR2_X1 U619 ( .A(n501), .B(n500), .ZN(n502) );
  INV_X1 U620 ( .A(n503), .ZN(n633) );
  NAND2_X1 U621 ( .A1(n505), .A2(n504), .ZN(n508) );
  NAND2_X1 U622 ( .A1(n508), .A2(G210), .ZN(n506) );
  XNOR2_X1 U623 ( .A(n506), .B(KEYINPUT93), .ZN(n507) );
  NAND2_X1 U624 ( .A1(n508), .A2(G214), .ZN(n715) );
  INV_X1 U625 ( .A(n590), .ZN(n509) );
  XNOR2_X1 U626 ( .A(n512), .B(n511), .ZN(n523) );
  XOR2_X1 U627 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n514) );
  XNOR2_X1 U628 ( .A(KEYINPUT12), .B(KEYINPUT99), .ZN(n513) );
  NAND2_X1 U629 ( .A1(G214), .A2(n515), .ZN(n516) );
  XNOR2_X1 U630 ( .A(n518), .B(n517), .ZN(n522) );
  NOR2_X1 U631 ( .A1(G902), .A2(n647), .ZN(n525) );
  XNOR2_X1 U632 ( .A(KEYINPUT13), .B(G475), .ZN(n524) );
  XNOR2_X1 U633 ( .A(n525), .B(n524), .ZN(n560) );
  INV_X1 U634 ( .A(n537), .ZN(n535) );
  XOR2_X1 U635 ( .A(KEYINPUT102), .B(G122), .Z(n527) );
  XNOR2_X1 U636 ( .A(n527), .B(n526), .ZN(n531) );
  XOR2_X1 U637 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n529) );
  XNOR2_X1 U638 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U639 ( .A1(G217), .A2(n532), .ZN(n533) );
  AND2_X1 U640 ( .A1(n535), .A2(n559), .ZN(n686) );
  INV_X1 U641 ( .A(n559), .ZN(n536) );
  NAND2_X1 U642 ( .A1(n537), .A2(n536), .ZN(n660) );
  INV_X1 U643 ( .A(KEYINPUT85), .ZN(n538) );
  NAND2_X1 U644 ( .A1(KEYINPUT85), .A2(KEYINPUT47), .ZN(n540) );
  NOR2_X1 U645 ( .A1(n719), .A2(n540), .ZN(n541) );
  NAND2_X1 U646 ( .A1(n539), .A2(n541), .ZN(n542) );
  OR2_X1 U647 ( .A1(n613), .A2(n547), .ZN(n548) );
  AND2_X1 U648 ( .A1(n560), .A2(n559), .ZN(n593) );
  AND2_X1 U649 ( .A1(n565), .A2(n550), .ZN(n683) );
  INV_X1 U650 ( .A(n683), .ZN(n551) );
  NAND2_X1 U651 ( .A1(n552), .A2(n452), .ZN(n554) );
  NOR2_X1 U652 ( .A1(n719), .A2(KEYINPUT47), .ZN(n555) );
  XNOR2_X1 U653 ( .A(n555), .B(KEYINPUT77), .ZN(n556) );
  OR2_X1 U654 ( .A1(n556), .A2(n679), .ZN(n557) );
  BUF_X1 U655 ( .A(n561), .Z(n562) );
  XOR2_X1 U656 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n563) );
  XNOR2_X1 U657 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n566) );
  NOR2_X1 U658 ( .A1(n660), .A2(n435), .ZN(n569) );
  BUF_X1 U659 ( .A(n567), .Z(n568) );
  NAND2_X1 U660 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U661 ( .A(n703), .B(KEYINPUT6), .ZN(n621) );
  NOR2_X1 U662 ( .A1(n570), .A2(n621), .ZN(n578) );
  XNOR2_X1 U663 ( .A(KEYINPUT36), .B(KEYINPUT89), .ZN(n571) );
  XNOR2_X1 U664 ( .A(n572), .B(n571), .ZN(n574) );
  INV_X1 U665 ( .A(KEYINPUT1), .ZN(n573) );
  BUF_X1 U666 ( .A(n584), .Z(n706) );
  NAND2_X1 U667 ( .A1(n574), .A2(n706), .ZN(n690) );
  INV_X1 U668 ( .A(KEYINPUT48), .ZN(n575) );
  AND2_X1 U669 ( .A1(n576), .A2(n686), .ZN(n693) );
  INV_X1 U670 ( .A(n706), .ZN(n577) );
  NAND2_X1 U671 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U672 ( .A(n579), .B(KEYINPUT43), .ZN(n580) );
  AND2_X1 U673 ( .A1(n407), .A2(n580), .ZN(n664) );
  NOR2_X1 U674 ( .A1(n693), .A2(n664), .ZN(n581) );
  INV_X1 U675 ( .A(KEYINPUT88), .ZN(n582) );
  INV_X1 U676 ( .A(n699), .ZN(n583) );
  XNOR2_X1 U677 ( .A(n585), .B(KEYINPUT33), .ZN(n722) );
  NOR2_X1 U678 ( .A1(n586), .A2(G898), .ZN(n588) );
  NOR2_X1 U679 ( .A1(n588), .A2(n587), .ZN(n589) );
  INV_X1 U680 ( .A(KEYINPUT67), .ZN(n591) );
  NOR2_X1 U681 ( .A1(n722), .A2(n617), .ZN(n592) );
  XNOR2_X1 U682 ( .A(n592), .B(KEYINPUT34), .ZN(n594) );
  NAND2_X1 U683 ( .A1(n594), .A2(n593), .ZN(n595) );
  OR2_X1 U684 ( .A1(n717), .A2(n699), .ZN(n596) );
  AND2_X1 U685 ( .A1(n706), .A2(n700), .ZN(n597) );
  AND2_X1 U686 ( .A1(n597), .A2(n621), .ZN(n598) );
  NAND2_X1 U687 ( .A1(n624), .A2(n598), .ZN(n602) );
  XNOR2_X1 U688 ( .A(KEYINPUT81), .B(KEYINPUT32), .ZN(n600) );
  INV_X1 U689 ( .A(KEYINPUT66), .ZN(n599) );
  XNOR2_X1 U690 ( .A(n600), .B(n599), .ZN(n601) );
  NOR2_X1 U691 ( .A1(n706), .A2(n603), .ZN(n604) );
  NAND2_X1 U692 ( .A1(n624), .A2(n604), .ZN(n606) );
  INV_X1 U693 ( .A(KEYINPUT107), .ZN(n605) );
  INV_X1 U694 ( .A(KEYINPUT44), .ZN(n608) );
  INV_X1 U695 ( .A(n408), .ZN(n614) );
  NOR2_X1 U696 ( .A1(n609), .A2(n614), .ZN(n712) );
  INV_X1 U697 ( .A(n617), .ZN(n610) );
  NAND2_X1 U698 ( .A1(n712), .A2(n610), .ZN(n611) );
  XNOR2_X1 U699 ( .A(n611), .B(KEYINPUT31), .ZN(n687) );
  NOR2_X1 U700 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n615), .A2(n614), .ZN(n616) );
  OR2_X1 U702 ( .A1(n687), .A2(n345), .ZN(n619) );
  INV_X1 U703 ( .A(n719), .ZN(n618) );
  NAND2_X1 U704 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U705 ( .A(n620), .B(KEYINPUT104), .ZN(n625) );
  OR2_X1 U706 ( .A1(n706), .A2(n700), .ZN(n622) );
  NOR2_X1 U707 ( .A1(n422), .A2(n622), .ZN(n623) );
  NAND2_X1 U708 ( .A1(n357), .A2(n623), .ZN(n673) );
  AND2_X1 U709 ( .A1(n625), .A2(n673), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n356), .A2(n633), .ZN(n629) );
  INV_X1 U712 ( .A(KEYINPUT86), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n629), .A2(n630), .ZN(n637) );
  OR2_X1 U714 ( .A1(n630), .A2(n376), .ZN(n631) );
  AND2_X1 U715 ( .A1(n633), .A2(KEYINPUT2), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n639), .B(n638), .ZN(n645) );
  OR2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n643) );
  INV_X1 U718 ( .A(KEYINPUT80), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n643), .B(n642), .ZN(n696) );
  INV_X1 U720 ( .A(n696), .ZN(n644) );
  AND2_X2 U721 ( .A1(n645), .A2(n644), .ZN(n744) );
  NAND2_X1 U722 ( .A1(n744), .A2(G475), .ZN(n648) );
  INV_X1 U723 ( .A(KEYINPUT59), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n648), .B(n369), .ZN(n651) );
  INV_X1 U725 ( .A(G952), .ZN(n649) );
  AND2_X1 U726 ( .A1(n649), .A2(G953), .ZN(n754) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(n653) );
  INV_X1 U728 ( .A(KEYINPUT60), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n653), .B(n652), .ZN(G60) );
  NAND2_X1 U730 ( .A1(n744), .A2(G217), .ZN(n656) );
  XOR2_X1 U731 ( .A(n406), .B(KEYINPUT122), .Z(n655) );
  XNOR2_X1 U732 ( .A(n656), .B(n655), .ZN(n657) );
  NOR2_X2 U733 ( .A1(n657), .A2(n754), .ZN(n659) );
  XNOR2_X1 U734 ( .A(n659), .B(n658), .ZN(G66) );
  NOR2_X1 U735 ( .A1(n679), .A2(n660), .ZN(n662) );
  XNOR2_X1 U736 ( .A(G146), .B(KEYINPUT115), .ZN(n661) );
  XNOR2_X1 U737 ( .A(n662), .B(n661), .ZN(G48) );
  XNOR2_X1 U738 ( .A(n664), .B(n663), .ZN(G42) );
  XNOR2_X1 U739 ( .A(n665), .B(G119), .ZN(G21) );
  NAND2_X1 U740 ( .A1(n744), .A2(G472), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X2 U742 ( .A1(n669), .A2(n754), .ZN(n672) );
  XNOR2_X1 U743 ( .A(KEYINPUT113), .B(KEYINPUT63), .ZN(n670) );
  XNOR2_X1 U744 ( .A(n670), .B(KEYINPUT90), .ZN(n671) );
  XNOR2_X1 U745 ( .A(n672), .B(n671), .ZN(G57) );
  XNOR2_X1 U746 ( .A(G101), .B(n673), .ZN(G3) );
  NAND2_X1 U747 ( .A1(n345), .A2(n684), .ZN(n674) );
  XNOR2_X1 U748 ( .A(n674), .B(G104), .ZN(G6) );
  XOR2_X1 U749 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n676) );
  NAND2_X1 U750 ( .A1(n345), .A2(n686), .ZN(n675) );
  XNOR2_X1 U751 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U752 ( .A(G107), .B(n677), .ZN(G9) );
  INV_X1 U753 ( .A(n686), .ZN(n678) );
  NOR2_X1 U754 ( .A1(n679), .A2(n678), .ZN(n681) );
  XNOR2_X1 U755 ( .A(KEYINPUT29), .B(KEYINPUT114), .ZN(n680) );
  XNOR2_X1 U756 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U757 ( .A(G128), .B(n682), .ZN(G30) );
  XOR2_X1 U758 ( .A(G143), .B(n683), .Z(G45) );
  NAND2_X1 U759 ( .A1(n687), .A2(n684), .ZN(n685) );
  XNOR2_X1 U760 ( .A(n685), .B(G113), .ZN(G15) );
  NAND2_X1 U761 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U762 ( .A(n688), .B(KEYINPUT116), .ZN(n689) );
  XNOR2_X1 U763 ( .A(G116), .B(n689), .ZN(G18) );
  XNOR2_X1 U764 ( .A(KEYINPUT37), .B(KEYINPUT117), .ZN(n691) );
  XNOR2_X1 U765 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U766 ( .A(G125), .B(n692), .ZN(G27) );
  XOR2_X1 U767 ( .A(G134), .B(n693), .Z(G36) );
  NOR2_X1 U768 ( .A1(n356), .A2(KEYINPUT2), .ZN(n694) );
  XOR2_X1 U769 ( .A(KEYINPUT83), .B(n694), .Z(n695) );
  NOR2_X1 U770 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U771 ( .A(KEYINPUT87), .B(n697), .ZN(n734) );
  NAND2_X1 U772 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U773 ( .A(KEYINPUT49), .B(n701), .ZN(n702) );
  NOR2_X1 U774 ( .A1(n408), .A2(n702), .ZN(n704) );
  XOR2_X1 U775 ( .A(KEYINPUT118), .B(n704), .Z(n710) );
  NOR2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U777 ( .A(KEYINPUT50), .B(n707), .Z(n708) );
  XNOR2_X1 U778 ( .A(KEYINPUT119), .B(n708), .ZN(n709) );
  NOR2_X1 U779 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U781 ( .A(KEYINPUT51), .B(n713), .Z(n714) );
  NOR2_X1 U782 ( .A1(n360), .A2(n714), .ZN(n725) );
  NOR2_X1 U783 ( .A1(n564), .A2(n715), .ZN(n716) );
  NOR2_X1 U784 ( .A1(n717), .A2(n716), .ZN(n721) );
  NOR2_X1 U785 ( .A1(n719), .A2(n359), .ZN(n720) );
  NOR2_X1 U786 ( .A1(n721), .A2(n720), .ZN(n723) );
  NOR2_X1 U787 ( .A1(n723), .A2(n729), .ZN(n724) );
  NOR2_X1 U788 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U789 ( .A(n726), .B(KEYINPUT52), .ZN(n727) );
  NOR2_X1 U790 ( .A1(n728), .A2(n727), .ZN(n731) );
  NOR2_X1 U791 ( .A1(n729), .A2(n360), .ZN(n730) );
  NOR2_X1 U792 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U793 ( .A(KEYINPUT120), .B(n732), .ZN(n733) );
  NAND2_X1 U794 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U795 ( .A(n736), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U796 ( .A1(n744), .A2(G210), .ZN(n740) );
  XOR2_X1 U797 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n737) );
  XNOR2_X1 U798 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U799 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X2 U800 ( .A1(n741), .A2(n754), .ZN(n743) );
  XOR2_X1 U801 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n742) );
  XNOR2_X1 U802 ( .A(n743), .B(n742), .ZN(G51) );
  NAND2_X1 U803 ( .A1(n750), .A2(G469), .ZN(n748) );
  XOR2_X1 U804 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n745) );
  NOR2_X1 U805 ( .A1(n754), .A2(n749), .ZN(G54) );
  NAND2_X1 U806 ( .A1(n750), .A2(G478), .ZN(n752) );
  XNOR2_X1 U807 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U808 ( .A1(n754), .A2(n753), .ZN(G63) );
  XNOR2_X1 U809 ( .A(n755), .B(KEYINPUT124), .ZN(n759) );
  NAND2_X1 U810 ( .A1(G953), .A2(G224), .ZN(n756) );
  XNOR2_X1 U811 ( .A(KEYINPUT61), .B(n756), .ZN(n757) );
  NAND2_X1 U812 ( .A1(n757), .A2(G898), .ZN(n758) );
  NAND2_X1 U813 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U814 ( .A(KEYINPUT126), .B(n760), .ZN(n769) );
  XNOR2_X1 U815 ( .A(n761), .B(KEYINPUT125), .ZN(n763) );
  XNOR2_X1 U816 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U817 ( .A(n764), .B(G101), .ZN(n767) );
  NOR2_X1 U818 ( .A1(n765), .A2(G898), .ZN(n766) );
  NOR2_X1 U819 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U820 ( .A(n769), .B(n768), .ZN(G69) );
  XNOR2_X1 U821 ( .A(n770), .B(n771), .ZN(n773) );
  XNOR2_X1 U822 ( .A(n773), .B(n772), .ZN(n776) );
  NOR2_X1 U823 ( .A1(n774), .A2(G953), .ZN(n775) );
  XNOR2_X1 U824 ( .A(n775), .B(KEYINPUT127), .ZN(n780) );
  XNOR2_X1 U825 ( .A(G227), .B(n776), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n777), .A2(G900), .ZN(n778) );
  NAND2_X1 U827 ( .A1(n778), .A2(G953), .ZN(n779) );
  NAND2_X1 U828 ( .A1(n780), .A2(n779), .ZN(G72) );
  XOR2_X1 U829 ( .A(n781), .B(G137), .Z(G39) );
  XOR2_X1 U830 ( .A(n782), .B(G131), .Z(G33) );
endmodule

