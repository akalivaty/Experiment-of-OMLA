//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT67), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT26), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT26), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(KEYINPUT67), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n202), .A2(KEYINPUT66), .A3(new_n215), .A4(new_n203), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n206), .A2(new_n213), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  AND2_X1   g017(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n214), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n207), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n220), .A2(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n207), .A2(new_n228), .A3(KEYINPUT23), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT25), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(new_n224), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n233), .B1(new_n207), .B2(KEYINPUT23), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(KEYINPUT24), .ZN(new_n237));
  NAND3_X1  g036(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n235), .B1(new_n220), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n217), .B1(new_n231), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G120gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G113gat), .ZN(new_n243));
  INV_X1    g042(.A(G113gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G120gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT1), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G134gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G127gat), .ZN(new_n250));
  INV_X1    g049(.A(G127gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G134gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n249), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n256), .A2(new_n257), .A3(new_n246), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n249), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(new_n247), .B2(new_n253), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT1), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT69), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n248), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT70), .B1(new_n241), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n257), .B1(new_n256), .B2(new_n246), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n263), .A2(KEYINPUT69), .A3(new_n254), .A4(new_n255), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n267), .A2(new_n268), .B1(new_n246), .B2(new_n247), .ZN(new_n269));
  OR2_X1    g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n222), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n207), .A2(new_n228), .A3(KEYINPUT23), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n228), .B1(new_n207), .B2(KEYINPUT23), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n272), .B(new_n232), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n233), .ZN(new_n276));
  INV_X1    g075(.A(new_n238), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n277), .A2(new_n236), .A3(KEYINPUT24), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(new_n271), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n232), .B(new_n234), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n269), .A2(new_n281), .A3(new_n282), .A4(new_n217), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n241), .A2(new_n265), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G227gat), .A2(G233gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT33), .ZN(new_n289));
  XNOR2_X1  g088(.A(G15gat), .B(G43gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(G71gat), .B(G99gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n288), .B(KEYINPUT32), .C1(new_n289), .C2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n267), .A2(new_n268), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n281), .A2(new_n217), .B1(new_n296), .B2(new_n248), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n269), .A2(new_n281), .A3(new_n217), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n297), .B1(KEYINPUT70), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n286), .B1(new_n299), .B2(new_n283), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n288), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n292), .B1(new_n288), .B2(new_n289), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n294), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT71), .B1(new_n288), .B2(KEYINPUT32), .ZN(new_n307));
  AOI211_X1 g106(.A(new_n295), .B(new_n301), .C1(new_n285), .C2(new_n287), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n294), .B(new_n305), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n293), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n299), .A2(new_n286), .A3(new_n283), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT34), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G141gat), .ZN(new_n316));
  INV_X1    g115(.A(G141gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G148gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT2), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G155gat), .ZN(new_n323));
  INV_X1    g122(.A(G162gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT75), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(G155gat), .B2(G162gat), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AND3_X1   g127(.A1(KEYINPUT74), .A2(G155gat), .A3(G162gat), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT74), .B1(G155gat), .B2(G162gat), .ZN(new_n330));
  OR2_X1    g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n322), .A2(new_n328), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n325), .B(new_n327), .C1(new_n329), .C2(new_n330), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n316), .A2(new_n318), .B1(KEYINPUT2), .B2(new_n320), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT76), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g139(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(G148gat), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n340), .B1(new_n343), .B2(new_n316), .ZN(new_n344));
  AND2_X1   g143(.A1(KEYINPUT78), .A2(G162gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(KEYINPUT78), .A2(G162gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT2), .B1(new_n347), .B2(new_n323), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n337), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT79), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n333), .A2(new_n336), .B1(new_n348), .B2(new_n344), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  XNOR2_X1  g154(.A(G197gat), .B(G204gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT22), .ZN(new_n357));
  INV_X1    g156(.A(G211gat), .ZN(new_n358));
  INV_X1    g157(.A(G218gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G211gat), .B(G218gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n355), .B1(new_n363), .B2(KEYINPUT29), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n351), .A2(new_n354), .A3(new_n364), .ZN(new_n365));
  AOI221_X4 g164(.A(KEYINPUT3), .B1(new_n344), .B2(new_n348), .C1(new_n333), .C2(new_n336), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n363), .B1(new_n366), .B2(KEYINPUT29), .ZN(new_n367));
  NAND2_X1  g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G22gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n362), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n361), .B(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n337), .A2(new_n355), .A3(new_n349), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n375), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n352), .B1(new_n377), .B2(new_n355), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n368), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n370), .A2(new_n371), .A3(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT86), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n370), .A2(new_n379), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(KEYINPUT85), .A3(G22gat), .ZN(new_n383));
  XOR2_X1   g182(.A(G78gat), .B(G106gat), .Z(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT31), .B(G50gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(G22gat), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT85), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n381), .A2(new_n383), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n380), .A2(KEYINPUT83), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n387), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n382), .A2(KEYINPUT83), .A3(G22gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n386), .B(KEYINPUT82), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n391), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AOI211_X1 g197(.A(KEYINPUT84), .B(new_n396), .C1(new_n393), .C2(new_n394), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n390), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT72), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n309), .ZN(new_n403));
  INV_X1    g202(.A(new_n313), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n293), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n314), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n351), .A2(new_n265), .A3(new_n354), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n269), .A2(new_n352), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n408), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n410), .B(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n351), .A2(KEYINPUT3), .A3(new_n354), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n366), .A2(new_n269), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(new_n418), .A3(new_n412), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n415), .A2(new_n418), .A3(new_n408), .A4(new_n412), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G1gat), .B(G29gat), .Z(new_n423));
  XNOR2_X1  g222(.A(G57gat), .B(G85gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n407), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n427), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n420), .A2(new_n431), .A3(new_n421), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(new_n420), .B2(new_n421), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n241), .A2(G226gat), .A3(G233gat), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n241), .A2(new_n375), .B1(G226gat), .B2(G233gat), .ZN(new_n438));
  OR3_X1    g237(.A1(new_n437), .A2(new_n438), .A3(new_n363), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n363), .B1(new_n437), .B2(new_n438), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(G8gat), .B(G36gat), .Z(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT73), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n445), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n439), .A2(new_n447), .A3(new_n440), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(KEYINPUT30), .A3(new_n448), .ZN(new_n449));
  OR3_X1    g248(.A1(new_n441), .A2(KEYINPUT30), .A3(new_n445), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT35), .B1(new_n406), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT89), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n427), .B(KEYINPUT87), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n422), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n429), .A3(new_n432), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n430), .A2(new_n458), .A3(new_n435), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT35), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n400), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n314), .A2(new_n405), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n454), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n404), .B1(new_n403), .B2(new_n293), .ZN(new_n466));
  INV_X1    g265(.A(new_n293), .ZN(new_n467));
  AOI211_X1 g266(.A(new_n313), .B(new_n467), .C1(new_n402), .C2(new_n309), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n434), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT81), .B1(new_n434), .B2(KEYINPUT6), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n461), .B1(new_n472), .B2(new_n458), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n469), .A2(new_n473), .A3(KEYINPUT89), .A4(new_n400), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n453), .A2(new_n465), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n412), .B1(new_n415), .B2(new_n418), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT39), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n455), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT39), .B1(new_n411), .B2(new_n413), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n482), .A2(KEYINPUT40), .B1(new_n422), .B2(new_n456), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n482), .B2(KEYINPUT40), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n449), .A2(new_n450), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT88), .B(new_n487), .C1(new_n479), .C2(new_n481), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n483), .A2(new_n485), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n447), .B1(new_n441), .B2(KEYINPUT37), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(KEYINPUT37), .B2(new_n441), .ZN(new_n491));
  INV_X1    g290(.A(new_n448), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(KEYINPUT38), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(KEYINPUT38), .B2(new_n491), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n489), .B(new_n400), .C1(new_n494), .C2(new_n459), .ZN(new_n495));
  INV_X1    g294(.A(new_n400), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n452), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n314), .A2(KEYINPUT36), .A3(new_n405), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT36), .B1(new_n314), .B2(new_n405), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n495), .B(new_n497), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n475), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G183gat), .B(G211gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT96), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(new_n323), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n503), .B(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G57gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n508), .A2(KEYINPUT95), .ZN(new_n509));
  INV_X1    g308(.A(G64gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G71gat), .A2(G78gat), .ZN(new_n512));
  OR2_X1    g311(.A1(G71gat), .A2(G78gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT9), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(new_n508), .B2(new_n510), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n513), .A2(new_n512), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n511), .A2(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G231gat), .A2(G233gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(G127gat), .ZN(new_n526));
  XOR2_X1   g325(.A(G15gat), .B(G22gat), .Z(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(G1gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529));
  INV_X1    g328(.A(G1gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(KEYINPUT16), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT90), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n532), .A2(KEYINPUT90), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n535), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n528), .A2(new_n531), .A3(new_n537), .A4(new_n533), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n536), .A2(KEYINPUT92), .A3(new_n538), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n541), .B(new_n542), .C1(new_n522), .C2(new_n521), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n526), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n526), .A2(new_n543), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n507), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n526), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n526), .A2(new_n543), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(new_n548), .A3(new_n506), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n551));
  XOR2_X1   g350(.A(KEYINPUT97), .B(G92gat), .Z(new_n552));
  INV_X1    g351(.A(G85gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n552), .A2(new_n553), .B1(KEYINPUT8), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT7), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G99gat), .B(G106gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT98), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT99), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT98), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n559), .B(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(new_n557), .A3(new_n555), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n564), .A2(KEYINPUT99), .A3(new_n557), .A4(new_n555), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G29gat), .ZN(new_n569));
  INV_X1    g368(.A(G36gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT14), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT14), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(G29gat), .B2(G36gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(G29gat), .A2(G36gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n571), .A2(new_n573), .A3(KEYINPUT15), .A4(new_n574), .ZN(new_n578));
  XNOR2_X1  g377(.A(G43gat), .B(G50gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n551), .B1(new_n568), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n580), .B2(new_n581), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n580), .A2(new_n584), .A3(new_n581), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n566), .B(new_n567), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(G190gat), .B(G218gat), .Z(new_n590));
  AND2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  XOR2_X1   g395(.A(new_n596), .B(KEYINPUT100), .Z(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n596), .ZN(new_n599));
  OAI22_X1  g398(.A1(new_n591), .A2(new_n592), .B1(KEYINPUT100), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT101), .B1(new_n550), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n546), .A2(new_n549), .ZN(new_n603));
  INV_X1    g402(.A(new_n601), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT91), .Z(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT13), .Z(new_n610));
  INV_X1    g409(.A(new_n542), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT92), .B1(new_n536), .B2(new_n538), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n611), .A2(new_n612), .A3(new_n582), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n541), .A2(new_n542), .B1(new_n580), .B2(new_n581), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n582), .B1(new_n611), .B2(new_n612), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n539), .B1(new_n587), .B2(new_n585), .ZN(new_n617));
  NOR2_X1   g416(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n616), .A2(new_n609), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G113gat), .B(G141gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G197gat), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT11), .B(G169gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n616), .A2(new_n609), .A3(new_n617), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n618), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n621), .A2(KEYINPUT94), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n628), .A2(new_n626), .A3(new_n615), .A4(new_n620), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT94), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n621), .A2(new_n628), .ZN(new_n634));
  INV_X1    g433(.A(new_n626), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(G230gat), .ZN(new_n638));
  INV_X1    g437(.A(G233gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n566), .A2(new_n567), .A3(new_n521), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n561), .A2(new_n520), .A3(new_n565), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT102), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n561), .A2(new_n645), .A3(new_n565), .A4(new_n520), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n641), .A2(new_n643), .A3(new_n644), .A4(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n568), .A2(KEYINPUT10), .A3(new_n520), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n640), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n640), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n643), .A2(new_n646), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n651), .B2(new_n641), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(new_n649), .B2(new_n652), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n607), .A2(new_n637), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n501), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n662), .A2(KEYINPUT103), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(KEYINPUT103), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n472), .A2(KEYINPUT104), .A3(new_n433), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n436), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g471(.A(new_n532), .B1(new_n665), .B2(new_n486), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  OAI211_X1 g473(.A(new_n486), .B(new_n674), .C1(new_n663), .C2(new_n664), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT42), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1325gat));
  AOI21_X1  g478(.A(G15gat), .B1(new_n665), .B2(new_n469), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n681));
  INV_X1    g480(.A(new_n498), .ZN(new_n682));
  INV_X1    g481(.A(new_n499), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT105), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G15gat), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT106), .Z(new_n689));
  AOI21_X1  g488(.A(new_n680), .B1(new_n665), .B2(new_n689), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n665), .A2(new_n496), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  NAND2_X1  g492(.A1(new_n501), .A2(new_n601), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n604), .B1(new_n475), .B2(new_n500), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT44), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n637), .A2(new_n603), .A3(new_n660), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n701), .B2(new_n669), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n697), .A2(new_n700), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n569), .A3(new_n670), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n703), .A2(new_n570), .A3(new_n486), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT46), .Z(new_n708));
  OAI21_X1  g507(.A(G36gat), .B1(new_n701), .B2(new_n451), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(G1329gat));
  NAND2_X1  g509(.A1(new_n682), .A2(new_n683), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n699), .A2(new_n712), .A3(new_n700), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G43gat), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n464), .A2(G43gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n703), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(KEYINPUT47), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(KEYINPUT108), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n696), .A2(new_n687), .A3(new_n700), .A4(new_n698), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(G43gat), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(G43gat), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(KEYINPUT108), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n717), .B1(new_n720), .B2(new_n723), .ZN(G1330gat));
  NAND2_X1  g523(.A1(new_n496), .A2(G50gat), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n703), .A2(new_n496), .ZN(new_n726));
  OAI22_X1  g525(.A1(new_n701), .A2(new_n725), .B1(G50gat), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT48), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  OAI221_X1 g528(.A(new_n729), .B1(G50gat), .B2(new_n726), .C1(new_n701), .C2(new_n725), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1331gat));
  NAND2_X1  g530(.A1(new_n633), .A2(new_n636), .ZN(new_n732));
  INV_X1    g531(.A(new_n660), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n607), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n501), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n669), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n508), .ZN(G1332gat));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT111), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n735), .B(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n451), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n740), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n747), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n739), .A3(new_n745), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1333gat));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n464), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(G71gat), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n687), .A2(G71gat), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n742), .B2(new_n754), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g555(.A1(new_n742), .A2(new_n496), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT112), .B(G78gat), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n603), .A2(new_n732), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n697), .A2(KEYINPUT51), .A3(new_n760), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n761), .A2(KEYINPUT113), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(KEYINPUT113), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  INV_X1    g563(.A(new_n760), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n694), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n762), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n767), .A2(new_n553), .A3(new_n660), .A4(new_n670), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n765), .A2(new_n733), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n699), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n669), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(G1336gat));
  NOR3_X1   g571(.A1(new_n733), .A2(new_n451), .A3(G92gat), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n767), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n696), .A2(new_n486), .A3(new_n698), .A4(new_n769), .ZN(new_n775));
  INV_X1    g574(.A(new_n552), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n766), .A2(new_n761), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n780), .A2(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n774), .A2(new_n779), .B1(new_n781), .B2(new_n778), .ZN(G1337gat));
  OAI21_X1  g581(.A(G99gat), .B1(new_n770), .B2(new_n686), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n464), .A2(G99gat), .A3(new_n733), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1338gat));
  NOR3_X1   g585(.A1(new_n400), .A2(G106gat), .A3(new_n733), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n767), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n696), .A2(new_n496), .A3(new_n698), .A4(new_n769), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT53), .B1(new_n789), .B2(G106gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n789), .A2(new_n792), .A3(G106gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n789), .B2(G106gat), .ZN(new_n794));
  INV_X1    g593(.A(new_n787), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n795), .B1(new_n766), .B2(new_n761), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n791), .B1(new_n797), .B2(new_n798), .ZN(G1339gat));
  NAND4_X1  g598(.A1(new_n602), .A2(new_n606), .A3(new_n637), .A4(new_n733), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n647), .A2(new_n640), .A3(new_n648), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n802), .A2(new_n649), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n649), .A2(new_n803), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n658), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n801), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n656), .B1(new_n649), .B2(new_n803), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n649), .A2(new_n803), .ZN(new_n809));
  OAI211_X1 g608(.A(KEYINPUT55), .B(new_n808), .C1(new_n809), .C2(new_n802), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n807), .A2(new_n657), .A3(new_n810), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n613), .A2(new_n614), .A3(new_n610), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n609), .B1(new_n616), .B2(new_n617), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n625), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n633), .A2(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n811), .A2(new_n604), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n633), .A2(new_n660), .A3(new_n814), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n633), .A2(new_n660), .A3(KEYINPUT115), .A4(new_n814), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n819), .B(new_n820), .C1(new_n637), .C2(new_n811), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n816), .B1(new_n821), .B2(new_n604), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n800), .B1(new_n822), .B2(new_n603), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n823), .A2(new_n469), .A3(new_n400), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n669), .A2(new_n486), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n637), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(new_n244), .ZN(G1340gat));
  NOR2_X1   g627(.A1(new_n826), .A2(new_n733), .ZN(new_n829));
  XNOR2_X1  g628(.A(KEYINPUT116), .B(G120gat), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n829), .B(new_n830), .ZN(G1341gat));
  NOR2_X1   g630(.A1(new_n826), .A2(new_n550), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(new_n251), .ZN(G1342gat));
  NAND3_X1  g632(.A1(new_n824), .A2(new_n601), .A3(new_n825), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(G134gat), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT56), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(G134gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1343gat));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n711), .A2(new_n825), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n400), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n800), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n817), .B1(new_n637), .B2(new_n811), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n604), .ZN(new_n846));
  INV_X1    g645(.A(new_n816), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n603), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n816), .B1(new_n604), .B2(new_n845), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT117), .B1(new_n851), .B2(new_n603), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n843), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT57), .B1(new_n823), .B2(new_n496), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n732), .B(new_n840), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n341), .A2(new_n342), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n670), .B1(new_n684), .B2(new_n685), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n823), .A2(new_n496), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(new_n451), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n823), .A2(new_n496), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n863), .A2(new_n686), .A3(KEYINPUT120), .A4(new_n670), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n732), .A2(new_n317), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n839), .B(new_n857), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n863), .A2(new_n670), .A3(new_n686), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n866), .A2(new_n486), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n868), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n859), .A2(new_n860), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(KEYINPUT118), .A3(new_n870), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n875), .A2(KEYINPUT119), .A3(KEYINPUT58), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT119), .B1(new_n875), .B2(KEYINPUT58), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n867), .B1(new_n876), .B2(new_n877), .ZN(G1344gat));
  OAI21_X1  g677(.A(new_n840), .B1(new_n853), .B2(new_n854), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n879), .A2(KEYINPUT59), .A3(new_n733), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n811), .A2(new_n604), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n815), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n882), .B2(new_n881), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n603), .B1(new_n884), .B2(new_n846), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n496), .B1(new_n885), .B2(new_n844), .ZN(new_n886));
  AOI22_X1  g685(.A1(new_n886), .A2(new_n841), .B1(new_n823), .B2(new_n842), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n840), .A2(new_n660), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT59), .B(G148gat), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n880), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n864), .A2(new_n861), .A3(new_n451), .A4(new_n660), .ZN(new_n891));
  AOI21_X1  g690(.A(G148gat), .B1(new_n891), .B2(KEYINPUT59), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT122), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n315), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n895), .A2(new_n896), .A3(new_n880), .A4(new_n889), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n893), .A2(new_n897), .ZN(G1345gat));
  OAI21_X1  g697(.A(G155gat), .B1(new_n879), .B2(new_n550), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n603), .A2(new_n323), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n865), .B2(new_n900), .ZN(G1346gat));
  AND2_X1   g700(.A1(new_n601), .A2(new_n347), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n862), .A2(new_n864), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT123), .ZN(new_n904));
  OAI22_X1  g703(.A1(new_n879), .A2(new_n604), .B1(new_n346), .B2(new_n345), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1347gat));
  AND2_X1   g705(.A1(new_n823), .A2(new_n669), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n406), .A2(new_n451), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT124), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(G169gat), .B1(new_n911), .B2(new_n732), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n907), .A2(new_n908), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT125), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n907), .A2(new_n915), .A3(new_n908), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n732), .A2(G169gat), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(G1348gat));
  INV_X1    g718(.A(G176gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n911), .A2(new_n920), .A3(new_n660), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n917), .A2(new_n660), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n920), .ZN(G1349gat));
  NAND3_X1  g722(.A1(new_n914), .A2(new_n603), .A3(new_n916), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G183gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n911), .A2(new_n202), .A3(new_n603), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT60), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(KEYINPUT60), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n925), .A2(new_n930), .A3(new_n926), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n911), .A2(new_n203), .A3(new_n601), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n914), .A2(new_n601), .A3(new_n916), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n934), .A2(new_n935), .A3(G190gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n934), .B2(G190gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(G1351gat));
  NOR2_X1   g737(.A1(new_n400), .A2(new_n451), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n907), .A2(new_n686), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n732), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n686), .A2(new_n486), .A3(new_n669), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n887), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n732), .A2(G197gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G1352gat));
  XOR2_X1   g744(.A(KEYINPUT127), .B(G204gat), .Z(new_n946));
  NAND3_X1  g745(.A1(new_n940), .A2(new_n660), .A3(new_n946), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT62), .Z(new_n948));
  NOR3_X1   g747(.A1(new_n887), .A2(new_n733), .A3(new_n942), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n946), .ZN(G1353gat));
  NAND3_X1  g749(.A1(new_n940), .A2(new_n358), .A3(new_n603), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n943), .A2(new_n603), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n952), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(G1354gat));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n359), .A3(new_n601), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n887), .A2(new_n604), .A3(new_n942), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n359), .ZN(G1355gat));
endmodule


