

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755;

  XNOR2_X1 U369 ( .A(KEYINPUT78), .B(KEYINPUT94), .ZN(n360) );
  NOR2_X1 U370 ( .A1(n725), .A2(n406), .ZN(n376) );
  NOR2_X1 U371 ( .A1(n679), .A2(n678), .ZN(n532) );
  AND2_X2 U372 ( .A1(n397), .A2(n375), .ZN(n713) );
  NOR2_X2 U373 ( .A1(n542), .A2(n541), .ZN(n661) );
  XNOR2_X2 U374 ( .A(n455), .B(KEYINPUT0), .ZN(n524) );
  NOR2_X2 U375 ( .A1(n560), .A2(n454), .ZN(n455) );
  NAND2_X2 U376 ( .A1(n400), .A2(n347), .ZN(n398) );
  XNOR2_X2 U377 ( .A(G119), .B(G116), .ZN(n403) );
  XNOR2_X2 U378 ( .A(n404), .B(n403), .ZN(n396) );
  XNOR2_X2 U379 ( .A(n432), .B(G113), .ZN(n404) );
  XNOR2_X2 U380 ( .A(n587), .B(KEYINPUT42), .ZN(n753) );
  XNOR2_X2 U381 ( .A(n490), .B(n440), .ZN(n500) );
  XNOR2_X2 U382 ( .A(n585), .B(n584), .ZN(n708) );
  NOR2_X2 U383 ( .A1(n694), .A2(n688), .ZN(n585) );
  NAND2_X1 U384 ( .A1(n382), .A2(n380), .ZN(n704) );
  INV_X1 U385 ( .A(n360), .ZN(n436) );
  XNOR2_X1 U386 ( .A(KEYINPUT79), .B(KEYINPUT95), .ZN(n435) );
  NAND2_X1 U387 ( .A1(n377), .A2(n620), .ZN(n397) );
  AND2_X1 U388 ( .A1(n385), .A2(n383), .ZN(n382) );
  NOR2_X1 U389 ( .A1(n751), .A2(n656), .ZN(n522) );
  NOR2_X1 U390 ( .A1(n576), .A2(n525), .ZN(n527) );
  XNOR2_X1 U391 ( .A(n557), .B(KEYINPUT114), .ZN(n599) );
  XNOR2_X1 U392 ( .A(n558), .B(n448), .ZN(n560) );
  BUF_X1 U393 ( .A(n573), .Z(n602) );
  XNOR2_X1 U394 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U395 ( .A(n388), .B(n387), .ZN(n718) );
  XNOR2_X1 U396 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U397 ( .A(n597), .B(n356), .ZN(n386) );
  NOR2_X2 U398 ( .A1(G953), .A2(G237), .ZN(n487) );
  INV_X2 U399 ( .A(KEYINPUT3), .ZN(n432) );
  XNOR2_X2 U400 ( .A(n405), .B(n486), .ZN(n736) );
  XNOR2_X2 U401 ( .A(G137), .B(G134), .ZN(n405) );
  XNOR2_X2 U402 ( .A(n602), .B(n583), .ZN(n692) );
  XOR2_X1 U403 ( .A(G122), .B(G104), .Z(n474) );
  NOR2_X1 U404 ( .A1(n649), .A2(n544), .ZN(n545) );
  NAND2_X1 U405 ( .A1(n381), .A2(KEYINPUT86), .ZN(n380) );
  INV_X1 U406 ( .A(n386), .ZN(n381) );
  XNOR2_X1 U407 ( .A(n444), .B(n443), .ZN(n573) );
  INV_X1 U408 ( .A(n673), .ZN(n484) );
  XNOR2_X1 U409 ( .A(n474), .B(KEYINPUT16), .ZN(n419) );
  XNOR2_X1 U410 ( .A(G119), .B(G128), .ZN(n502) );
  XNOR2_X1 U411 ( .A(KEYINPUT99), .B(G110), .ZN(n503) );
  NAND2_X1 U412 ( .A1(n508), .A2(G221), .ZN(n391) );
  XNOR2_X1 U413 ( .A(G137), .B(KEYINPUT100), .ZN(n504) );
  XNOR2_X1 U414 ( .A(n379), .B(KEYINPUT24), .ZN(n505) );
  INV_X1 U415 ( .A(KEYINPUT23), .ZN(n379) );
  XNOR2_X1 U416 ( .A(n365), .B(n364), .ZN(n508) );
  INV_X1 U417 ( .A(KEYINPUT8), .ZN(n364) );
  NAND2_X1 U418 ( .A1(n741), .A2(G234), .ZN(n365) );
  INV_X1 U419 ( .A(n617), .ZN(n406) );
  XOR2_X1 U420 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n472) );
  XNOR2_X1 U421 ( .A(KEYINPUT105), .B(KEYINPUT104), .ZN(n471) );
  XNOR2_X1 U422 ( .A(n425), .B(n470), .ZN(n424) );
  XOR2_X1 U423 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n470) );
  XNOR2_X1 U424 ( .A(n468), .B(n469), .ZN(n425) );
  XNOR2_X1 U425 ( .A(G143), .B(KEYINPUT11), .ZN(n469) );
  XNOR2_X1 U426 ( .A(G113), .B(G131), .ZN(n475) );
  XNOR2_X1 U427 ( .A(n390), .B(G140), .ZN(n389) );
  INV_X1 U428 ( .A(KEYINPUT10), .ZN(n390) );
  XNOR2_X1 U429 ( .A(n369), .B(KEYINPUT33), .ZN(n709) );
  INV_X1 U430 ( .A(KEYINPUT113), .ZN(n372) );
  NOR2_X1 U431 ( .A1(n561), .A2(n676), .ZN(n562) );
  BUF_X1 U432 ( .A(n524), .Z(n537) );
  BUF_X1 U433 ( .A(n571), .Z(n676) );
  XNOR2_X1 U434 ( .A(n513), .B(n512), .ZN(n514) );
  NOR2_X1 U435 ( .A1(n718), .A2(G902), .ZN(n515) );
  NOR2_X1 U436 ( .A1(n384), .A2(n670), .ZN(n383) );
  NOR2_X1 U437 ( .A1(n605), .A2(n606), .ZN(n384) );
  INV_X1 U438 ( .A(G237), .ZN(n442) );
  INV_X1 U439 ( .A(n572), .ZN(n399) );
  INV_X1 U440 ( .A(KEYINPUT6), .ZN(n409) );
  XOR2_X1 U441 ( .A(G107), .B(G122), .Z(n457) );
  XNOR2_X1 U442 ( .A(G116), .B(G134), .ZN(n456) );
  XOR2_X1 U443 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n459) );
  XNOR2_X1 U444 ( .A(G902), .B(KEYINPUT15), .ZN(n614) );
  INV_X1 U445 ( .A(G131), .ZN(n486) );
  NAND2_X1 U446 ( .A1(G234), .A2(G237), .ZN(n449) );
  OR2_X1 U447 ( .A1(n674), .A2(n572), .ZN(n554) );
  INV_X1 U448 ( .A(G902), .ZN(n478) );
  XNOR2_X1 U449 ( .A(KEYINPUT73), .B(G110), .ZN(n439) );
  XNOR2_X1 U450 ( .A(n736), .B(G146), .ZN(n493) );
  XNOR2_X1 U451 ( .A(n366), .B(n441), .ZN(n637) );
  NOR2_X1 U452 ( .A1(n558), .A2(KEYINPUT36), .ZN(n414) );
  XNOR2_X1 U453 ( .A(n418), .B(n354), .ZN(n520) );
  NOR2_X1 U454 ( .A1(n694), .A2(n484), .ZN(n485) );
  INV_X1 U455 ( .A(KEYINPUT1), .ZN(n368) );
  XNOR2_X1 U456 ( .A(n506), .B(n507), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n391), .B(n739), .ZN(n388) );
  NAND2_X1 U458 ( .A1(n362), .A2(n407), .ZN(n375) );
  XNOR2_X1 U459 ( .A(n426), .B(n361), .ZN(n630) );
  XNOR2_X1 U460 ( .A(n476), .B(n473), .ZN(n426) );
  XNOR2_X1 U461 ( .A(n424), .B(n739), .ZN(n361) );
  BUF_X1 U462 ( .A(n713), .Z(n717) );
  NAND2_X1 U463 ( .A1(n710), .A2(n741), .ZN(n430) );
  XNOR2_X1 U464 ( .A(n423), .B(KEYINPUT117), .ZN(n749) );
  NAND2_X1 U465 ( .A1(n373), .A2(n412), .ZN(n423) );
  AND2_X1 U466 ( .A1(n374), .A2(n350), .ZN(n373) );
  NAND2_X1 U467 ( .A1(n411), .A2(n414), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n363), .B(KEYINPUT34), .ZN(n525) );
  INV_X1 U469 ( .A(n576), .ZN(n577) );
  AND2_X1 U470 ( .A1(n565), .A2(n586), .ZN(n662) );
  NOR2_X1 U471 ( .A1(n536), .A2(n367), .ZN(n538) );
  XNOR2_X1 U472 ( .A(n428), .B(n427), .ZN(G75) );
  INV_X1 U473 ( .A(KEYINPUT53), .ZN(n427) );
  NAND2_X1 U474 ( .A1(n711), .A2(n429), .ZN(n428) );
  NOR2_X1 U475 ( .A1(n712), .A2(n430), .ZN(n429) );
  AND2_X1 U476 ( .A1(n563), .A2(n349), .ZN(n347) );
  XNOR2_X1 U477 ( .A(n571), .B(n409), .ZN(n555) );
  INV_X1 U478 ( .A(n555), .ZN(n370) );
  AND2_X1 U479 ( .A1(n748), .A2(n528), .ZN(n348) );
  AND2_X1 U480 ( .A1(n674), .A2(n399), .ZN(n349) );
  AND2_X1 U481 ( .A1(n559), .A2(n413), .ZN(n350) );
  AND2_X1 U482 ( .A1(n605), .A2(n606), .ZN(n351) );
  NOR2_X1 U483 ( .A1(n679), .A2(n674), .ZN(n352) );
  AND2_X1 U484 ( .A1(n417), .A2(n545), .ZN(n353) );
  XOR2_X1 U485 ( .A(KEYINPUT65), .B(KEYINPUT22), .Z(n354) );
  XOR2_X1 U486 ( .A(KEYINPUT115), .B(KEYINPUT30), .Z(n355) );
  XOR2_X1 U487 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n356) );
  XOR2_X1 U488 ( .A(n622), .B(n621), .Z(n357) );
  NAND2_X1 U489 ( .A1(n612), .A2(n613), .ZN(n358) );
  XNOR2_X1 U490 ( .A(n401), .B(n355), .ZN(n400) );
  XNOR2_X1 U491 ( .A(n396), .B(n489), .ZN(n402) );
  XNOR2_X1 U492 ( .A(n378), .B(n619), .ZN(n377) );
  NAND2_X1 U493 ( .A1(n359), .A2(n353), .ZN(n416) );
  XNOR2_X1 U494 ( .A(n522), .B(n521), .ZN(n359) );
  INV_X1 U495 ( .A(n725), .ZN(n620) );
  NOR2_X2 U496 ( .A1(n520), .A2(n370), .ZN(n530) );
  NOR2_X1 U497 ( .A1(n749), .A2(n568), .ZN(n393) );
  NAND2_X1 U498 ( .A1(n376), .A2(n408), .ZN(n362) );
  NAND2_X1 U499 ( .A1(n537), .A2(n709), .ZN(n363) );
  NAND2_X1 U500 ( .A1(n578), .A2(n577), .ZN(n628) );
  XNOR2_X1 U501 ( .A(n420), .B(n728), .ZN(n366) );
  NOR2_X1 U502 ( .A1(n633), .A2(n721), .ZN(n634) );
  NOR2_X1 U503 ( .A1(n640), .A2(n721), .ZN(n642) );
  XNOR2_X2 U504 ( .A(n737), .B(G101), .ZN(n490) );
  XNOR2_X2 U505 ( .A(n464), .B(KEYINPUT4), .ZN(n737) );
  XNOR2_X2 U506 ( .A(G143), .B(G128), .ZN(n464) );
  INV_X1 U507 ( .A(n563), .ZN(n367) );
  XNOR2_X2 U508 ( .A(n563), .B(n368), .ZN(n679) );
  XNOR2_X2 U509 ( .A(n501), .B(G469), .ZN(n563) );
  NAND2_X1 U510 ( .A1(n371), .A2(n370), .ZN(n369) );
  XNOR2_X1 U511 ( .A(n532), .B(n372), .ZN(n371) );
  NAND2_X1 U512 ( .A1(n599), .A2(KEYINPUT36), .ZN(n374) );
  NAND2_X1 U513 ( .A1(n618), .A2(KEYINPUT2), .ZN(n378) );
  NAND2_X1 U514 ( .A1(n386), .A2(n351), .ZN(n385) );
  XNOR2_X2 U515 ( .A(n477), .B(n389), .ZN(n739) );
  XNOR2_X1 U516 ( .A(n392), .B(KEYINPUT69), .ZN(n596) );
  NAND2_X1 U517 ( .A1(n394), .A2(n393), .ZN(n392) );
  XNOR2_X1 U518 ( .A(n395), .B(n582), .ZN(n394) );
  NAND2_X1 U519 ( .A1(n580), .A2(n581), .ZN(n395) );
  XNOR2_X1 U520 ( .A(n419), .B(n396), .ZN(n728) );
  NAND2_X1 U521 ( .A1(n707), .A2(n397), .ZN(n711) );
  XNOR2_X2 U522 ( .A(n398), .B(KEYINPUT75), .ZN(n588) );
  NOR2_X2 U523 ( .A1(n571), .A2(n570), .ZN(n401) );
  XNOR2_X1 U524 ( .A(n493), .B(n402), .ZN(n491) );
  NAND2_X1 U525 ( .A1(n416), .A2(n415), .ZN(n546) );
  OR2_X2 U526 ( .A1(n645), .A2(G902), .ZN(n501) );
  NAND2_X1 U527 ( .A1(n617), .A2(n358), .ZN(n407) );
  XNOR2_X1 U528 ( .A(n704), .B(n608), .ZN(n408) );
  XNOR2_X2 U529 ( .A(n410), .B(n492), .ZN(n571) );
  OR2_X2 U530 ( .A1(n622), .A2(G902), .ZN(n410) );
  INV_X1 U531 ( .A(n599), .ZN(n411) );
  NAND2_X1 U532 ( .A1(n558), .A2(KEYINPUT36), .ZN(n413) );
  NAND2_X1 U533 ( .A1(n348), .A2(n545), .ZN(n415) );
  INV_X1 U534 ( .A(n748), .ZN(n417) );
  NAND2_X1 U535 ( .A1(n530), .A2(n352), .ZN(n517) );
  NAND2_X1 U536 ( .A1(n524), .A2(n485), .ZN(n418) );
  XNOR2_X1 U537 ( .A(n421), .B(n438), .ZN(n420) );
  XNOR2_X1 U538 ( .A(n437), .B(n422), .ZN(n421) );
  INV_X1 U539 ( .A(n477), .ZN(n422) );
  BUF_X1 U540 ( .A(n704), .Z(n740) );
  XOR2_X1 U541 ( .A(n593), .B(KEYINPUT64), .Z(n431) );
  INV_X1 U542 ( .A(KEYINPUT74), .ZN(n608) );
  INV_X1 U543 ( .A(KEYINPUT91), .ZN(n446) );
  INV_X1 U544 ( .A(KEYINPUT41), .ZN(n584) );
  INV_X1 U545 ( .A(KEYINPUT116), .ZN(n574) );
  INV_X1 U546 ( .A(n721), .ZN(n625) );
  NAND2_X1 U547 ( .A1(n708), .A2(n586), .ZN(n587) );
  XNOR2_X1 U548 ( .A(n575), .B(n574), .ZN(n578) );
  XOR2_X2 U549 ( .A(G146), .B(G125), .Z(n477) );
  XOR2_X1 U550 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n434) );
  INV_X2 U551 ( .A(G953), .ZN(n741) );
  NAND2_X1 U552 ( .A1(G224), .A2(n741), .ZN(n433) );
  XNOR2_X1 U553 ( .A(n434), .B(n433), .ZN(n438) );
  XNOR2_X1 U554 ( .A(n439), .B(G107), .ZN(n729) );
  XNOR2_X1 U555 ( .A(n729), .B(KEYINPUT71), .ZN(n440) );
  INV_X1 U556 ( .A(n500), .ZN(n441) );
  NAND2_X1 U557 ( .A1(n637), .A2(n614), .ZN(n444) );
  NAND2_X1 U558 ( .A1(n478), .A2(n442), .ZN(n445) );
  AND2_X1 U559 ( .A1(n445), .A2(G210), .ZN(n443) );
  NAND2_X1 U560 ( .A1(n445), .A2(G214), .ZN(n691) );
  NAND2_X1 U561 ( .A1(n573), .A2(n691), .ZN(n447) );
  XNOR2_X2 U562 ( .A(n447), .B(n446), .ZN(n558) );
  INV_X1 U563 ( .A(KEYINPUT19), .ZN(n448) );
  XNOR2_X1 U564 ( .A(n449), .B(KEYINPUT14), .ZN(n450) );
  NAND2_X1 U565 ( .A1(G952), .A2(n450), .ZN(n703) );
  NOR2_X1 U566 ( .A1(G953), .A2(n703), .ZN(n550) );
  NAND2_X1 U567 ( .A1(G902), .A2(n450), .ZN(n547) );
  XOR2_X1 U568 ( .A(G898), .B(KEYINPUT96), .Z(n724) );
  NAND2_X1 U569 ( .A1(G953), .A2(n724), .ZN(n731) );
  NOR2_X1 U570 ( .A1(n547), .A2(n731), .ZN(n451) );
  XOR2_X1 U571 ( .A(KEYINPUT97), .B(n451), .Z(n452) );
  NOR2_X1 U572 ( .A1(n550), .A2(n452), .ZN(n453) );
  XNOR2_X1 U573 ( .A(n453), .B(KEYINPUT98), .ZN(n454) );
  XNOR2_X1 U574 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U575 ( .A(KEYINPUT9), .B(KEYINPUT111), .ZN(n458) );
  XNOR2_X1 U576 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U577 ( .A(n461), .B(n460), .Z(n463) );
  NAND2_X1 U578 ( .A1(G217), .A2(n508), .ZN(n462) );
  XNOR2_X1 U579 ( .A(n463), .B(n462), .ZN(n466) );
  XNOR2_X1 U580 ( .A(n464), .B(KEYINPUT7), .ZN(n465) );
  XNOR2_X1 U581 ( .A(n466), .B(n465), .ZN(n715) );
  NAND2_X1 U582 ( .A1(n715), .A2(n478), .ZN(n467) );
  XNOR2_X1 U583 ( .A(n467), .B(G478), .ZN(n542) );
  INV_X1 U584 ( .A(n542), .ZN(n523) );
  NAND2_X1 U585 ( .A1(n487), .A2(G214), .ZN(n468) );
  XNOR2_X1 U586 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U587 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U588 ( .A1(n630), .A2(n478), .ZN(n480) );
  XNOR2_X1 U589 ( .A(KEYINPUT13), .B(G475), .ZN(n479) );
  XNOR2_X1 U590 ( .A(n480), .B(n479), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n523), .A2(n539), .ZN(n694) );
  NAND2_X1 U592 ( .A1(n614), .A2(G234), .ZN(n481) );
  XNOR2_X1 U593 ( .A(n481), .B(KEYINPUT20), .ZN(n509) );
  NAND2_X1 U594 ( .A1(G221), .A2(n509), .ZN(n483) );
  INV_X1 U595 ( .A(KEYINPUT21), .ZN(n482) );
  XNOR2_X1 U596 ( .A(n483), .B(n482), .ZN(n673) );
  NAND2_X1 U597 ( .A1(n487), .A2(G210), .ZN(n488) );
  XNOR2_X1 U598 ( .A(n488), .B(KEYINPUT5), .ZN(n489) );
  XNOR2_X1 U599 ( .A(n491), .B(n490), .ZN(n622) );
  INV_X1 U600 ( .A(G472), .ZN(n492) );
  INV_X1 U601 ( .A(n493), .ZN(n498) );
  NAND2_X1 U602 ( .A1(n741), .A2(G227), .ZN(n494) );
  XNOR2_X1 U603 ( .A(n494), .B(G104), .ZN(n496) );
  XNOR2_X1 U604 ( .A(KEYINPUT77), .B(G140), .ZN(n495) );
  XNOR2_X1 U605 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U606 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U607 ( .A(n500), .B(n499), .ZN(n645) );
  XNOR2_X1 U608 ( .A(n503), .B(n502), .ZN(n507) );
  XNOR2_X1 U609 ( .A(n505), .B(n504), .ZN(n506) );
  NAND2_X1 U610 ( .A1(n509), .A2(G217), .ZN(n513) );
  XNOR2_X1 U611 ( .A(KEYINPUT101), .B(KEYINPUT25), .ZN(n511) );
  INV_X1 U612 ( .A(KEYINPUT76), .ZN(n510) );
  XNOR2_X1 U613 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X2 U614 ( .A(n515), .B(n514), .ZN(n674) );
  INV_X1 U615 ( .A(KEYINPUT32), .ZN(n516) );
  XNOR2_X1 U616 ( .A(n517), .B(n516), .ZN(n751) );
  INV_X1 U617 ( .A(n676), .ZN(n531) );
  NOR2_X1 U618 ( .A1(n674), .A2(n531), .ZN(n518) );
  NAND2_X1 U619 ( .A1(n679), .A2(n518), .ZN(n519) );
  NOR2_X1 U620 ( .A1(n520), .A2(n519), .ZN(n656) );
  INV_X1 U621 ( .A(KEYINPUT44), .ZN(n528) );
  NAND2_X1 U622 ( .A1(n528), .A2(KEYINPUT90), .ZN(n521) );
  OR2_X1 U623 ( .A1(n523), .A2(n539), .ZN(n576) );
  NAND2_X1 U624 ( .A1(n674), .A2(n673), .ZN(n678) );
  XNOR2_X1 U625 ( .A(KEYINPUT85), .B(KEYINPUT35), .ZN(n526) );
  XNOR2_X1 U626 ( .A(n527), .B(n526), .ZN(n748) );
  AND2_X1 U627 ( .A1(n679), .A2(n674), .ZN(n529) );
  AND2_X1 U628 ( .A1(n530), .A2(n529), .ZN(n649) );
  NAND2_X1 U629 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U630 ( .A(KEYINPUT102), .B(n533), .Z(n685) );
  NAND2_X1 U631 ( .A1(n524), .A2(n685), .ZN(n534) );
  XOR2_X1 U632 ( .A(KEYINPUT31), .B(n534), .Z(n667) );
  INV_X1 U633 ( .A(n678), .ZN(n535) );
  NAND2_X1 U634 ( .A1(n535), .A2(n676), .ZN(n536) );
  NAND2_X1 U635 ( .A1(n538), .A2(n537), .ZN(n652) );
  NAND2_X1 U636 ( .A1(n667), .A2(n652), .ZN(n543) );
  XNOR2_X1 U637 ( .A(n539), .B(KEYINPUT108), .ZN(n541) );
  AND2_X1 U638 ( .A1(n541), .A2(n542), .ZN(n540) );
  XNOR2_X1 U639 ( .A(n540), .B(KEYINPUT112), .ZN(n658) );
  OR2_X1 U640 ( .A1(n658), .A2(n661), .ZN(n690) );
  AND2_X1 U641 ( .A1(n543), .A2(n690), .ZN(n544) );
  XNOR2_X2 U642 ( .A(n546), .B(KEYINPUT45), .ZN(n725) );
  OR2_X1 U643 ( .A1(n741), .A2(n547), .ZN(n548) );
  NOR2_X1 U644 ( .A1(G900), .A2(n548), .ZN(n549) );
  NOR2_X1 U645 ( .A1(n550), .A2(n549), .ZN(n552) );
  INV_X1 U646 ( .A(KEYINPUT80), .ZN(n551) );
  XNOR2_X1 U647 ( .A(n552), .B(n551), .ZN(n553) );
  NAND2_X1 U648 ( .A1(n553), .A2(n673), .ZN(n572) );
  XNOR2_X1 U649 ( .A(n554), .B(KEYINPUT70), .ZN(n561) );
  NOR2_X1 U650 ( .A1(n561), .A2(n555), .ZN(n556) );
  NAND2_X1 U651 ( .A1(n556), .A2(n661), .ZN(n557) );
  INV_X1 U652 ( .A(n679), .ZN(n559) );
  INV_X1 U653 ( .A(n560), .ZN(n565) );
  XNOR2_X1 U654 ( .A(n562), .B(KEYINPUT28), .ZN(n564) );
  AND2_X1 U655 ( .A1(n564), .A2(n563), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n662), .A2(n690), .ZN(n569) );
  INV_X1 U657 ( .A(KEYINPUT67), .ZN(n566) );
  XNOR2_X1 U658 ( .A(n566), .B(KEYINPUT47), .ZN(n567) );
  NOR2_X1 U659 ( .A1(n569), .A2(n567), .ZN(n568) );
  NAND2_X1 U660 ( .A1(n569), .A2(KEYINPUT47), .ZN(n581) );
  INV_X1 U661 ( .A(n691), .ZN(n570) );
  NAND2_X1 U662 ( .A1(n588), .A2(n602), .ZN(n575) );
  INV_X1 U663 ( .A(KEYINPUT83), .ZN(n579) );
  XNOR2_X1 U664 ( .A(n628), .B(n579), .ZN(n580) );
  INV_X1 U665 ( .A(KEYINPUT82), .ZN(n582) );
  INV_X1 U666 ( .A(KEYINPUT38), .ZN(n583) );
  NAND2_X1 U667 ( .A1(n692), .A2(n691), .ZN(n688) );
  NAND2_X1 U668 ( .A1(n588), .A2(n692), .ZN(n591) );
  XNOR2_X1 U669 ( .A(KEYINPUT39), .B(KEYINPUT72), .ZN(n589) );
  XOR2_X1 U670 ( .A(n589), .B(KEYINPUT89), .Z(n590) );
  XNOR2_X1 U671 ( .A(n591), .B(n590), .ZN(n607) );
  NAND2_X1 U672 ( .A1(n607), .A2(n661), .ZN(n592) );
  XNOR2_X1 U673 ( .A(n592), .B(KEYINPUT40), .ZN(n754) );
  NAND2_X1 U674 ( .A1(n753), .A2(n754), .ZN(n594) );
  XNOR2_X1 U675 ( .A(KEYINPUT46), .B(KEYINPUT88), .ZN(n593) );
  XNOR2_X1 U676 ( .A(n594), .B(n431), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U678 ( .A1(n679), .A2(n691), .ZN(n598) );
  NOR2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n601) );
  INV_X1 U680 ( .A(KEYINPUT43), .ZN(n600) );
  XNOR2_X1 U681 ( .A(n601), .B(n600), .ZN(n604) );
  INV_X1 U682 ( .A(n602), .ZN(n603) );
  AND2_X1 U683 ( .A1(n604), .A2(n603), .ZN(n671) );
  INV_X1 U684 ( .A(n671), .ZN(n605) );
  INV_X1 U685 ( .A(KEYINPUT86), .ZN(n606) );
  AND2_X1 U686 ( .A1(n607), .A2(n658), .ZN(n670) );
  NAND2_X1 U687 ( .A1(KEYINPUT2), .A2(KEYINPUT66), .ZN(n612) );
  INV_X1 U688 ( .A(KEYINPUT2), .ZN(n609) );
  OR2_X1 U689 ( .A1(n614), .A2(n609), .ZN(n611) );
  INV_X1 U690 ( .A(KEYINPUT66), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n613) );
  INV_X1 U692 ( .A(n613), .ZN(n616) );
  INV_X1 U693 ( .A(n614), .ZN(n615) );
  OR2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  INV_X1 U695 ( .A(n704), .ZN(n618) );
  INV_X1 U696 ( .A(KEYINPUT84), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n713), .A2(G472), .ZN(n623) );
  XNOR2_X1 U698 ( .A(KEYINPUT118), .B(KEYINPUT62), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n623), .B(n357), .ZN(n626) );
  INV_X1 U700 ( .A(G952), .ZN(n624) );
  AND2_X1 U701 ( .A1(n624), .A2(G953), .ZN(n721) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n627), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U704 ( .A(n628), .B(G143), .ZN(G45) );
  NAND2_X1 U705 ( .A1(n713), .A2(G475), .ZN(n632) );
  XOR2_X1 U706 ( .A(KEYINPUT93), .B(KEYINPUT59), .Z(n629) );
  XNOR2_X1 U707 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n634), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U709 ( .A1(n713), .A2(G210), .ZN(n639) );
  XNOR2_X1 U710 ( .A(KEYINPUT92), .B(KEYINPUT54), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(KEYINPUT55), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U713 ( .A(n639), .B(n638), .ZN(n640) );
  XOR2_X1 U714 ( .A(KEYINPUT87), .B(KEYINPUT56), .Z(n641) );
  XNOR2_X1 U715 ( .A(n642), .B(n641), .ZN(G51) );
  NAND2_X1 U716 ( .A1(n717), .A2(G469), .ZN(n647) );
  XNOR2_X1 U717 ( .A(KEYINPUT125), .B(KEYINPUT57), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n643), .B(KEYINPUT58), .ZN(n644) );
  XNOR2_X1 U719 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X1 U721 ( .A1(n648), .A2(n721), .ZN(G54) );
  XOR2_X1 U722 ( .A(G101), .B(n649), .Z(G3) );
  INV_X1 U723 ( .A(n661), .ZN(n665) );
  NOR2_X1 U724 ( .A1(n665), .A2(n652), .ZN(n651) );
  XNOR2_X1 U725 ( .A(G104), .B(KEYINPUT119), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n651), .B(n650), .ZN(G6) );
  INV_X1 U727 ( .A(n658), .ZN(n668) );
  NOR2_X1 U728 ( .A1(n668), .A2(n652), .ZN(n654) );
  XNOR2_X1 U729 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U731 ( .A(G107), .B(n655), .ZN(G9) );
  XOR2_X1 U732 ( .A(G110), .B(n656), .Z(n657) );
  XNOR2_X1 U733 ( .A(KEYINPUT120), .B(n657), .ZN(G12) );
  XOR2_X1 U734 ( .A(G128), .B(KEYINPUT29), .Z(n660) );
  NAND2_X1 U735 ( .A1(n662), .A2(n658), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n660), .B(n659), .ZN(G30) );
  XOR2_X1 U737 ( .A(G146), .B(KEYINPUT121), .Z(n664) );
  NAND2_X1 U738 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n664), .B(n663), .ZN(G48) );
  NOR2_X1 U740 ( .A1(n665), .A2(n667), .ZN(n666) );
  XOR2_X1 U741 ( .A(G113), .B(n666), .Z(G15) );
  NOR2_X1 U742 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U743 ( .A(G116), .B(n669), .Z(G18) );
  XOR2_X1 U744 ( .A(G134), .B(n670), .Z(G36) );
  XOR2_X1 U745 ( .A(G140), .B(n671), .Z(n672) );
  XNOR2_X1 U746 ( .A(KEYINPUT122), .B(n672), .ZN(G42) );
  NOR2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n675), .B(KEYINPUT49), .ZN(n677) );
  AND2_X1 U749 ( .A1(n677), .A2(n676), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n680), .B(KEYINPUT50), .ZN(n681) );
  AND2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U753 ( .A(KEYINPUT123), .B(n683), .Z(n684) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U755 ( .A(n686), .B(KEYINPUT51), .ZN(n687) );
  NAND2_X1 U756 ( .A1(n687), .A2(n708), .ZN(n700) );
  INV_X1 U757 ( .A(n688), .ZN(n689) );
  NAND2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n697) );
  NOR2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U761 ( .A(KEYINPUT124), .B(n695), .Z(n696) );
  NAND2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U763 ( .A1(n698), .A2(n709), .ZN(n699) );
  NAND2_X1 U764 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U765 ( .A(KEYINPUT52), .B(n701), .Z(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n712) );
  NOR2_X1 U767 ( .A1(n725), .A2(n740), .ZN(n705) );
  NOR2_X1 U768 ( .A1(n705), .A2(KEYINPUT2), .ZN(n706) );
  XNOR2_X1 U769 ( .A(n706), .B(KEYINPUT81), .ZN(n707) );
  NAND2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U771 ( .A1(n713), .A2(G478), .ZN(n714) );
  XOR2_X1 U772 ( .A(n715), .B(n714), .Z(n716) );
  NOR2_X1 U773 ( .A1(n721), .A2(n716), .ZN(G63) );
  NAND2_X1 U774 ( .A1(n717), .A2(G217), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U776 ( .A1(n721), .A2(n720), .ZN(G66) );
  NAND2_X1 U777 ( .A1(G953), .A2(G224), .ZN(n722) );
  XOR2_X1 U778 ( .A(KEYINPUT61), .B(n722), .Z(n723) );
  NOR2_X1 U779 ( .A1(n724), .A2(n723), .ZN(n727) );
  NOR2_X1 U780 ( .A1(G953), .A2(n725), .ZN(n726) );
  NOR2_X1 U781 ( .A1(n727), .A2(n726), .ZN(n734) );
  XNOR2_X1 U782 ( .A(G101), .B(n728), .ZN(n730) );
  XNOR2_X1 U783 ( .A(n730), .B(n729), .ZN(n732) );
  NAND2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U786 ( .A(KEYINPUT126), .B(n735), .ZN(G69) );
  XNOR2_X1 U787 ( .A(n737), .B(n736), .ZN(n738) );
  XNOR2_X1 U788 ( .A(n739), .B(n738), .ZN(n743) );
  XNOR2_X1 U789 ( .A(n740), .B(n743), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n742), .A2(n741), .ZN(n747) );
  XNOR2_X1 U791 ( .A(n743), .B(G227), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n744), .A2(G900), .ZN(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(G953), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n747), .A2(n746), .ZN(G72) );
  XOR2_X1 U795 ( .A(n748), .B(G122), .Z(G24) );
  XNOR2_X1 U796 ( .A(G125), .B(n749), .ZN(n750) );
  XNOR2_X1 U797 ( .A(n750), .B(KEYINPUT37), .ZN(G27) );
  BUF_X1 U798 ( .A(n751), .Z(n752) );
  XOR2_X1 U799 ( .A(G119), .B(n752), .Z(G21) );
  XNOR2_X1 U800 ( .A(G137), .B(n753), .ZN(G39) );
  XOR2_X1 U801 ( .A(G131), .B(n754), .Z(n755) );
  XNOR2_X1 U802 ( .A(KEYINPUT127), .B(n755), .ZN(G33) );
endmodule

