//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND2_X1   g0009(.A1(KEYINPUT64), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(KEYINPUT64), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n215), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n206), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n209), .B(new_n220), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n242), .B(KEYINPUT65), .Z(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G97), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G1), .A3(G13), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n251));
  AND3_X1   g0051(.A1(new_n249), .A2(G238), .A3(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G226), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n222), .A2(G1698), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n255), .B(new_n256), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G97), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n249), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n252), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT13), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT66), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G41), .A2(G45), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(G1), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n250), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  INV_X1    g0070(.A(new_n213), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(new_n248), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n269), .A2(KEYINPUT67), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(KEYINPUT67), .B1(new_n269), .B2(new_n272), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n263), .B(new_n264), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT66), .B1(new_n279), .B2(new_n250), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n266), .A2(new_n265), .A3(G1), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n272), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n269), .A2(KEYINPUT67), .A3(new_n272), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n264), .B1(new_n286), .B2(new_n263), .ZN(new_n287));
  OAI21_X1  g0087(.A(G169), .B1(new_n276), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n276), .A2(new_n287), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n288), .A2(KEYINPUT14), .B1(new_n289), .B2(G179), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n263), .B1(new_n273), .B2(new_n274), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT13), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n291), .B1(new_n293), .B2(new_n275), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT74), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT14), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n295), .B1(new_n294), .B2(new_n296), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n290), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n213), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n212), .A2(G33), .ZN(new_n302));
  INV_X1    g0102(.A(G77), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G20), .ZN(new_n305));
  INV_X1    g0105(.A(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n307), .A2(new_n202), .B1(new_n305), .B2(G68), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n301), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT11), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT71), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n250), .A2(KEYINPUT71), .A3(G13), .A4(G20), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n301), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n250), .A2(G20), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G68), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n311), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n314), .A2(new_n315), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT12), .B1(new_n320), .B2(G68), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n305), .A2(KEYINPUT12), .A3(G68), .ZN(new_n322));
  INV_X1    g0122(.A(G13), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(G1), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n309), .B2(new_n310), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n299), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n293), .A2(G190), .A3(new_n275), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n328), .B(new_n331), .C1(new_n289), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n301), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT8), .B(G58), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(G33), .A3(new_n212), .ZN(new_n338));
  INV_X1    g0138(.A(new_n307), .ZN(new_n339));
  AOI22_X1  g0139(.A1(G150), .A2(new_n339), .B1(new_n203), .B2(G20), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n335), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT9), .ZN(new_n343));
  INV_X1    g0143(.A(new_n312), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n202), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT68), .ZN(new_n346));
  INV_X1    g0146(.A(new_n317), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n202), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n344), .A2(new_n301), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n317), .A2(KEYINPUT68), .A3(G50), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n342), .A2(new_n343), .A3(new_n345), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n345), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT9), .B1(new_n353), .B2(new_n341), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT3), .B(G33), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(G222), .A3(new_n254), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(G223), .A3(G1698), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n357), .B(new_n358), .C1(new_n303), .C2(new_n356), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n262), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n249), .A2(new_n251), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G226), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n286), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G200), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n286), .A2(new_n360), .A3(G190), .A4(new_n362), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n355), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT10), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n355), .A2(KEYINPUT72), .ZN(new_n368));
  XOR2_X1   g0168(.A(KEYINPUT73), .B(KEYINPUT10), .Z(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n352), .A2(new_n370), .A3(new_n354), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n364), .A2(new_n365), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT15), .B(G87), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n302), .A2(new_n375), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n212), .A2(new_n303), .B1(new_n336), .B2(new_n307), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n301), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n316), .A2(G77), .A3(new_n317), .ZN(new_n379));
  INV_X1    g0179(.A(new_n320), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n303), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n257), .A2(new_n258), .ZN(new_n384));
  INV_X1    g0184(.A(G107), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n249), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G232), .A2(G1698), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n254), .A2(G238), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n356), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n386), .A2(new_n389), .B1(new_n361), .B2(G244), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n286), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT70), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n286), .A2(KEYINPUT70), .A3(new_n390), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n383), .B1(new_n395), .B2(new_n332), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n393), .B2(new_n394), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n353), .A2(new_n341), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n363), .B2(new_n291), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT69), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n402), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n363), .A2(G179), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G179), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n395), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n393), .A2(new_n291), .A3(new_n394), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n382), .A3(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n374), .A2(new_n399), .A3(new_n406), .A4(new_n410), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n249), .A2(G232), .A3(new_n251), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n253), .A2(G1698), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(G223), .B2(G1698), .ZN(new_n414));
  INV_X1    g0214(.A(G87), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n414), .A2(new_n384), .B1(new_n306), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n412), .B1(new_n416), .B2(new_n262), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(new_n407), .C1(new_n274), .C2(new_n273), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(G169), .B1(new_n286), .B2(new_n417), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT77), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n336), .B1(new_n250), .B2(G20), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n349), .B1(new_n344), .B2(new_n336), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT75), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G58), .A2(G68), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n305), .B1(new_n217), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G159), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n307), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n424), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(G58), .A2(G68), .ZN(new_n430));
  OAI21_X1  g0230(.A(G20), .B1(new_n430), .B2(new_n201), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(KEYINPUT75), .C1(new_n427), .C2(new_n307), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT7), .B1(new_n356), .B2(G20), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT7), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n212), .A2(new_n384), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n436), .A3(G68), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(KEYINPUT16), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n301), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT64), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n305), .ZN(new_n443));
  NAND2_X1  g0243(.A1(KEYINPUT64), .A2(G20), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT7), .B1(new_n445), .B2(new_n356), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n384), .A2(new_n435), .A3(new_n305), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(G68), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n426), .A2(new_n428), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n441), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n423), .B1(new_n439), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n417), .B1(new_n274), .B2(new_n273), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n291), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT77), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n418), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n421), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT18), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT18), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n421), .A2(new_n458), .A3(new_n455), .A4(new_n451), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n448), .A2(new_n449), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n301), .B(new_n438), .C1(new_n460), .C2(new_n441), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n286), .A2(G190), .A3(new_n417), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n452), .A2(G200), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n461), .A2(new_n423), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT17), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n463), .A2(new_n462), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n467), .A2(KEYINPUT17), .A3(new_n461), .A4(new_n423), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n457), .A2(new_n459), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n334), .A2(new_n411), .A3(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(G244), .B(new_n254), .C1(new_n257), .C2(new_n258), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT4), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G250), .A2(G1698), .ZN(new_n476));
  NAND2_X1  g0276(.A1(KEYINPUT4), .A2(G244), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(G1698), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n356), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT79), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(new_n479), .A3(KEYINPUT79), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n262), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT81), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT80), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(new_n277), .A3(KEYINPUT5), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(KEYINPUT80), .B2(G41), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n278), .A2(G1), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n249), .A2(G274), .ZN(new_n492));
  OR2_X1    g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n249), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n224), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n484), .A2(new_n485), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n485), .B1(new_n484), .B2(new_n496), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n291), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT78), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT6), .ZN(new_n501));
  AND2_X1   g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  NOR2_X1   g0302(.A1(G97), .A2(G107), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n385), .A2(KEYINPUT6), .A3(G97), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n212), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n307), .A2(new_n303), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n507), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n385), .A2(KEYINPUT6), .A3(G97), .ZN(new_n510));
  XNOR2_X1  g0310(.A(G97), .B(G107), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(new_n501), .ZN(new_n512));
  OAI211_X1 g0312(.A(KEYINPUT78), .B(new_n509), .C1(new_n512), .C2(new_n212), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n446), .A2(G107), .A3(new_n447), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n508), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n301), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n312), .A2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n250), .A2(G33), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n335), .A2(new_n312), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n517), .B1(new_n520), .B2(G97), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n249), .B1(new_n480), .B2(new_n481), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n495), .B1(new_n522), .B2(new_n483), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n516), .A2(new_n521), .B1(new_n523), .B2(new_n407), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n499), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n473), .A2(new_n479), .A3(KEYINPUT79), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT79), .B1(new_n473), .B2(new_n479), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n526), .A2(new_n527), .A3(new_n249), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT81), .B1(new_n528), .B2(new_n495), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n484), .A2(new_n485), .A3(new_n496), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(G190), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n516), .A2(new_n521), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n332), .B1(new_n484), .B2(new_n496), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(G238), .B(new_n254), .C1(new_n257), .C2(new_n258), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT82), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT82), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n356), .A2(new_n538), .A3(G238), .A4(new_n254), .ZN(new_n539));
  INV_X1    g0339(.A(G116), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT83), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT83), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G116), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G33), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n356), .A2(G244), .A3(G1698), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n537), .A2(new_n539), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n262), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n250), .A2(G45), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n549), .A2(G250), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n249), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n492), .B2(new_n549), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G200), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n552), .B1(new_n547), .B2(new_n262), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G190), .ZN(new_n557));
  INV_X1    g0357(.A(new_n375), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n320), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n519), .A2(new_n415), .ZN(new_n560));
  OR2_X1    g0360(.A1(KEYINPUT85), .A2(G87), .ZN(new_n561));
  NAND2_X1  g0361(.A1(KEYINPUT85), .A2(G87), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n503), .A3(new_n562), .ZN(new_n563));
  OR2_X1    g0363(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n564));
  NAND2_X1  g0364(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n260), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n563), .B1(new_n566), .B2(new_n445), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n443), .A2(G33), .A3(G97), .A4(new_n444), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n564), .A3(new_n565), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n212), .A2(new_n356), .A3(G68), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI211_X1 g0371(.A(new_n559), .B(new_n560), .C1(new_n571), .C2(new_n301), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n555), .A2(new_n557), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n556), .A2(new_n407), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n301), .ZN(new_n575));
  INV_X1    g0375(.A(new_n559), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n520), .A2(new_n558), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n574), .B(new_n578), .C1(G169), .C2(new_n556), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n525), .A2(new_n535), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n306), .A2(G97), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n443), .A2(new_n582), .A3(new_n444), .A4(new_n474), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n541), .A2(new_n543), .A3(G20), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n301), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(new_n584), .A3(KEYINPUT20), .A4(new_n301), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g0389(.A(KEYINPUT83), .B(G116), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n540), .B1(new_n250), .B2(G33), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n380), .A2(new_n590), .B1(new_n316), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G257), .B(new_n254), .C1(new_n257), .C2(new_n258), .ZN(new_n594));
  OAI211_X1 g0394(.A(G264), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n595));
  INV_X1    g0395(.A(G303), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n594), .B(new_n595), .C1(new_n596), .C2(new_n356), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n262), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n491), .A2(G270), .A3(new_n249), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n493), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(G169), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT86), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT21), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT21), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n593), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n598), .A2(G179), .A3(new_n493), .A4(new_n599), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n600), .A2(G200), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n607), .B(new_n611), .C1(new_n397), .C2(new_n600), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n604), .A2(new_n606), .A3(new_n610), .A4(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n443), .B(new_n444), .C1(new_n257), .C2(new_n258), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT22), .B1(new_n614), .B2(new_n415), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT22), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n212), .A2(new_n356), .A3(new_n616), .A4(G87), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT24), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n590), .A2(G20), .A3(new_n306), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT23), .B1(new_n305), .B2(G107), .ZN(new_n621));
  OR2_X1    g0421(.A1(KEYINPUT23), .A2(G107), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n212), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n618), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n301), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n344), .A2(new_n385), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n628), .B(KEYINPUT25), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(G107), .B2(new_n520), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(G257), .B(G1698), .C1(new_n257), .C2(new_n258), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT87), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n356), .A2(KEYINPUT87), .A3(G257), .A4(G1698), .ZN(new_n635));
  NAND2_X1  g0435(.A1(G33), .A2(G294), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n356), .A2(G250), .A3(new_n254), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n634), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n262), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n491), .A2(G264), .A3(new_n249), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n639), .A2(G179), .A3(new_n493), .A4(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n491), .A2(new_n492), .ZN(new_n642));
  INV_X1    g0442(.A(new_n640), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n642), .B(new_n643), .C1(new_n638), .C2(new_n262), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n641), .B(KEYINPUT88), .C1(new_n644), .C2(new_n291), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT88), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n646), .A3(G179), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n631), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n644), .A2(G200), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n643), .B1(new_n638), .B2(new_n262), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n650), .A2(new_n397), .A3(new_n493), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n627), .B(new_n630), .C1(new_n649), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n581), .A2(new_n613), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n470), .A2(new_n654), .ZN(G372));
  INV_X1    g0455(.A(new_n406), .ZN(new_n656));
  INV_X1    g0456(.A(new_n333), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n410), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n329), .B2(new_n299), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n468), .A2(new_n466), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n457), .B(new_n459), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n656), .B1(new_n661), .B2(new_n374), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n559), .B1(new_n571), .B2(new_n301), .ZN(new_n663));
  INV_X1    g0463(.A(new_n560), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n663), .B(new_n664), .C1(new_n556), .C2(new_n332), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT89), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n555), .A2(KEYINPUT89), .A3(new_n572), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n668), .A3(new_n557), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n525), .A2(new_n535), .A3(new_n669), .A4(new_n652), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n609), .B1(new_n603), .B2(KEYINPUT21), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n648), .A2(new_n606), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n579), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n573), .A2(new_n579), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n525), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(G169), .B1(new_n529), .B2(new_n530), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n523), .A2(new_n407), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n532), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n579), .A3(new_n669), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n676), .B1(new_n674), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n470), .B1(new_n673), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n662), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT90), .Z(G369));
  NAND2_X1  g0485(.A1(new_n212), .A2(new_n324), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT91), .ZN(new_n688));
  OAI21_X1  g0488(.A(G213), .B1(new_n686), .B2(KEYINPUT27), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n607), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n613), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n671), .A2(new_n606), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n692), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n696), .B(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n648), .A2(new_n691), .ZN(new_n699));
  INV_X1    g0499(.A(new_n691), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n631), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n648), .A2(new_n701), .A3(new_n652), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n698), .A2(G330), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n694), .A2(new_n691), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n706), .A2(new_n653), .B1(new_n648), .B2(new_n700), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n705), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n207), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n250), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n563), .A2(G116), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n711), .A2(new_n712), .B1(new_n219), .B2(new_n710), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT28), .Z(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT26), .B1(new_n680), .B2(new_n580), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n557), .B1(new_n665), .B2(new_n666), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT89), .B1(new_n555), .B2(new_n572), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n579), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n525), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n715), .B1(KEYINPUT26), .B2(new_n719), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT29), .B(new_n691), .C1(new_n720), .C2(new_n673), .ZN(new_n721));
  INV_X1    g0521(.A(new_n579), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n497), .A2(new_n498), .A3(new_n397), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n516), .B(new_n521), .C1(new_n523), .C2(new_n332), .ZN(new_n724));
  OAI22_X1  g0524(.A1(new_n723), .A2(new_n724), .B1(new_n677), .B2(new_n679), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n669), .A2(new_n652), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n648), .A2(new_n671), .A3(new_n606), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n722), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n680), .A2(KEYINPUT26), .A3(new_n580), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n719), .B2(KEYINPUT26), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n700), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n721), .B1(new_n732), .B2(KEYINPUT29), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  INV_X1    g0534(.A(new_n608), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n529), .A2(new_n530), .A3(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n556), .A2(new_n650), .A3(KEYINPUT93), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT93), .B1(new_n556), .B2(new_n650), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n734), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n497), .A2(new_n498), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n556), .A2(new_n650), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT93), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n556), .A2(new_n650), .A3(KEYINPUT93), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n741), .A2(new_n746), .A3(KEYINPUT30), .A4(new_n735), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT94), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n644), .B1(new_n748), .B2(new_n554), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n600), .A2(new_n407), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n523), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n749), .B(new_n751), .C1(new_n748), .C2(new_n554), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n740), .A2(new_n747), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n700), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT31), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n653), .A2(new_n613), .ZN(new_n758));
  INV_X1    g0558(.A(new_n725), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n758), .A2(new_n759), .A3(new_n580), .A4(new_n691), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n756), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G330), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n733), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT95), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n733), .A2(KEYINPUT95), .A3(new_n762), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n714), .B1(new_n767), .B2(G1), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT96), .Z(G364));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n213), .B1(G20), .B2(new_n291), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n356), .A2(new_n207), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT97), .ZN(new_n776));
  INV_X1    g0576(.A(G355), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n776), .A2(new_n777), .B1(G116), .B2(new_n207), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n709), .A2(new_n356), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G45), .B2(new_n218), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n242), .B2(G45), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n774), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n445), .A2(new_n323), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G45), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n711), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n212), .A2(new_n407), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G190), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G311), .ZN(new_n791));
  INV_X1    g0591(.A(G283), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n332), .A2(G179), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n445), .A2(new_n397), .A3(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n790), .A2(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G179), .A2(G200), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n445), .A2(new_n397), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n795), .B1(G329), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n793), .A2(G20), .A3(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n356), .B1(new_n801), .B2(G303), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n796), .A2(G190), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n445), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n788), .A2(G190), .A3(new_n332), .ZN(new_n807));
  INV_X1    g0607(.A(G322), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n802), .B1(new_n805), .B2(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n788), .A2(G200), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n397), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(KEYINPUT100), .B(KEYINPUT33), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(G317), .Z(new_n815));
  AOI21_X1  g0615(.A(new_n809), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n811), .A2(G190), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT99), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G326), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n799), .B(new_n816), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT101), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n817), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G50), .A2(new_n824), .B1(new_n813), .B2(G68), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n797), .A2(new_n427), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT32), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n807), .B(KEYINPUT98), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G58), .ZN(new_n829));
  INV_X1    g0629(.A(new_n794), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G107), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n804), .A2(G97), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n561), .A2(new_n562), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n384), .B1(new_n801), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n790), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(G77), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n825), .A2(new_n827), .A3(new_n829), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n821), .A2(new_n822), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n823), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n787), .B1(new_n840), .B2(new_n773), .ZN(new_n841));
  INV_X1    g0641(.A(new_n772), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n696), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n698), .A2(G330), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n785), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n698), .A2(G330), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT102), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  NOR2_X1   g0649(.A1(new_n410), .A2(new_n700), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n396), .A2(new_n398), .B1(new_n383), .B2(new_n691), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n410), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n732), .B(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(new_n762), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT105), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n786), .B1(new_n853), .B2(new_n762), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n773), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n771), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n786), .B1(G77), .B2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n824), .A2(G137), .B1(new_n836), .B2(G159), .ZN(new_n861));
  INV_X1    g0661(.A(G150), .ZN(new_n862));
  INV_X1    g0662(.A(G143), .ZN(new_n863));
  INV_X1    g0663(.A(new_n828), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n861), .B1(new_n862), .B2(new_n812), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT34), .Z(new_n866));
  NAND2_X1  g0666(.A1(new_n830), .A2(G68), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n798), .A2(G132), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n804), .A2(G58), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n384), .B1(new_n801), .B2(G50), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n832), .B1(new_n807), .B2(new_n806), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT103), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n384), .B1(new_n800), .B2(new_n385), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n790), .A2(new_n590), .B1(new_n415), .B2(new_n794), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n874), .B(new_n875), .C1(G311), .C2(new_n798), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n876), .B1(new_n792), .B2(new_n812), .C1(new_n596), .C2(new_n817), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n866), .A2(new_n871), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n860), .B1(new_n878), .B2(new_n773), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n771), .B2(new_n852), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT104), .Z(new_n881));
  NOR2_X1   g0681(.A1(new_n857), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(G384));
  NOR2_X1   g0683(.A1(new_n783), .A2(new_n250), .ZN(new_n884));
  INV_X1    g0684(.A(G330), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT107), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n328), .A2(new_n691), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n293), .A2(G179), .A3(new_n275), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n294), .B2(new_n296), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT74), .B1(new_n288), .B2(KEYINPUT14), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n333), .B(new_n888), .C1(new_n893), .C2(new_n328), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n290), .B(new_n333), .C1(new_n297), .C2(new_n298), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(KEYINPUT106), .A3(new_n887), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT106), .B1(new_n895), .B2(new_n887), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n886), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n898), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n900), .A2(KEYINPUT107), .A3(new_n894), .A4(new_n896), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n852), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n654), .A2(new_n691), .B1(new_n754), .B2(new_n755), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n904), .B2(new_n757), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT112), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT112), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n902), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n441), .B1(new_n433), .B2(new_n437), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n423), .B1(new_n439), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n421), .A2(new_n455), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n690), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n464), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT37), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT109), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(KEYINPUT110), .B(KEYINPUT37), .Z(new_n919));
  NAND2_X1  g0719(.A1(new_n451), .A2(new_n690), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n456), .A2(new_n464), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(KEYINPUT109), .B(KEYINPUT37), .C1(new_n913), .C2(new_n915), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n918), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n914), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n469), .A2(KEYINPUT108), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT108), .B1(new_n469), .B2(new_n924), .ZN(new_n926));
  OAI211_X1 g0726(.A(KEYINPUT38), .B(new_n923), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n456), .A2(new_n464), .A3(new_n920), .ZN(new_n928));
  INV_X1    g0728(.A(new_n919), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n921), .ZN(new_n931));
  INV_X1    g0731(.A(new_n469), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n931), .B1(new_n932), .B2(new_n920), .ZN(new_n933));
  XNOR2_X1  g0733(.A(KEYINPUT111), .B(KEYINPUT38), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n910), .B1(new_n927), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n907), .A2(new_n909), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n469), .A2(new_n924), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT108), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n469), .A2(KEYINPUT108), .A3(new_n924), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT38), .B1(new_n942), .B2(new_n923), .ZN(new_n943));
  INV_X1    g0743(.A(new_n927), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n910), .B1(new_n945), .B2(new_n906), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n937), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n761), .A2(new_n470), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n885), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n947), .B2(new_n948), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n690), .B1(new_n457), .B2(new_n459), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n691), .B(new_n852), .C1(new_n682), .C2(new_n673), .ZN(new_n952));
  INV_X1    g0752(.A(new_n850), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n902), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT38), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n927), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n951), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(KEYINPUT39), .A3(new_n927), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n927), .A2(new_n935), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT39), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n330), .A2(new_n700), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n961), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n721), .B(new_n470), .C1(new_n732), .C2(KEYINPUT29), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n662), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n968), .B(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n884), .B1(new_n950), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n971), .B2(new_n950), .ZN(new_n973));
  INV_X1    g0773(.A(new_n512), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT35), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(KEYINPUT35), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n975), .A2(G116), .A3(new_n214), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT36), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n219), .A2(G77), .A3(new_n425), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(G50), .B2(new_n216), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(G1), .A3(new_n323), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n973), .A2(new_n978), .A3(new_n981), .ZN(G367));
  INV_X1    g0782(.A(new_n779), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n774), .B1(new_n207), .B2(new_n375), .C1(new_n238), .C2(new_n983), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n984), .A2(new_n786), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n691), .A2(new_n572), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n669), .A2(new_n986), .A3(new_n579), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n579), .B2(new_n986), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n794), .A2(new_n303), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n202), .B2(new_n790), .ZN(new_n991));
  INV_X1    g0791(.A(new_n807), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n991), .B1(G150), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n798), .A2(G137), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n804), .A2(G68), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n384), .B1(new_n801), .B2(G58), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(new_n813), .B2(G159), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n993), .B(new_n998), .C1(new_n819), .C2(new_n863), .ZN(new_n999));
  XOR2_X1   g0799(.A(KEYINPUT113), .B(G311), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n819), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT114), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n794), .A2(new_n223), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n356), .B(new_n1003), .C1(G317), .C2(new_n798), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1001), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n801), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n800), .A2(new_n590), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1007), .B1(new_n1008), .B2(KEYINPUT46), .C1(new_n385), .C2(new_n805), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G283), .B2(new_n836), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n806), .B2(new_n812), .C1(new_n864), .C2(new_n596), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n999), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  OAI221_X1 g0813(.A(new_n985), .B1(new_n842), .B2(new_n988), .C1(new_n1013), .C2(new_n858), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n700), .A2(new_n532), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n759), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n680), .A2(new_n700), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n706), .A2(new_n653), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n525), .B1(new_n1016), .B2(new_n648), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1020), .A2(KEYINPUT42), .B1(new_n1021), .B2(new_n691), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(KEYINPUT42), .B2(new_n1020), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n704), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1027), .B(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n784), .A2(G1), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT45), .ZN(new_n1032));
  OR3_X1    g0832(.A1(new_n1028), .A2(new_n1032), .A3(new_n707), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(new_n1028), .B2(new_n707), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1028), .A2(new_n707), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT44), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1028), .A2(KEYINPUT44), .A3(new_n707), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n705), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1035), .A2(new_n1040), .A3(new_n704), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n706), .A2(new_n699), .A3(new_n702), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n653), .B2(new_n706), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n844), .B(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n767), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n710), .B(KEYINPUT41), .Z(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1031), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1014), .B1(new_n1030), .B2(new_n1051), .ZN(G387));
  AOI21_X1  g0852(.A(new_n1047), .B1(new_n765), .B2(new_n766), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n710), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1047), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n767), .B2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G294), .A2(new_n801), .B1(new_n804), .B2(G283), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n812), .A2(new_n1000), .B1(new_n596), .B2(new_n790), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n819), .A2(new_n808), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(G317), .C2(new_n828), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1058), .B1(new_n1061), .B2(KEYINPUT48), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(KEYINPUT48), .B2(new_n1061), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT49), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n384), .B1(new_n797), .B2(new_n820), .C1(new_n590), .C2(new_n794), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n807), .A2(new_n202), .B1(new_n790), .B2(new_n216), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n805), .A2(new_n375), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n801), .A2(G77), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(new_n356), .A3(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1003), .B(new_n1071), .C1(new_n337), .C2(new_n813), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n427), .B2(new_n817), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1067), .B(new_n1073), .C1(G150), .C2(new_n798), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT116), .Z(new_n1075));
  OAI21_X1  g0875(.A(new_n773), .B1(new_n1066), .B2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n712), .B(KEYINPUT115), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n278), .B1(new_n216), .B2(new_n303), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n336), .A2(G50), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT50), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n1080), .B2(new_n1079), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n779), .B1(new_n1077), .B2(new_n1082), .C1(new_n235), .C2(new_n278), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(G107), .B2(new_n207), .C1(new_n712), .C2(new_n776), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n785), .B1(new_n1084), .B2(new_n774), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1076), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n699), .A2(new_n702), .A3(new_n772), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1086), .A2(new_n1087), .B1(new_n1031), .B2(new_n1056), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1057), .A2(new_n1088), .ZN(G393));
  NAND2_X1  g0889(.A1(new_n246), .A2(new_n779), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n773), .B(new_n772), .C1(G97), .C2(new_n709), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n785), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n790), .A2(new_n336), .B1(new_n863), .B2(new_n797), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n805), .A2(new_n303), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n384), .B(new_n1094), .C1(G68), .C2(new_n801), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n415), .B2(new_n794), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1093), .B(new_n1096), .C1(G50), .C2(new_n813), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n817), .A2(new_n862), .B1(new_n427), .B2(new_n807), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT51), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n824), .A2(G317), .B1(G311), .B2(new_n992), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT52), .Z(new_n1101));
  OAI22_X1  g0901(.A1(new_n790), .A2(new_n806), .B1(new_n808), .B2(new_n797), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n356), .B1(new_n801), .B2(G283), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n831), .B(new_n1103), .C1(new_n590), .C2(new_n805), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1102), .B(new_n1104), .C1(G303), .C2(new_n813), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1097), .A2(new_n1099), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1092), .B1(new_n858), .B2(new_n1106), .C1(new_n1018), .C2(new_n842), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1031), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1107), .B1(new_n1044), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1044), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1110), .A2(new_n1053), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1054), .B1(new_n1110), .B2(new_n1053), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(G390));
  NAND3_X1  g0914(.A1(new_n902), .A2(new_n905), .A3(G330), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n851), .A2(new_n410), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n691), .B(new_n1116), .C1(new_n720), .C2(new_n673), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1117), .A2(new_n953), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n761), .A2(G330), .A3(new_n852), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1119), .A2(new_n899), .A3(new_n901), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1115), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n954), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n761), .A2(new_n470), .A3(G330), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n969), .A2(new_n662), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT117), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT117), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n969), .A2(new_n1128), .A3(new_n662), .A4(new_n1125), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT118), .B1(new_n1124), .B2(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1115), .A2(new_n1120), .A3(new_n1118), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n902), .B(new_n1119), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n1122), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT118), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1131), .A2(KEYINPUT119), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1115), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n966), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n965), .A2(new_n962), .B1(new_n955), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n963), .A2(new_n1140), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n899), .A2(new_n901), .B1(new_n1117), .B2(new_n953), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1139), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n962), .A2(new_n965), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n955), .A2(new_n1140), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n1149), .A3(new_n1115), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1138), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1131), .A2(new_n1137), .A3(new_n1153), .A4(KEYINPUT119), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n710), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1151), .A2(new_n1031), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n786), .B1(new_n337), .B2(new_n859), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n384), .B1(new_n800), .B2(new_n415), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1158), .B(new_n1094), .C1(G68), .C2(new_n830), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n385), .B2(new_n812), .C1(new_n792), .C2(new_n817), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n992), .A2(G116), .B1(new_n836), .B2(G97), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n806), .B2(new_n797), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n813), .A2(G137), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n824), .A2(G128), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n801), .A2(G150), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(KEYINPUT53), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1165), .A2(KEYINPUT53), .B1(G159), .B2(new_n804), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n384), .B1(new_n830), .B2(G50), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1169), .A2(KEYINPUT120), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT54), .B(G143), .Z(new_n1171));
  AOI22_X1  g0971(.A1(new_n992), .A2(G132), .B1(new_n836), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(KEYINPUT120), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n798), .A2(G125), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1170), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1160), .A2(new_n1162), .B1(new_n1168), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1157), .B1(new_n1176), .B2(new_n773), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1146), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1177), .B1(new_n1178), .B2(new_n771), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1156), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1155), .A2(new_n1181), .ZN(G378));
  OAI211_X1 g0982(.A(new_n902), .B(new_n905), .C1(new_n943), .C2(new_n944), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n885), .B1(new_n1183), .B2(new_n910), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n374), .A2(new_n406), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n690), .B1(new_n341), .B2(new_n353), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1187), .B(new_n1188), .Z(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1184), .A2(new_n937), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1184), .B2(new_n937), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n968), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n946), .A2(G330), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n909), .A2(new_n936), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n908), .B1(new_n902), .B2(new_n905), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1189), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n968), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1184), .A2(new_n937), .A3(new_n1190), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1193), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1031), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n786), .B1(G50), .B2(new_n859), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n992), .A2(G128), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n804), .A2(G150), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n801), .A2(new_n1171), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(G125), .ZN(new_n1209));
  INV_X1    g1009(.A(G132), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n1209), .A2(new_n817), .B1(new_n812), .B2(new_n1210), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1208), .B(new_n1211), .C1(G137), .C2(new_n836), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n830), .A2(G159), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n798), .C2(G124), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n812), .A2(new_n223), .B1(new_n375), .B2(new_n790), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT121), .Z(new_n1220));
  OAI21_X1  g1020(.A(new_n995), .B1(new_n817), .B2(new_n540), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT122), .Z(new_n1222));
  NOR2_X1   g1022(.A1(new_n794), .A2(new_n215), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n356), .A2(G41), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1070), .B(new_n1224), .C1(new_n807), .C2(new_n385), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G283), .C2(new_n798), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1220), .A2(new_n1222), .A3(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(KEYINPUT58), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(KEYINPUT58), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1224), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1231), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1218), .A2(new_n1229), .A3(new_n1230), .A4(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1204), .B1(new_n1233), .B2(new_n773), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1190), .B2(new_n771), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1203), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1202), .A2(KEYINPUT57), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1153), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(new_n1130), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n710), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1124), .A2(KEYINPUT118), .A3(new_n1130), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1136), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1151), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1132), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT57), .B1(new_n1244), .B2(new_n1202), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1236), .B1(new_n1240), .B2(new_n1245), .ZN(G375));
  OAI21_X1  g1046(.A(new_n786), .B1(G68), .B2(new_n859), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n992), .A2(G283), .B1(G303), .B2(new_n798), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n385), .B2(new_n790), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n356), .B(new_n1068), .C1(G97), .C2(new_n801), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n824), .A2(G294), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(new_n1251), .A3(new_n990), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1249), .B(new_n1252), .C1(new_n544), .C2(new_n813), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1253), .A2(KEYINPUT123), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(KEYINPUT123), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G132), .A2(new_n824), .B1(new_n813), .B2(new_n1171), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n828), .A2(G137), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n356), .B1(new_n800), .B2(new_n427), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1258), .B(new_n1223), .C1(G50), .C2(new_n804), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n836), .A2(G150), .B1(G128), .B2(new_n798), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1256), .A2(new_n1257), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1254), .A2(new_n1255), .A3(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1247), .B1(new_n1262), .B2(new_n773), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n902), .B2(new_n771), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1124), .B2(new_n1108), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1131), .A2(new_n1137), .A3(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1268), .B2(new_n1049), .ZN(G381));
  INV_X1    g1069(.A(G387), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(G393), .A2(G396), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1270), .A2(new_n1271), .A3(new_n882), .A4(new_n1113), .ZN(new_n1272));
  OR4_X1    g1072(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1272), .ZN(G407));
  INV_X1    g1073(.A(G343), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(G213), .ZN(new_n1275));
  OR3_X1    g1075(.A1(G375), .A2(G378), .A3(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(G407), .A2(G213), .A3(new_n1276), .ZN(G409));
  INV_X1    g1077(.A(KEYINPUT125), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1268), .A2(KEYINPUT60), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n710), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1279), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(G384), .B1(new_n1284), .B2(new_n1266), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1282), .B1(new_n1268), .B2(KEYINPUT60), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1286), .A2(new_n882), .A3(new_n1265), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1278), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1284), .A2(G384), .A3(new_n1266), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n882), .B1(new_n1286), .B2(new_n1265), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1289), .A2(KEYINPUT125), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G378), .B(new_n1236), .C1(new_n1240), .C2(new_n1245), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1054), .B1(new_n1138), .B2(new_n1151), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1180), .B1(new_n1294), .B2(new_n1154), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1202), .B(new_n1050), .C1(new_n1130), .C2(new_n1238), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1235), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1193), .A2(new_n1201), .A3(KEYINPUT124), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1031), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT124), .B1(new_n1193), .B2(new_n1201), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1295), .B1(new_n1297), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1293), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1292), .A2(new_n1303), .A3(new_n1275), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1303), .A2(new_n1275), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1289), .A2(KEYINPUT125), .A3(new_n1290), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT125), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1309));
  INV_X1    g1109(.A(G2897), .ZN(new_n1310));
  OAI22_X1  g1110(.A1(new_n1308), .A2(new_n1309), .B1(new_n1310), .B2(new_n1275), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1275), .A2(new_n1310), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1307), .A2(new_n1311), .A3(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(G393), .B(G396), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(G387), .A2(new_n1113), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(G387), .A2(new_n1113), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1315), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n848), .B1(new_n1057), .B2(new_n1088), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1271), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1270), .A2(G390), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(new_n1322), .A3(new_n1316), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1319), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  AOI22_X1  g1125(.A1(new_n1293), .A2(new_n1302), .B1(G213), .B2(new_n1274), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1305), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1325), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1306), .A2(new_n1314), .A3(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT126), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1306), .A2(new_n1314), .A3(new_n1328), .A4(KEYINPUT126), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT61), .B1(new_n1304), .B2(KEYINPUT62), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT62), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1326), .A2(new_n1335), .A3(new_n1292), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1334), .A2(new_n1314), .A3(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1333), .A2(new_n1339), .ZN(G405));
  NAND2_X1  g1140(.A1(G375), .A2(new_n1295), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1293), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT127), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1341), .A2(KEYINPUT127), .A3(new_n1293), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1344), .A2(new_n1292), .A3(new_n1345), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n1341), .B(new_n1293), .C1(new_n1285), .C2(new_n1287), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  XNOR2_X1  g1148(.A(new_n1348), .B(new_n1338), .ZN(G402));
endmodule


