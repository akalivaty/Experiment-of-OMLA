//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  AND2_X1   g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(G197gat), .B(G204gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n212), .A3(new_n205), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  INV_X1    g021(.A(G155gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT80), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT80), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G155gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n222), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n218), .B(new_n221), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT78), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(new_n228), .ZN(new_n232));
  OR2_X1    g031(.A1(G141gat), .A2(G148gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(G141gat), .A2(G148gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(KEYINPUT79), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT79), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n219), .B2(new_n220), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n232), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n231), .B1(G155gat), .B2(G162gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n217), .A2(KEYINPUT78), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n216), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n229), .B(new_n230), .C1(new_n238), .C2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT29), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n214), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT3), .B1(new_n214), .B2(new_n243), .ZN(new_n245));
  INV_X1    g044(.A(new_n232), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n219), .A2(new_n220), .A3(new_n236), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT79), .B1(new_n233), .B2(new_n234), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n241), .ZN(new_n250));
  INV_X1    g049(.A(new_n217), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n233), .B(new_n234), .C1(new_n251), .C2(new_n215), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT80), .B(G155gat), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT2), .B1(new_n254), .B2(new_n222), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n249), .A2(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n245), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n202), .B1(new_n244), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT88), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g059(.A(KEYINPUT88), .B(new_n202), .C1(new_n244), .C2(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n202), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(new_n245), .B2(new_n256), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n214), .B(KEYINPUT75), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n242), .A2(new_n243), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G22gat), .ZN(new_n270));
  INV_X1    g069(.A(G78gat), .ZN(new_n271));
  INV_X1    g070(.A(G22gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n262), .A2(new_n272), .A3(new_n268), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n272), .B1(new_n262), .B2(new_n268), .ZN(new_n275));
  AOI211_X1 g074(.A(G22gat), .B(new_n267), .C1(new_n260), .C2(new_n261), .ZN(new_n276));
  OAI21_X1  g075(.A(G78gat), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT31), .B(G50gat), .ZN(new_n278));
  INV_X1    g077(.A(G106gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n274), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n280), .B1(new_n274), .B2(new_n277), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n285), .A2(KEYINPUT26), .ZN(new_n286));
  INV_X1    g085(.A(G169gat), .ZN(new_n287));
  INV_X1    g086(.A(G176gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n290));
  AOI211_X1 g089(.A(new_n284), .B(new_n286), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT27), .B(G183gat), .ZN(new_n292));
  INV_X1    g091(.A(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n295), .A2(KEYINPUT65), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(KEYINPUT65), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  OAI22_X1  g098(.A1(new_n299), .A2(KEYINPUT66), .B1(new_n295), .B2(new_n294), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n292), .A2(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n291), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n285), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n284), .A2(new_n309), .B1(G169gat), .B2(G176gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(G183gat), .B(G190gat), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n308), .B(new_n310), .C1(new_n309), .C2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT25), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G183gat), .B(G190gat), .Z(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT24), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n316), .A2(KEYINPUT25), .A3(new_n308), .A4(new_n310), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n304), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n243), .ZN(new_n320));
  NAND2_X1  g119(.A1(G226gat), .A2(G233gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT64), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n314), .A2(new_n323), .A3(new_n317), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n314), .B2(new_n317), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n304), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n321), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(KEYINPUT76), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT76), .B1(new_n326), .B2(new_n327), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n214), .B(new_n322), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n318), .A2(KEYINPUT64), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n323), .A3(new_n317), .ZN(new_n333));
  INV_X1    g132(.A(new_n294), .ZN(new_n334));
  AOI22_X1  g133(.A1(KEYINPUT28), .A2(new_n334), .B1(new_n301), .B2(new_n302), .ZN(new_n335));
  INV_X1    g134(.A(new_n303), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n332), .A2(new_n333), .B1(new_n337), .B2(new_n291), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n243), .ZN(new_n339));
  OAI221_X1 g138(.A(new_n265), .B1(new_n319), .B2(new_n321), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(G8gat), .B(G36gat), .Z(new_n341));
  XNOR2_X1  g140(.A(G64gat), .B(G92gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n331), .A2(KEYINPUT30), .A3(new_n340), .A4(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n340), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(new_n338), .B2(new_n321), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n347), .A2(new_n328), .B1(new_n321), .B2(new_n320), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n345), .B1(new_n348), .B2(new_n214), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n344), .B1(new_n349), .B2(new_n343), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n331), .A2(new_n340), .A3(new_n343), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n351), .A3(new_n353), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n350), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G113gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(G120gat), .ZN(new_n359));
  INV_X1    g158(.A(G120gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(G113gat), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT68), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(G113gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(G120gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT68), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(G127gat), .A2(G134gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(G127gat), .A2(G134gat), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT1), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n362), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n372));
  OAI21_X1  g171(.A(G127gat), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G113gat), .B(G120gat), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n373), .B(new_n367), .C1(KEYINPUT1), .C2(new_n374), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n370), .A2(new_n375), .A3(KEYINPUT81), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT81), .B1(new_n370), .B2(new_n375), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n224), .A2(new_n226), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n228), .B1(new_n379), .B2(G162gat), .ZN(new_n380));
  OAI22_X1  g179(.A1(new_n238), .A2(new_n241), .B1(new_n380), .B2(new_n252), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n365), .B1(new_n363), .B2(new_n364), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT1), .ZN(new_n385));
  AND2_X1   g184(.A1(G127gat), .A2(G134gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(G127gat), .A2(G134gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT67), .B(G134gat), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n387), .B1(new_n390), .B2(G127gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n385), .B1(new_n359), .B2(new_n361), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n389), .A2(new_n366), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n256), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n382), .A2(new_n383), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n396), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(KEYINPUT39), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n370), .A2(new_n375), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n381), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n249), .A2(new_n250), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n393), .A2(new_n403), .A3(KEYINPUT4), .A4(new_n229), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n235), .A2(new_n237), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n241), .B1(new_n408), .B2(new_n246), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n380), .A2(new_n252), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT3), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n401), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n370), .A2(new_n375), .A3(KEYINPUT81), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n411), .A2(new_n242), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT82), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n378), .A2(new_n417), .A3(new_n242), .A4(new_n411), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n383), .B1(new_n407), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n399), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G1gat), .B(G29gat), .Z(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT39), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n420), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n422), .A2(KEYINPUT40), .A3(new_n428), .A4(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT5), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n382), .A2(new_n394), .ZN(new_n433));
  INV_X1    g232(.A(new_n383), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n402), .A2(new_n404), .A3(new_n383), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n419), .B2(new_n438), .ZN(new_n439));
  AOI211_X1 g238(.A(KEYINPUT83), .B(new_n437), .C1(new_n416), .C2(new_n418), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n434), .A2(KEYINPUT5), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n407), .A2(new_n419), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n428), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n428), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(new_n421), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n283), .B1(new_n357), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT38), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT37), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n349), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n343), .B1(new_n349), .B2(new_n452), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI22_X1  g254(.A1(new_n338), .A2(new_n339), .B1(new_n321), .B2(new_n319), .ZN(new_n456));
  INV_X1    g255(.A(new_n265), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n348), .B2(new_n214), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT38), .B1(new_n459), .B2(KEYINPUT37), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n352), .ZN(new_n462));
  XOR2_X1   g261(.A(KEYINPUT87), .B(KEYINPUT6), .Z(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n462), .B1(new_n444), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n441), .A2(KEYINPUT86), .A3(new_n428), .A4(new_n443), .ZN(new_n466));
  INV_X1    g265(.A(new_n443), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n419), .A2(new_n438), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT83), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n419), .A2(new_n436), .A3(new_n438), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n467), .B1(new_n471), .B2(new_n435), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n466), .B(new_n463), .C1(new_n472), .C2(new_n428), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT86), .B1(new_n472), .B2(new_n428), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n461), .B(new_n465), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n455), .B1(new_n475), .B2(KEYINPUT90), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n441), .A2(new_n443), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(new_n427), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(new_n445), .A3(new_n466), .A4(new_n463), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT90), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n461), .A4(new_n465), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n450), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n326), .A2(new_n393), .ZN(new_n484));
  INV_X1    g283(.A(G227gat), .ZN(new_n485));
  INV_X1    g284(.A(G233gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n304), .B(new_n401), .C1(new_n324), .C2(new_n325), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT69), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT69), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n484), .A2(new_n491), .A3(new_n487), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n494), .A2(KEYINPUT32), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G15gat), .B(G43gat), .Z(new_n497));
  XNOR2_X1  g296(.A(G71gat), .B(G99gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n484), .A2(new_n488), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n485), .B2(new_n486), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n505), .A2(KEYINPUT34), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(KEYINPUT34), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT32), .B1(new_n501), .B2(new_n494), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n490), .B2(new_n492), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT72), .ZN(new_n512));
  AOI211_X1 g311(.A(new_n512), .B(new_n509), .C1(new_n490), .C2(new_n492), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n503), .B(new_n508), .C1(new_n511), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT74), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n510), .B(KEYINPUT72), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT74), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n508), .A4(new_n503), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n503), .B1(new_n511), .B2(new_n513), .ZN(new_n519));
  INV_X1    g318(.A(new_n508), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n515), .A2(new_n518), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n519), .B1(KEYINPUT73), .B2(new_n508), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n508), .A2(KEYINPUT73), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(new_n516), .A3(new_n503), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n526), .A3(KEYINPUT36), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n343), .B1(new_n331), .B2(new_n340), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n462), .B2(KEYINPUT30), .ZN(new_n529));
  INV_X1    g328(.A(new_n356), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(new_n354), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n444), .A2(new_n464), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n480), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n523), .B(new_n527), .C1(new_n533), .C2(new_n283), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT35), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n274), .A2(new_n277), .ZN(new_n536));
  INV_X1    g335(.A(new_n280), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n274), .A2(new_n277), .A3(new_n280), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n540), .B1(new_n524), .B2(new_n526), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n535), .B1(new_n541), .B2(new_n533), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT35), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n532), .B1(new_n473), .B2(new_n474), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n544), .A3(new_n357), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n515), .A2(new_n518), .A3(new_n521), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI22_X1  g346(.A1(new_n483), .A2(new_n534), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT100), .ZN(new_n549));
  NAND2_X1  g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552));
  INV_X1    g351(.A(G85gat), .ZN(new_n553));
  INV_X1    g352(.A(G92gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(KEYINPUT8), .A2(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT98), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G99gat), .B(G106gat), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n556), .B(KEYINPUT98), .ZN(new_n561));
  INV_X1    g360(.A(new_n559), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR3_X1   g363(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n565), .A2(KEYINPUT92), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(KEYINPUT92), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G29gat), .A2(G36gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT91), .ZN(new_n572));
  XNOR2_X1  g371(.A(G43gat), .B(G50gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT15), .ZN(new_n574));
  XOR2_X1   g373(.A(G43gat), .B(G50gat), .Z(new_n575));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n570), .A2(new_n572), .A3(new_n574), .A4(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n569), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n572), .B1(new_n579), .B2(new_n565), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(KEYINPUT15), .A3(new_n573), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n564), .A2(new_n582), .B1(KEYINPUT41), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n578), .A2(KEYINPUT17), .A3(new_n581), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n586), .A2(new_n560), .A3(new_n563), .A4(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G190gat), .B(G218gat), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT97), .ZN(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n590), .B1(new_n584), .B2(new_n588), .ZN(new_n598));
  OR3_X1    g397(.A1(new_n592), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n592), .B2(new_n598), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G71gat), .B(G78gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT94), .Z(new_n603));
  INV_X1    g402(.A(KEYINPUT9), .ZN(new_n604));
  INV_X1    g403(.A(G71gat), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n604), .B1(new_n605), .B2(new_n271), .ZN(new_n606));
  INV_X1    g405(.A(G64gat), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n607), .A2(G57gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(G57gat), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT95), .B(G57gat), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n608), .B1(new_n612), .B2(G64gat), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n602), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n602), .A2(new_n614), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n606), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n611), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(G127gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G15gat), .B(G22gat), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT16), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n625), .B1(new_n626), .B2(G1gat), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(G1gat), .B2(new_n625), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G8gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n618), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(KEYINPUT21), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n624), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n223), .ZN(new_n634));
  XNOR2_X1  g433(.A(G183gat), .B(G211gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n624), .A2(new_n631), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n631), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n640), .A3(new_n636), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n601), .B1(new_n638), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n564), .A2(new_n630), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n618), .A2(new_n560), .A3(new_n563), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n646), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n643), .A2(new_n650), .A3(new_n644), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n564), .A2(KEYINPUT10), .A3(new_n630), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  NAND3_X1  g456(.A1(new_n648), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n647), .B2(new_n653), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(new_n660), .A3(KEYINPUT99), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT99), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n662), .B(new_n659), .C1(new_n647), .C2(new_n653), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(G8gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n628), .B(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n586), .A2(new_n666), .A3(new_n587), .ZN(new_n667));
  NAND2_X1  g466(.A1(G229gat), .A2(G233gat), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n582), .A2(new_n629), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT18), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n668), .B(KEYINPUT13), .Z(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n666), .A2(new_n581), .A3(new_n578), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n669), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n677), .A2(KEYINPUT93), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(KEYINPUT93), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n672), .B(new_n673), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G113gat), .B(G141gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G197gat), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT11), .B(G169gat), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT12), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n678), .A2(new_n679), .ZN(new_n687));
  INV_X1    g486(.A(new_n685), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n687), .A2(new_n688), .A3(new_n672), .A4(new_n673), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n642), .A2(new_n664), .A3(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n548), .A2(new_n549), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n549), .B1(new_n548), .B2(new_n691), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n544), .B(KEYINPUT101), .Z(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT102), .B(G1gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1324gat));
  INV_X1    g498(.A(new_n694), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n665), .B1(new_n700), .B2(new_n531), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n626), .A2(new_n665), .ZN(new_n702));
  NOR2_X1   g501(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n703));
  NOR4_X1   g502(.A1(new_n694), .A2(new_n357), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT42), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n705), .B1(KEYINPUT42), .B2(new_n704), .ZN(G1325gat));
  OR3_X1    g505(.A1(new_n694), .A2(G15gat), .A3(new_n546), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n523), .A2(new_n527), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n708), .A2(KEYINPUT103), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(KEYINPUT103), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G15gat), .B1(new_n694), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n707), .A2(new_n712), .ZN(G1326gat));
  NOR2_X1   g512(.A1(new_n694), .A2(new_n283), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  AND2_X1   g515(.A1(new_n548), .A2(new_n601), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n638), .A2(new_n641), .ZN(new_n718));
  INV_X1    g517(.A(new_n664), .ZN(new_n719));
  INV_X1    g518(.A(new_n690), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n722), .A2(G29gat), .A3(new_n696), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT45), .Z(new_n724));
  XOR2_X1   g523(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n725));
  AND3_X1   g524(.A1(new_n548), .A2(new_n601), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n548), .B2(new_n601), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(new_n695), .A3(new_n721), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G29gat), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n724), .A2(new_n731), .ZN(G1328gat));
  NOR3_X1   g531(.A1(new_n722), .A2(G36gat), .A3(new_n357), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n729), .A2(new_n531), .A3(new_n721), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G36gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(G1329gat));
  INV_X1    g536(.A(new_n708), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n729), .A2(new_n738), .A3(new_n721), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G43gat), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n722), .A2(G43gat), .A3(new_n546), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(KEYINPUT47), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n711), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n744), .B(new_n721), .C1(new_n726), .C2(new_n728), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n745), .A2(KEYINPUT105), .A3(G43gat), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT105), .B1(new_n745), .B2(G43gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n746), .A2(new_n747), .A3(new_n741), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n743), .B1(new_n748), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g548(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n750));
  INV_X1    g549(.A(new_n722), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n283), .A2(G50gat), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n540), .B(new_n721), .C1(new_n726), .C2(new_n728), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G50gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1331gat));
  AND2_X1   g557(.A1(new_n642), .A2(new_n720), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n548), .A2(new_n719), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n695), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(new_n612), .Z(G1332gat));
  AOI21_X1  g561(.A(new_n357), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT107), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT108), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n764), .B(new_n767), .ZN(G1333gat));
  AOI21_X1  g567(.A(new_n605), .B1(new_n760), .B2(new_n744), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n546), .A2(G71gat), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n760), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g571(.A1(new_n760), .A2(new_n540), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT109), .B(G78gat), .Z(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1335gat));
  NOR2_X1   g574(.A1(new_n718), .A2(new_n690), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n548), .A2(new_n601), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n548), .A2(KEYINPUT51), .A3(new_n601), .A4(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n781), .A2(KEYINPUT110), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(KEYINPUT110), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n696), .A2(G85gat), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n782), .A2(new_n719), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n718), .A2(new_n664), .A3(new_n690), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n729), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n695), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n788), .B2(new_n553), .ZN(G1336gat));
  OAI211_X1 g588(.A(new_n531), .B(new_n786), .C1(new_n726), .C2(new_n728), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n554), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n791), .B2(new_n790), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n719), .A2(new_n554), .A3(new_n531), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n779), .B2(new_n780), .ZN(new_n795));
  XNOR2_X1  g594(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n790), .A2(G92gat), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n799), .B2(new_n795), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1337gat));
  NAND2_X1  g600(.A1(new_n787), .A2(new_n744), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G99gat), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n546), .A2(G99gat), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n782), .A2(new_n719), .A3(new_n783), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(G1338gat));
  NOR3_X1   g605(.A1(new_n283), .A2(G106gat), .A3(new_n664), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n779), .B2(new_n780), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n540), .B(new_n786), .C1(new_n726), .C2(new_n728), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(G106gat), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n810), .B2(G106gat), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n811), .A2(new_n813), .A3(KEYINPUT53), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  AOI221_X4 g614(.A(new_n809), .B1(new_n812), .B2(new_n815), .C1(G106gat), .C2(new_n810), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n814), .A2(new_n816), .ZN(G1339gat));
  NAND2_X1  g616(.A1(new_n759), .A2(new_n664), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n667), .A2(new_n669), .ZN(new_n819));
  INV_X1    g618(.A(new_n668), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT115), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n819), .A2(new_n823), .A3(new_n820), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n669), .A2(new_n676), .A3(new_n675), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT116), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n822), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n684), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(new_n689), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830));
  AOI211_X1 g629(.A(KEYINPUT54), .B(new_n649), .C1(new_n651), .C2(new_n652), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n657), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n653), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(KEYINPUT114), .A3(new_n659), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n651), .A2(new_n652), .A3(new_n649), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n653), .A2(new_n833), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n832), .A2(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n829), .B(new_n601), .C1(new_n838), .C2(KEYINPUT55), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n836), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n831), .A2(new_n830), .A3(new_n657), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT114), .B1(new_n834), .B2(new_n659), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n658), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n661), .A2(new_n828), .A3(new_n663), .A4(new_n689), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT117), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n829), .A2(new_n849), .A3(new_n663), .A4(new_n661), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n690), .B1(new_n838), .B2(KEYINPUT55), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n848), .B(new_n850), .C1(new_n845), .C2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n601), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n846), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n818), .B1(new_n854), .B2(new_n718), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT118), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n818), .B(new_n857), .C1(new_n854), .C2(new_n718), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n856), .A2(new_n283), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n546), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n696), .A2(new_n531), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n720), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n856), .A2(new_n858), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n541), .A2(new_n357), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n695), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n690), .A2(new_n358), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT119), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n863), .B1(new_n866), .B2(new_n868), .ZN(G1340gat));
  INV_X1    g668(.A(new_n866), .ZN(new_n870));
  AOI21_X1  g669(.A(G120gat), .B1(new_n870), .B2(new_n719), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n862), .A2(new_n360), .A3(new_n664), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(G1341gat));
  NAND3_X1  g672(.A1(new_n870), .A2(new_n623), .A3(new_n718), .ZN(new_n874));
  INV_X1    g673(.A(new_n718), .ZN(new_n875));
  OAI21_X1  g674(.A(G127gat), .B1(new_n862), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1342gat));
  OR2_X1    g676(.A1(new_n853), .A2(new_n390), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT56), .B1(new_n866), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(KEYINPUT120), .B(KEYINPUT56), .C1(new_n866), .C2(new_n878), .ZN(new_n882));
  OR3_X1    g681(.A1(new_n866), .A2(KEYINPUT56), .A3(new_n878), .ZN(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n862), .B2(new_n853), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n884), .ZN(G1343gat));
  NAND2_X1  g684(.A1(new_n861), .A2(new_n708), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n847), .B1(new_n845), .B2(new_n851), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n846), .B1(new_n853), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n818), .B1(new_n888), .B2(new_n718), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n540), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n886), .B1(new_n890), .B2(KEYINPUT57), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n856), .A2(new_n892), .A3(new_n540), .A4(new_n858), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n891), .A2(new_n893), .A3(new_n690), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT58), .B1(new_n894), .B2(G141gat), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n711), .A2(new_n540), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n864), .A2(new_n896), .A3(new_n898), .A4(new_n695), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n856), .A2(new_n695), .A3(new_n858), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT121), .B1(new_n900), .B2(new_n897), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n357), .A3(new_n901), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n720), .A2(G141gat), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n895), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n720), .A2(G141gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n357), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n900), .A2(new_n897), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n908), .B1(G141gat), .B2(new_n894), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n904), .B1(new_n905), .B2(new_n909), .ZN(G1344gat));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n891), .A2(new_n893), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n911), .B(G148gat), .C1(new_n912), .C2(new_n664), .ZN(new_n913));
  INV_X1    g712(.A(G148gat), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n856), .A2(KEYINPUT57), .A3(new_n540), .A4(new_n858), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n890), .A2(new_n892), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n886), .A2(new_n664), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n913), .B1(new_n919), .B2(new_n911), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n719), .A2(new_n914), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n902), .B2(new_n921), .ZN(G1345gat));
  NAND2_X1  g721(.A1(new_n718), .A2(new_n379), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT122), .Z(new_n924));
  NOR2_X1   g723(.A1(new_n912), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n899), .A2(new_n901), .A3(new_n357), .A4(new_n718), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n254), .ZN(G1346gat));
  NOR3_X1   g726(.A1(new_n912), .A2(new_n222), .A3(new_n853), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n899), .A2(new_n901), .A3(new_n357), .A4(new_n601), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(new_n222), .ZN(G1347gat));
  NOR2_X1   g729(.A1(new_n695), .A2(new_n357), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n859), .A2(new_n860), .A3(new_n690), .A4(new_n931), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT123), .B1(new_n932), .B2(G169gat), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n524), .A2(new_n526), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n859), .A2(new_n935), .A3(new_n931), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n690), .A2(new_n287), .ZN(new_n937));
  OAI22_X1  g736(.A1(new_n933), .A2(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1348gat));
  NAND4_X1  g737(.A1(new_n856), .A2(new_n283), .A3(new_n858), .A4(new_n931), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(new_n546), .A3(new_n664), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n719), .A2(new_n288), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n940), .A2(new_n288), .B1(new_n936), .B2(new_n941), .ZN(G1349gat));
  AND2_X1   g741(.A1(new_n718), .A2(new_n292), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n859), .A2(new_n935), .A3(new_n931), .A4(new_n943), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n939), .A2(new_n546), .A3(new_n875), .ZN(new_n945));
  INV_X1    g744(.A(G183gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g747(.A1(new_n859), .A2(new_n860), .A3(new_n601), .A4(new_n931), .ZN(new_n949));
  NOR2_X1   g748(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n293), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n601), .A2(new_n293), .ZN(new_n954));
  OAI22_X1  g753(.A1(new_n952), .A2(new_n953), .B1(new_n936), .B2(new_n954), .ZN(G1351gat));
  NAND2_X1  g754(.A1(new_n711), .A2(new_n931), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n917), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n720), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n856), .A2(new_n540), .A3(new_n858), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n960), .A2(new_n956), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n720), .A2(G197gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT125), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n961), .A2(KEYINPUT125), .A3(new_n962), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  OAI21_X1  g764(.A(G204gat), .B1(new_n958), .B2(new_n664), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n664), .A2(G204gat), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n960), .A2(new_n956), .A3(new_n968), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT126), .A3(new_n967), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT126), .B1(new_n969), .B2(new_n967), .ZN(new_n971));
  OAI221_X1 g770(.A(new_n966), .B1(new_n967), .B2(new_n969), .C1(new_n970), .C2(new_n971), .ZN(G1353gat));
  INV_X1    g771(.A(G211gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n961), .A2(new_n973), .A3(new_n718), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n917), .A2(new_n718), .A3(new_n957), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  NAND2_X1  g777(.A1(new_n601), .A2(G218gat), .ZN(new_n979));
  XOR2_X1   g778(.A(new_n979), .B(KEYINPUT127), .Z(new_n980));
  NOR2_X1   g779(.A1(new_n958), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(G218gat), .B1(new_n961), .B2(new_n601), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


