//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT70), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT71), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G120gat), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G113gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n205), .B(new_n206), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n204), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G127gat), .B(G134gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n204), .A2(new_n211), .A3(new_n213), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G148gat), .ZN(new_n219));
  INV_X1    g018(.A(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n219), .A2(new_n221), .B1(KEYINPUT2), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n224));
  INV_X1    g023(.A(new_n222), .ZN(new_n225));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G155gat), .ZN(new_n228));
  INV_X1    g027(.A(G162gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(KEYINPUT80), .A3(new_n222), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n223), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n222), .ZN(new_n233));
  XNOR2_X1  g032(.A(G141gat), .B(G148gat), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n224), .B(new_n233), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n202), .B1(new_n217), .B2(new_n237), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n204), .A2(new_n211), .A3(new_n213), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n213), .B1(new_n204), .B2(new_n211), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n202), .B(new_n237), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT5), .ZN(new_n244));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(new_n239), .B2(new_n240), .ZN(new_n247));
  INV_X1    g046(.A(new_n237), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT81), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT3), .B1(new_n232), .B2(new_n236), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n247), .A2(new_n249), .A3(new_n250), .A4(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n243), .A2(new_n244), .A3(new_n245), .A4(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n247), .A2(new_n250), .A3(new_n248), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n217), .A2(new_n237), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT82), .ZN(new_n258));
  INV_X1    g057(.A(new_n245), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n253), .B(new_n245), .C1(new_n238), .C2(new_n242), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT5), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n254), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(G1gat), .B(G29gat), .Z(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT0), .ZN(new_n266));
  XNOR2_X1  g065(.A(G57gat), .B(G85gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(KEYINPUT6), .A3(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n268), .B(new_n254), .C1(new_n262), .C2(new_n263), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n268), .B(KEYINPUT90), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n259), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT82), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n277), .A2(KEYINPUT5), .A3(new_n260), .A4(new_n261), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n275), .B1(new_n278), .B2(new_n254), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n270), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT35), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G211gat), .A2(G218gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT22), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(G197gat), .A2(G204gat), .ZN(new_n286));
  AND2_X1   g085(.A1(G197gat), .A2(G204gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G211gat), .B(G218gat), .Z(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G211gat), .B(G218gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(G197gat), .B(G204gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n292), .A3(new_n285), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n290), .A2(KEYINPUT75), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT75), .B1(new_n290), .B2(new_n293), .ZN(new_n295));
  OAI22_X1  g094(.A1(new_n251), .A2(KEYINPUT29), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT29), .B1(new_n290), .B2(new_n293), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n248), .B1(KEYINPUT3), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G228gat), .ZN(new_n300));
  INV_X1    g099(.A(G233gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT84), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT84), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n299), .A2(new_n306), .A3(new_n303), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n288), .A2(new_n289), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n291), .B1(new_n285), .B2(new_n292), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT3), .B1(new_n311), .B2(KEYINPUT85), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT85), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n237), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n294), .A2(new_n295), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n237), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n302), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT86), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n311), .A2(KEYINPUT85), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n317), .B1(new_n297), .B2(new_n313), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n248), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n302), .A4(new_n296), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n305), .A2(new_n307), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT87), .ZN(new_n327));
  OAI21_X1  g126(.A(G22gat), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n305), .A2(new_n307), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(new_n325), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n329), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT88), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n330), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT87), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n326), .A2(new_n327), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT88), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .A4(G22gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G22gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n326), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G78gat), .B(G106gat), .ZN(new_n341));
  INV_X1    g140(.A(G50gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n338), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n333), .A2(G22gat), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n346), .B1(new_n350), .B2(new_n340), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n282), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT65), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT66), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n358), .A2(KEYINPUT66), .A3(new_n361), .ZN(new_n365));
  AND2_X1   g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(KEYINPUT23), .B2(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n369));
  INV_X1    g168(.A(G169gat), .ZN(new_n370));
  INV_X1    g169(.A(G176gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n369), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(KEYINPUT68), .A2(KEYINPUT25), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n368), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT68), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n368), .B2(new_n374), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n364), .B(new_n365), .C1(new_n376), .C2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G183gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT27), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT27), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G183gat), .ZN(new_n383));
  INV_X1    g182(.A(G190gat), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n372), .B1(new_n366), .B2(KEYINPUT26), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT26), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n367), .A2(new_n388), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n385), .A2(new_n386), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n381), .A2(new_n383), .A3(new_n384), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT28), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(KEYINPUT69), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n391), .A2(new_n393), .B1(G183gat), .B2(G190gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n361), .A2(new_n354), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n374), .A3(new_n368), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n390), .A2(new_n394), .B1(new_n396), .B2(KEYINPUT25), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n217), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n379), .A2(new_n397), .A3(new_n216), .A4(new_n215), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT34), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT34), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n402), .B(KEYINPUT64), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n401), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT32), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT72), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n401), .B2(new_n407), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n399), .A2(KEYINPUT72), .A3(new_n406), .A4(new_n400), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT73), .B(KEYINPUT33), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n412), .B2(new_n413), .ZN(new_n416));
  XOR2_X1   g215(.A(G15gat), .B(G43gat), .Z(new_n417));
  XNOR2_X1  g216(.A(G71gat), .B(G99gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n414), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  AOI221_X4 g220(.A(new_n410), .B1(new_n415), .B2(new_n419), .C1(new_n412), .C2(new_n413), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n409), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n412), .A2(new_n413), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT32), .ZN(new_n425));
  INV_X1    g224(.A(new_n415), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n427), .A3(new_n419), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n414), .B1(new_n416), .B2(new_n420), .ZN(new_n429));
  INV_X1    g228(.A(new_n409), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT74), .B1(new_n423), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n433), .A2(KEYINPUT74), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G8gat), .B(G36gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G64gat), .B(G92gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(G226gat), .A2(G233gat), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n441), .B1(new_n398), .B2(new_n308), .ZN(new_n442));
  INV_X1    g241(.A(new_n316), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n379), .A2(new_n397), .A3(KEYINPUT76), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT76), .B1(new_n379), .B2(new_n397), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n445), .B1(new_n448), .B2(new_n441), .ZN(new_n449));
  NOR4_X1   g248(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT78), .A4(new_n440), .ZN(new_n450));
  OAI211_X1 g249(.A(KEYINPUT79), .B(new_n444), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n441), .B1(new_n448), .B2(new_n308), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n398), .A2(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT77), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT77), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n398), .A2(new_n455), .A3(new_n441), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n443), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n448), .A2(new_n445), .A3(new_n441), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT76), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n398), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n379), .A2(new_n397), .A3(KEYINPUT76), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n441), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT78), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT79), .B1(new_n466), .B2(new_n444), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n439), .B1(new_n459), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n444), .B1(new_n449), .B2(new_n450), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT79), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n471), .A2(new_n458), .A3(new_n451), .A4(new_n438), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(KEYINPUT30), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n459), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n471), .A4(new_n438), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n473), .A2(KEYINPUT89), .A3(new_n476), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n353), .A2(new_n435), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n268), .B1(new_n278), .B2(new_n254), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n270), .B1(new_n273), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n347), .B1(new_n332), .B2(new_n337), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n431), .B(new_n423), .C1(new_n485), .C2(new_n351), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT35), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n243), .A2(new_n253), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n259), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(KEYINPUT39), .C1(new_n259), .C2(new_n257), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT91), .B(KEYINPUT39), .Z(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n259), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT92), .A3(new_n275), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT92), .B1(new_n493), .B2(new_n275), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT93), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT40), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n499), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(new_n491), .C1(new_n495), .C2(new_n496), .ZN(new_n502));
  INV_X1    g301(.A(new_n279), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n504), .B1(new_n479), .B2(new_n480), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n349), .A2(new_n352), .ZN(new_n506));
  INV_X1    g305(.A(new_n472), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n280), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT29), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n454), .B(new_n456), .C1(new_n510), .C2(new_n441), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n511), .B2(new_n316), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n442), .A2(new_n316), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n466), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT38), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n471), .A2(new_n458), .A3(new_n451), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n515), .B(new_n439), .C1(new_n516), .C2(KEYINPUT37), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT38), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n439), .A2(KEYINPUT37), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n468), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(KEYINPUT37), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n506), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n505), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n432), .B2(new_n434), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n423), .A2(KEYINPUT36), .A3(new_n431), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n485), .A2(new_n351), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n484), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n488), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n534), .A2(KEYINPUT96), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n535), .A2(G1gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(G1gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT16), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(G8gat), .Z(new_n541));
  INV_X1    g340(.A(G43gat), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT15), .B1(new_n542), .B2(G50gat), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(new_n542), .B2(G50gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT95), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n342), .B2(G43gat), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT94), .B1(new_n542), .B2(G50gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(new_n342), .A3(G43gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(KEYINPUT95), .A3(G50gat), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n546), .A2(new_n547), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT15), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G29gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n555));
  AND2_X1   g354(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n555), .B1(new_n558), .B2(G36gat), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n544), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n559), .A2(new_n544), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT17), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n541), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n540), .B(G8gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n562), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n567), .A2(KEYINPUT18), .A3(new_n568), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n565), .B(new_n562), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n568), .B(KEYINPUT13), .Z(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n571), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(G197gat), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT11), .B(G169gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n580), .B(KEYINPUT12), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n571), .A2(new_n583), .A3(new_n572), .A4(new_n575), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n533), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G57gat), .B(G64gat), .Z(new_n587));
  INV_X1    g386(.A(KEYINPUT9), .ZN(new_n588));
  INV_X1    g387(.A(G71gat), .ZN(new_n589));
  INV_X1    g388(.A(G78gat), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G71gat), .B(G78gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n587), .A2(new_n593), .A3(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G183gat), .B(G211gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n595), .A2(new_n596), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n565), .B1(KEYINPUT21), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(KEYINPUT41), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G134gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(new_n229), .ZN(new_n619));
  NAND2_X1  g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT7), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(G85gat), .ZN(new_n623));
  INV_X1    g422(.A(G92gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G99gat), .B(G106gat), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n629));
  INV_X1    g428(.A(new_n627), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(new_n621), .A3(new_n625), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n626), .A2(KEYINPUT99), .A3(new_n627), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT100), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n563), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n634), .A2(new_n562), .B1(KEYINPUT41), .B2(new_n616), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G190gat), .B(G218gat), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n619), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n638), .A2(new_n639), .ZN(new_n643));
  OR3_X1    g442(.A1(new_n642), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n640), .B2(new_n643), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n615), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n608), .B1(new_n633), .B2(new_n632), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n597), .B1(new_n628), .B2(new_n631), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n634), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT102), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n657), .A3(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(G230gat), .A2(G233gat), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n651), .A2(new_n652), .A3(new_n659), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT103), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n660), .A2(new_n669), .A3(new_n666), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n659), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n653), .B2(new_n654), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n665), .B1(new_n673), .B2(new_n661), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n649), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n660), .A2(new_n669), .A3(new_n666), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n669), .B1(new_n660), .B2(new_n666), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n649), .B(new_n674), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n648), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n586), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n483), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT105), .B(G1gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1324gat));
  AND3_X1   g486(.A1(new_n473), .A2(KEYINPUT89), .A3(new_n476), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT89), .B1(new_n473), .B2(new_n476), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n586), .A2(new_n691), .A3(new_n683), .ZN(new_n692));
  AND2_X1   g491(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n692), .A2(G8gat), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT42), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(KEYINPUT42), .B2(new_n695), .ZN(G1325gat));
  OAI21_X1  g497(.A(G15gat), .B1(new_n684), .B2(new_n529), .ZN(new_n699));
  INV_X1    g498(.A(new_n435), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n700), .A2(G15gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n684), .B2(new_n701), .ZN(G1326gat));
  NOR2_X1   g501(.A1(new_n684), .A2(new_n506), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT43), .B(G22gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  NOR3_X1   g504(.A1(new_n614), .A2(new_n646), .A3(new_n680), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n586), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n707), .A2(G29gat), .A3(new_n483), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT45), .Z(new_n709));
  AND3_X1   g508(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(new_n688), .B2(new_n689), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n316), .B1(new_n452), .B2(new_n457), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n514), .A2(KEYINPUT37), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n519), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n468), .B2(new_n520), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n472), .B(new_n270), .C1(new_n273), .C2(new_n279), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n439), .B1(new_n516), .B2(KEYINPUT37), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n509), .B1(new_n474), .B2(new_n471), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT38), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n530), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n711), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n527), .A2(new_n528), .B1(new_n484), .B2(new_n530), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n723), .B1(new_n722), .B2(new_n724), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n488), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n646), .A2(KEYINPUT44), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n533), .A2(new_n647), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n727), .A2(new_n728), .B1(new_n729), .B2(KEYINPUT44), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n615), .A2(new_n585), .A3(new_n681), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n730), .A2(new_n483), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n709), .B1(new_n554), .B2(new_n732), .ZN(G1328gat));
  NOR3_X1   g532(.A1(new_n730), .A2(new_n690), .A3(new_n731), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(KEYINPUT107), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(KEYINPUT107), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(G36gat), .A3(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n707), .A2(G36gat), .A3(new_n690), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT46), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1329gat));
  NOR2_X1   g539(.A1(new_n730), .A2(new_n731), .ZN(new_n741));
  INV_X1    g540(.A(new_n529), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n542), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n744), .B2(new_n743), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n707), .A2(G43gat), .A3(new_n700), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n542), .B1(new_n741), .B2(new_n742), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n748), .B1(new_n751), .B2(new_n747), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1330gat));
  NOR3_X1   g552(.A1(new_n707), .A2(G50gat), .A3(new_n506), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n741), .A2(new_n530), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(G50gat), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g556(.A(new_n488), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT106), .B1(new_n525), .B2(new_n532), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n722), .A2(new_n724), .A3(new_n723), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n585), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n648), .A2(new_n762), .A3(new_n680), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n483), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g568(.A(new_n764), .B(KEYINPUT109), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n766), .A2(KEYINPUT110), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n773), .A3(new_n691), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT49), .B(G64gat), .Z(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(G1333gat));
  NOR2_X1   g576(.A1(new_n529), .A2(new_n589), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n772), .A2(new_n773), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n589), .B1(new_n770), .B2(new_n700), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n779), .A2(KEYINPUT50), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT50), .B1(new_n779), .B2(new_n780), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(G1334gat));
  NAND3_X1  g582(.A1(new_n772), .A2(new_n773), .A3(new_n530), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n615), .A2(new_n762), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n681), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n786), .B1(new_n730), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n728), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n759), .A2(new_n760), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n488), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n533), .B2(new_n647), .ZN(new_n795));
  OAI211_X1 g594(.A(KEYINPUT111), .B(new_n788), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(G85gat), .B1(new_n797), .B2(new_n483), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n787), .A2(new_n646), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n761), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n727), .A2(KEYINPUT51), .A3(new_n800), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n680), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n767), .A2(new_n623), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n798), .B1(new_n806), .B2(new_n807), .ZN(G1336gat));
  NOR2_X1   g607(.A1(new_n690), .A2(G92gat), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n681), .B(new_n810), .C1(new_n802), .C2(new_n804), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n788), .B1(new_n793), .B2(new_n795), .ZN(new_n813));
  OAI21_X1  g612(.A(G92gat), .B1(new_n813), .B2(new_n690), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n790), .A2(new_n691), .A3(new_n796), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G92gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n812), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n817), .B1(new_n820), .B2(KEYINPUT52), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n811), .B1(new_n818), .B2(G92gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n822), .A2(KEYINPUT112), .A3(new_n815), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n816), .B1(new_n821), .B2(new_n823), .ZN(G1337gat));
  OAI21_X1  g623(.A(G99gat), .B1(new_n797), .B2(new_n529), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n700), .A2(G99gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n806), .B2(new_n826), .ZN(G1338gat));
  OAI21_X1  g626(.A(G106gat), .B1(new_n813), .B2(new_n506), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n506), .A2(G106gat), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n828), .B(new_n829), .C1(new_n806), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n806), .A2(new_n830), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n790), .A2(new_n530), .A3(new_n796), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(G106gat), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n831), .B1(new_n834), .B2(new_n829), .ZN(G1339gat));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT54), .B1(new_n655), .B2(new_n659), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n672), .B1(new_n655), .B2(KEYINPUT102), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n658), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n664), .B1(new_n673), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n836), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n660), .ZN(new_n844));
  OAI211_X1 g643(.A(KEYINPUT55), .B(new_n841), .C1(new_n844), .C2(new_n837), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n671), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n671), .A2(new_n843), .A3(new_n848), .A4(new_n845), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n567), .A2(new_n568), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n573), .A2(new_n574), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n580), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n584), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n644), .A2(new_n645), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n847), .A2(new_n585), .A3(new_n849), .ZN(new_n858));
  INV_X1    g657(.A(new_n679), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n854), .B1(new_n675), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n647), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT114), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n860), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n863), .A2(new_n646), .B1(new_n850), .B2(new_n855), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n862), .A2(new_n866), .A3(new_n615), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n648), .A2(new_n762), .A3(new_n681), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n483), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n691), .A2(new_n486), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(G113gat), .B1(new_n872), .B2(new_n585), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n615), .B1(new_n864), .B2(new_n865), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n857), .A2(new_n861), .A3(KEYINPUT114), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n868), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n876), .A2(KEYINPUT115), .A3(new_n506), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT115), .B1(new_n876), .B2(new_n506), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n690), .A2(new_n767), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n700), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n762), .A2(new_n207), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n873), .B1(new_n884), .B2(new_n885), .ZN(G1340gat));
  NAND3_X1  g685(.A1(new_n880), .A2(new_n680), .A3(new_n882), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(G120gat), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n887), .B2(G120gat), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n680), .A2(new_n209), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT117), .Z(new_n892));
  OAI22_X1  g691(.A1(new_n889), .A2(new_n890), .B1(new_n871), .B2(new_n892), .ZN(G1341gat));
  OAI21_X1  g692(.A(G127gat), .B1(new_n883), .B2(new_n615), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n615), .A2(G127gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n871), .B2(new_n895), .ZN(G1342gat));
  NOR2_X1   g695(.A1(new_n646), .A2(G134gat), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  OR3_X1    g697(.A1(new_n871), .A2(KEYINPUT118), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT118), .B1(new_n871), .B2(new_n898), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G134gat), .B1(new_n883), .B2(new_n646), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n901), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(KEYINPUT56), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT119), .B(new_n900), .C1(new_n899), .C2(new_n901), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n902), .B(new_n903), .C1(new_n906), .C2(new_n907), .ZN(G1343gat));
  NOR2_X1   g707(.A1(new_n742), .A2(new_n506), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n869), .A2(new_n690), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n218), .A3(new_n585), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n860), .B1(new_n762), .B2(new_n846), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n646), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n856), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n615), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n868), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(KEYINPUT57), .A3(new_n530), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n506), .B1(new_n867), .B2(new_n868), .ZN(new_n918));
  XNOR2_X1  g717(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n917), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n742), .A2(new_n881), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n921), .A2(new_n585), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n911), .B1(new_n923), .B2(new_n218), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n926));
  INV_X1    g725(.A(new_n846), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n855), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT121), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n614), .B1(new_n929), .B2(KEYINPUT121), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n930), .A2(new_n931), .B1(new_n683), .B2(new_n762), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n926), .B1(new_n932), .B2(new_n506), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n920), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n922), .A2(new_n680), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT59), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n921), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n910), .B2(new_n680), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n939), .B(new_n941), .C1(G148gat), .C2(new_n942), .ZN(G1345gat));
  NAND3_X1  g742(.A1(new_n910), .A2(new_n228), .A3(new_n614), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n921), .A2(new_n614), .A3(new_n922), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n228), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n946), .B(new_n947), .ZN(G1346gat));
  AOI21_X1  g747(.A(new_n920), .B1(new_n876), .B2(new_n530), .ZN(new_n949));
  INV_X1    g748(.A(new_n917), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n647), .B(new_n922), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n921), .A2(KEYINPUT123), .A3(new_n647), .A4(new_n922), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(G162gat), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n910), .A2(new_n229), .A3(new_n647), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(KEYINPUT124), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1347gat));
  NOR2_X1   g760(.A1(new_n690), .A2(new_n767), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AOI211_X1 g762(.A(new_n486), .B(new_n963), .C1(new_n867), .C2(new_n868), .ZN(new_n964));
  AOI21_X1  g763(.A(G169gat), .B1(new_n964), .B2(new_n585), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n435), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n879), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n762), .A2(new_n370), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(G1348gat));
  NAND3_X1  g768(.A1(new_n964), .A2(new_n371), .A3(new_n680), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n967), .A2(new_n680), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n970), .B1(new_n972), .B2(new_n371), .ZN(G1349gat));
  INV_X1    g772(.A(new_n966), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n614), .B(new_n974), .C1(new_n877), .C2(new_n878), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n614), .A2(new_n381), .A3(new_n383), .ZN(new_n976));
  AOI22_X1  g775(.A1(new_n975), .A2(G183gat), .B1(new_n964), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n977), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n978));
  NOR2_X1   g777(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n979));
  AND2_X1   g778(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n978), .A2(new_n981), .ZN(G1350gat));
  NAND3_X1  g781(.A1(new_n964), .A2(new_n384), .A3(new_n647), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n647), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n984), .B1(new_n985), .B2(G190gat), .ZN(new_n986));
  AOI211_X1 g785(.A(KEYINPUT61), .B(new_n384), .C1(new_n967), .C2(new_n647), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(G1351gat));
  AND3_X1   g787(.A1(new_n876), .A2(new_n909), .A3(new_n962), .ZN(new_n989));
  INV_X1    g788(.A(G197gat), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n989), .A2(new_n990), .A3(new_n585), .ZN(new_n991));
  XOR2_X1   g790(.A(new_n991), .B(KEYINPUT126), .Z(new_n992));
  AOI211_X1 g791(.A(new_n742), .B(new_n963), .C1(new_n933), .C2(new_n934), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n993), .A2(new_n585), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n992), .B1(new_n994), .B2(new_n990), .ZN(G1352gat));
  INV_X1    g794(.A(G204gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n989), .A2(new_n996), .A3(new_n680), .ZN(new_n997));
  XOR2_X1   g796(.A(new_n997), .B(KEYINPUT62), .Z(new_n998));
  AND2_X1   g797(.A1(new_n993), .A2(new_n680), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n998), .B1(new_n999), .B2(new_n996), .ZN(G1353gat));
  INV_X1    g799(.A(G211gat), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n989), .A2(new_n1001), .A3(new_n614), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n963), .A2(new_n742), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n935), .A2(new_n614), .A3(new_n1003), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(G1354gat));
  OAI21_X1  g806(.A(new_n647), .B1(new_n993), .B2(KEYINPUT127), .ZN(new_n1008));
  AND3_X1   g807(.A1(new_n935), .A2(KEYINPUT127), .A3(new_n1003), .ZN(new_n1009));
  OAI21_X1  g808(.A(G218gat), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g809(.A(G218gat), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n989), .A2(new_n1011), .A3(new_n647), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1010), .A2(new_n1012), .ZN(G1355gat));
endmodule


