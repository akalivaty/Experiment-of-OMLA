//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT65), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT67), .Z(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT68), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n473), .A3(KEYINPUT3), .ZN(new_n474));
  OR2_X1    g049(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  INV_X1    g052(.A(G101), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n471), .A2(new_n473), .ZN(new_n479));
  OAI22_X1  g054(.A1(new_n476), .A2(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n469), .B1(new_n480), .B2(new_n465), .ZN(G160));
  NOR2_X1   g056(.A1(new_n476), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n476), .A2(new_n465), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(new_n465), .B2(G112), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n483), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n466), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n474), .A2(KEYINPUT4), .A3(new_n475), .A4(new_n491), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n474), .A2(new_n475), .A3(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n498), .A2(KEYINPUT69), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT69), .B1(new_n498), .B2(new_n500), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n496), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  OR2_X1    g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n507), .A2(G62), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n512), .B1(new_n508), .B2(new_n509), .ZN(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT70), .B1(KEYINPUT71), .B2(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT70), .A2(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT6), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n519), .A2(new_n507), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT72), .B(G88), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n519), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n514), .A2(new_n522), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  XOR2_X1   g101(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n507), .ZN(new_n530));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  OR3_X1    g106(.A1(new_n530), .A2(KEYINPUT74), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT74), .B1(new_n530), .B2(new_n531), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n523), .A2(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n520), .A2(G89), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT76), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(new_n523), .A2(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n520), .A2(G90), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G651), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND2_X1  g123(.A1(new_n523), .A2(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n520), .A2(G81), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n545), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  AND2_X1   g135(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n519), .A2(G53), .A3(G543), .ZN(new_n562));
  NOR2_X1   g137(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n561), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n565), .B1(new_n564), .B2(new_n562), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n519), .A2(G91), .A3(new_n507), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n519), .A2(KEYINPUT79), .A3(G91), .A4(new_n507), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n530), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n569), .A2(new_n570), .B1(G651), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n566), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G168), .ZN(G286));
  NAND4_X1  g151(.A1(new_n516), .A2(new_n518), .A3(G49), .A4(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n516), .A2(new_n518), .A3(G87), .A4(new_n507), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G288));
  NAND3_X1  g159(.A1(new_n519), .A2(G48), .A3(G543), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n516), .A2(new_n518), .A3(G86), .A4(new_n507), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n545), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n523), .A2(G47), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n520), .A2(G85), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n545), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n516), .A2(new_n518), .A3(G92), .A4(new_n507), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(KEYINPUT81), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(KEYINPUT81), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n598), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n530), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n523), .A2(G54), .B1(G651), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n595), .B1(new_n608), .B2(G868), .ZN(G284));
  XOR2_X1   g184(.A(G284), .B(KEYINPUT82), .Z(G321));
  NOR2_X1   g185(.A1(G299), .A2(G868), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g187(.A(new_n611), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n608), .B1(new_n614), .B2(G860), .ZN(G148));
  NOR2_X1   g190(.A1(new_n554), .A2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n608), .A2(new_n614), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g195(.A1(new_n479), .A2(G2105), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n466), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n482), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n484), .A2(G123), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n628), .A2(new_n629), .B1(new_n630), .B2(G2105), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n629), .B2(new_n628), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n626), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n625), .A2(new_n634), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT85), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  AOI21_X1  g215(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT86), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(G14), .B1(new_n642), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n642), .B2(new_n649), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT87), .Z(new_n654));
  NOR2_X1   g229(.A1(G2072), .A2(G2078), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n442), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n652), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(KEYINPUT17), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n657), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n652), .B(new_n653), .C1(new_n442), .C2(new_n655), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT18), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n654), .A2(new_n658), .A3(new_n652), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT88), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2100), .ZN(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n671), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  AOI211_X1 g250(.A(new_n673), .B(new_n675), .C1(new_n668), .C2(new_n672), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  INV_X1    g255(.A(G1981), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G229));
  MUX2_X1   g258(.A(G6), .B(G305), .S(G16), .Z(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT91), .Z(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT32), .B(G1981), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT90), .B(G16), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n689), .A2(G22), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1971), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G23), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(G16), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G288), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT33), .ZN(new_n697));
  INV_X1    g272(.A(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n693), .B(new_n699), .C1(new_n686), .C2(new_n685), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G25), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n482), .A2(G131), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n484), .A2(G119), .ZN(new_n706));
  OR2_X1    g281(.A1(G95), .A2(G2105), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n707), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n710), .B2(new_n703), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT35), .B(G1991), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT89), .Z(new_n713));
  OAI21_X1  g288(.A(KEYINPUT92), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(G24), .B(G290), .S(new_n689), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1986), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n714), .B(new_n716), .C1(new_n713), .C2(new_n711), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n701), .A2(new_n702), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n689), .A2(G19), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n554), .B2(new_n689), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT93), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1341), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n703), .A2(G27), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G164), .B2(new_n703), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT97), .B(G2078), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n703), .A2(G35), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G162), .B2(new_n703), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n733));
  INV_X1    g308(.A(G2090), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n732), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n482), .A2(G140), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n484), .A2(G128), .ZN(new_n738));
  NOR2_X1   g313(.A1(G104), .A2(G2105), .ZN(new_n739));
  OAI21_X1  g314(.A(G2104), .B1(new_n465), .B2(G116), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n737), .B(new_n738), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n703), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G2067), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT24), .ZN(new_n748));
  INV_X1    g323(.A(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G160), .B2(new_n703), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(G2084), .ZN(new_n753));
  INV_X1    g328(.A(G28), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(KEYINPUT30), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n754), .B2(KEYINPUT30), .ZN(new_n756));
  OR2_X1    g331(.A1(KEYINPUT31), .A2(G11), .ZN(new_n757));
  NAND2_X1  g332(.A1(KEYINPUT31), .A2(G11), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n755), .A2(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n633), .B2(new_n703), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G2084), .B2(new_n752), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n736), .A2(new_n747), .A3(new_n753), .A4(new_n761), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n726), .A2(new_n730), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n703), .A2(G32), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n482), .A2(G141), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n484), .A2(G129), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT26), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n621), .A2(G105), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n765), .A2(new_n766), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT96), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n764), .B1(new_n777), .B2(new_n703), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT27), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1996), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n688), .A2(G20), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT23), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1956), .Z(new_n784));
  MUX2_X1   g359(.A(G4), .B(new_n607), .S(G16), .Z(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(G1348), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n785), .A2(G1348), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G21), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(G16), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G286), .B2(G16), .ZN(new_n791));
  INV_X1    g366(.A(G1966), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NOR2_X1   g369(.A1(G29), .A2(G33), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT94), .Z(new_n796));
  NAND3_X1  g371(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT25), .Z(new_n798));
  AOI22_X1  g373(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n482), .A2(KEYINPUT95), .A3(G139), .ZN(new_n800));
  AOI21_X1  g375(.A(KEYINPUT95), .B1(new_n482), .B2(G139), .ZN(new_n801));
  OAI221_X1 g376(.A(new_n798), .B1(new_n465), .B2(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(new_n703), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(G2072), .Z(new_n804));
  INV_X1    g379(.A(G5), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(G16), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G301), .B2(G16), .ZN(new_n807));
  INV_X1    g382(.A(G1961), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n793), .A2(new_n794), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n763), .A2(new_n780), .A3(new_n788), .A4(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n721), .A2(new_n722), .A3(new_n811), .ZN(G311));
  INV_X1    g387(.A(G311), .ZN(G150));
  NAND2_X1  g388(.A1(new_n523), .A2(G55), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n520), .A2(G93), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n814), .B(new_n815), .C1(new_n545), .C2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n553), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT38), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n608), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n822), .A2(new_n823), .A3(G860), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n817), .A2(G860), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT37), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n824), .A2(new_n826), .ZN(G145));
  NAND2_X1  g402(.A1(new_n484), .A2(G130), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT99), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n482), .A2(G142), .ZN(new_n830));
  NOR2_X1   g405(.A1(G106), .A2(G2105), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(new_n465), .B2(G118), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n623), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n494), .A2(new_n495), .A3(new_n498), .A4(new_n500), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n802), .B(new_n835), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n834), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n776), .B(new_n741), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n709), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n633), .B(G160), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G162), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n837), .A2(new_n839), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G37), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n842), .B1(new_n840), .B2(new_n843), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT100), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n847), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n849), .A2(new_n850), .A3(new_n845), .A4(new_n844), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(KEYINPUT42), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n818), .B(new_n617), .ZN(new_n857));
  INV_X1    g432(.A(G299), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n607), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n608), .A2(G299), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT101), .B1(new_n608), .B2(G299), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n858), .A2(new_n607), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n865), .A3(new_n860), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT41), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT102), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n866), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT41), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n856), .B(new_n862), .C1(new_n874), .C2(new_n857), .ZN(new_n875));
  INV_X1    g450(.A(new_n872), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n868), .B2(KEYINPUT102), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n857), .B1(new_n877), .B2(new_n871), .ZN(new_n878));
  INV_X1    g453(.A(new_n862), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n855), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G303), .B(G290), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n583), .B(G305), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n854), .B2(KEYINPUT42), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n875), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n875), .B2(new_n880), .ZN(new_n886));
  OAI21_X1  g461(.A(G868), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G868), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n817), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(G295));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n887), .A2(new_n891), .A3(new_n889), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n887), .B2(new_n889), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(G331));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  NAND2_X1  g470(.A1(G301), .A2(KEYINPUT105), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n542), .A2(new_n543), .A3(new_n897), .A4(new_n546), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(G168), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n538), .A2(new_n896), .A3(new_n540), .A4(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n818), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n904), .A2(new_n861), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(new_n818), .A3(new_n901), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n900), .A2(new_n818), .A3(KEYINPUT107), .A4(new_n901), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n904), .A2(new_n906), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n873), .A2(KEYINPUT106), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT106), .B1(new_n873), .B2(new_n911), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n883), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n883), .B(new_n910), .C1(new_n912), .C2(new_n913), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n845), .A4(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n908), .A2(new_n904), .A3(new_n909), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT41), .B1(new_n859), .B2(new_n860), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n863), .A2(new_n865), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n860), .A2(KEYINPUT41), .ZN(new_n923));
  OAI22_X1  g498(.A1(new_n921), .A2(KEYINPUT108), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n921), .A2(KEYINPUT108), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n905), .A2(new_n906), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(G37), .B1(new_n928), .B2(new_n915), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n918), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n895), .B1(new_n919), .B2(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n918), .A2(new_n929), .A3(new_n917), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n916), .A2(new_n845), .A3(new_n918), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(KEYINPUT43), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n895), .B2(new_n935), .ZN(G397));
  INV_X1    g511(.A(KEYINPUT123), .ZN(new_n937));
  INV_X1    g512(.A(G8), .ZN(new_n938));
  NOR2_X1   g513(.A1(G168), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(KEYINPUT51), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n498), .A2(new_n500), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT69), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n498), .A2(KEYINPUT69), .A3(new_n500), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n945), .B2(new_n496), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT50), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT114), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G2084), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n503), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT50), .ZN(new_n953));
  NAND2_X1  g528(.A1(G160), .A2(G40), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n835), .A2(new_n950), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n947), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n948), .A2(new_n949), .A3(new_n953), .A4(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n951), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G40), .ZN(new_n961));
  AOI211_X1 g536(.A(new_n961), .B(new_n469), .C1(new_n480), .C2(new_n465), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n956), .B2(KEYINPUT45), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n792), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n938), .B1(new_n958), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT122), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n940), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI211_X1 g542(.A(KEYINPUT122), .B(new_n938), .C1(new_n958), .C2(new_n964), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n937), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n958), .A2(new_n964), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(G8), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT122), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n965), .A2(new_n966), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n972), .A2(KEYINPUT123), .A3(new_n973), .A4(new_n940), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT51), .B1(new_n965), .B2(new_n939), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n969), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT62), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n970), .A2(new_n939), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n948), .A2(new_n953), .A3(new_n957), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n808), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n960), .A2(new_n963), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G2078), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n962), .B1(new_n959), .B2(new_n955), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT112), .B1(new_n951), .B2(new_n959), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n991), .B(KEYINPUT45), .C1(new_n503), .C2(new_n950), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n989), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n991), .B1(new_n946), .B2(KEYINPUT45), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n951), .A2(KEYINPUT112), .A3(new_n959), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n998), .A2(KEYINPUT113), .A3(new_n989), .ZN(new_n999));
  AOI21_X1  g574(.A(G2078), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n987), .B1(new_n1000), .B2(KEYINPUT53), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G171), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1971), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n995), .A2(new_n999), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n962), .B1(new_n956), .B2(new_n947), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n947), .B2(new_n946), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n734), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n938), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G303), .A2(G8), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT55), .Z(new_n1011));
  NOR2_X1   g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n980), .A2(G2090), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1005), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(G8), .A3(new_n1011), .ZN(new_n1016));
  OAI21_X1  g591(.A(G8), .B1(new_n954), .B2(new_n955), .ZN(new_n1017));
  AOI211_X1 g592(.A(new_n698), .B(new_n579), .C1(new_n581), .C2(new_n582), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n583), .B2(G1976), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(KEYINPUT115), .B(new_n1020), .C1(new_n583), .C2(G1976), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT52), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G305), .A2(G1981), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n585), .A2(new_n588), .A3(new_n681), .A4(new_n586), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT49), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1017), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1027), .A2(KEYINPUT49), .A3(new_n1028), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1025), .A2(new_n1026), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1003), .A2(new_n1013), .A3(new_n1016), .A4(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT125), .B1(new_n979), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1016), .B(new_n1037), .C1(new_n1011), .C2(new_n1009), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(new_n1002), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT125), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n976), .A2(new_n978), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1041), .B(new_n1042), .C1(KEYINPUT62), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(KEYINPUT62), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT126), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1039), .A2(new_n1044), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1016), .A2(new_n1037), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(new_n1012), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT45), .B1(new_n955), .B2(KEYINPUT109), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(KEYINPUT109), .B2(new_n955), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n989), .A2(new_n1053), .A3(new_n984), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n981), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1056), .B(G301), .C1(new_n1000), .C2(KEYINPUT53), .ZN(new_n1057));
  INV_X1    g632(.A(G2078), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT113), .B1(new_n998), .B2(new_n989), .ZN(new_n1059));
  AOI211_X1 g634(.A(new_n994), .B(new_n988), .C1(new_n996), .C2(new_n997), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n986), .B1(new_n1061), .B2(new_n983), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1057), .B1(new_n1062), .B2(G301), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n987), .B(G301), .C1(new_n1000), .C2(KEYINPUT53), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1055), .B1(new_n1061), .B2(new_n983), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1066), .B(KEYINPUT54), .C1(new_n1067), .C2(G301), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1043), .A2(new_n1051), .A3(new_n1065), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT54), .B1(new_n1002), .B2(new_n1057), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(new_n1040), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1073), .A2(KEYINPUT124), .A3(new_n1043), .A4(new_n1068), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT56), .B(G2072), .Z(new_n1075));
  NOR2_X1   g650(.A1(new_n993), .A2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1076), .B(KEYINPUT121), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n858), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(G299), .A2(KEYINPUT120), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1080), .A2(KEYINPUT57), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT119), .B(G1956), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1007), .A2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1077), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1086), .B1(new_n1077), .B2(new_n1089), .ZN(new_n1091));
  INV_X1    g666(.A(G1348), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n954), .A2(new_n955), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n980), .A2(new_n1092), .B1(new_n746), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(new_n607), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1090), .A2(new_n1091), .A3(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT58), .B(G1341), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n993), .A2(G1996), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n554), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT59), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT61), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1094), .A2(new_n607), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT60), .B1(new_n1102), .B2(new_n1095), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1094), .A2(new_n1104), .A3(new_n608), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1100), .A2(KEYINPUT61), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1096), .A2(new_n1106), .B1(new_n1090), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1071), .A2(new_n1074), .A3(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G305), .A2(G1981), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n583), .A2(new_n698), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT116), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI22_X1  g689(.A1(new_n1016), .A2(new_n1035), .B1(new_n1017), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n965), .A2(G168), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT118), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1051), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n938), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1119), .B(new_n1035), .C1(new_n1121), .C2(new_n1011), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1122), .B(new_n1117), .C1(new_n1011), .C2(new_n1121), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1115), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1049), .A2(new_n1109), .A3(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1053), .A2(new_n954), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G290), .A2(G1986), .ZN(new_n1127));
  XOR2_X1   g702(.A(new_n1127), .B(KEYINPUT110), .Z(new_n1128));
  AND2_X1   g703(.A1(G290), .A2(G1986), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT111), .ZN(new_n1131));
  INV_X1    g706(.A(G1996), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n776), .B(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n741), .B(new_n746), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n709), .B(new_n713), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1126), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1131), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1125), .A2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1053), .A2(G1996), .A3(new_n954), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1140), .A2(KEYINPUT46), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(KEYINPUT46), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1134), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1126), .B1(new_n1143), .B2(new_n776), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT47), .Z(new_n1146));
  NAND2_X1  g721(.A1(new_n1128), .A2(new_n1126), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT127), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT48), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1150), .A2(new_n1137), .A3(new_n1151), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n709), .A2(new_n713), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1135), .A2(new_n1153), .B1(G2067), .B2(new_n741), .ZN(new_n1154));
  AOI211_X1 g729(.A(new_n1146), .B(new_n1152), .C1(new_n1126), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1139), .A2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g731(.A1(G229), .A2(new_n463), .A3(G401), .A4(G227), .ZN(new_n1158));
  NAND2_X1  g732(.A1(new_n1158), .A2(new_n852), .ZN(new_n1159));
  NOR2_X1   g733(.A1(new_n935), .A2(new_n1159), .ZN(G308));
  OR2_X1    g734(.A1(new_n935), .A2(new_n1159), .ZN(G225));
endmodule


