//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n631, new_n632, new_n635, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1236, new_n1237, new_n1239;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g047(.A(KEYINPUT67), .B(G125), .C1(new_n463), .C2(new_n464), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n469), .B1(new_n475), .B2(G2105), .ZN(G160));
  NOR2_X1   g051(.A1(new_n463), .A2(new_n464), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(new_n462), .ZN(new_n478));
  MUX2_X1   g053(.A(G100), .B(G112), .S(G2105), .Z(new_n479));
  AOI22_X1  g054(.A1(new_n478), .A2(G124), .B1(G2104), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n477), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n481), .A2(new_n482), .A3(G136), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n481), .B2(G136), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND2_X1  g061(.A1(new_n462), .A2(G102), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n466), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n463), .B2(new_n464), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT69), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(new_n490), .C1(new_n463), .C2(new_n464), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n489), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT3), .B(G2104), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n498), .A2(new_n499), .A3(G138), .A4(new_n462), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n511), .A2(new_n517), .ZN(G166));
  OR2_X1    g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n505), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(G51), .B1(new_n508), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n508), .A2(new_n512), .A3(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n527), .B1(new_n524), .B2(new_n526), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n523), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g107(.A(KEYINPUT71), .B(new_n523), .C1(new_n528), .C2(new_n529), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n510), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n513), .A2(new_n537), .B1(new_n515), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  AND2_X1   g116(.A1(KEYINPUT5), .A2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(KEYINPUT5), .A2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT72), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n548), .B(new_n541), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(G651), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n508), .A2(new_n512), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G81), .B1(G43), .B2(new_n521), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND3_X1  g135(.A1(new_n512), .A2(G53), .A3(G543), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT74), .B1(new_n561), .B2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n521), .A2(new_n563), .A3(new_n564), .A4(G53), .ZN(new_n565));
  AOI211_X1 g140(.A(KEYINPUT73), .B(new_n564), .C1(new_n521), .C2(G53), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n561), .B2(KEYINPUT9), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n562), .B(new_n565), .C1(new_n566), .C2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT75), .B1(new_n513), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n508), .A2(new_n512), .A3(new_n572), .A4(G91), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n506), .B2(new_n507), .ZN(new_n575));
  AND2_X1   g150(.A1(G78), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND3_X1   g152(.A1(new_n571), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n569), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND2_X1  g157(.A1(new_n521), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n513), .ZN(G288));
  AOI22_X1  g161(.A1(new_n551), .A2(G86), .B1(G48), .B2(new_n521), .ZN(new_n587));
  OAI21_X1  g162(.A(G61), .B1(new_n542), .B2(new_n543), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT76), .B1(new_n590), .B2(G651), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n592));
  AOI211_X1 g167(.A(new_n592), .B(new_n510), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n587), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(KEYINPUT77), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n592), .B1(new_n597), .B2(new_n510), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n590), .A2(KEYINPUT76), .A3(G651), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n596), .B1(new_n600), .B2(new_n587), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n595), .A2(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n510), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n508), .A2(new_n512), .A3(G85), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n512), .A2(G47), .A3(G543), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n605), .A2(new_n606), .A3(KEYINPUT78), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT78), .B1(new_n605), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(KEYINPUT79), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n611), .B(new_n604), .C1(new_n607), .C2(new_n608), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n612), .ZN(G290));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n513), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n508), .A2(new_n512), .A3(KEYINPUT10), .A4(G92), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G79), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT80), .B1(new_n619), .B2(new_n505), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n621), .A2(G79), .A3(G543), .ZN(new_n622));
  INV_X1    g197(.A(G66), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n622), .C1(new_n544), .C2(new_n623), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n624), .A2(G651), .B1(G54), .B2(new_n521), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  MUX2_X1   g201(.A(new_n626), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g202(.A(new_n626), .B(G301), .S(G868), .Z(G321));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  OR3_X1    g204(.A1(G168), .A2(KEYINPUT81), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g205(.A1(G168), .A2(new_n629), .ZN(new_n631));
  AOI21_X1  g206(.A(KEYINPUT81), .B1(G299), .B2(new_n629), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(G297));
  OAI21_X1  g208(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(G280));
  INV_X1    g209(.A(new_n626), .ZN(new_n635));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G860), .ZN(G148));
  NOR2_X1   g212(.A1(new_n553), .A2(G868), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n626), .A2(G559), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n638), .B1(G868), .B2(new_n639), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n478), .A2(G123), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT83), .ZN(new_n643));
  MUX2_X1   g218(.A(G99), .B(G111), .S(G2105), .Z(new_n644));
  AOI22_X1  g219(.A1(new_n481), .A2(G135), .B1(G2104), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT84), .B(G2096), .Z(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n481), .A2(G2104), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT13), .B(G2100), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n646), .A2(new_n647), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n648), .A2(new_n653), .A3(new_n654), .ZN(G156));
  INV_X1    g230(.A(KEYINPUT14), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT15), .B(G2435), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2427), .ZN(new_n659));
  INV_X1    g234(.A(G2430), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n656), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n662), .A2(new_n668), .ZN(new_n670));
  AND3_X1   g245(.A1(new_n669), .A2(G14), .A3(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  INV_X1    g253(.A(new_n674), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n679), .A2(KEYINPUT17), .A3(new_n672), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n672), .B1(new_n679), .B2(KEYINPUT17), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n676), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n673), .A2(new_n676), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n679), .B1(new_n683), .B2(KEYINPUT17), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n678), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G2096), .Z(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(G2100), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n690), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n690), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n701), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(G229));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(G23), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G288), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(G22), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT85), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G166), .B2(new_n707), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(G1971), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(G1971), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n711), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT32), .B(G1981), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n594), .A2(KEYINPUT77), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n600), .A2(new_n596), .A3(new_n587), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n707), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G6), .A2(G16), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n718), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n718), .ZN(new_n726));
  NOR3_X1   g301(.A1(new_n721), .A2(new_n723), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n717), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(KEYINPUT34), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n717), .B(new_n730), .C1(new_n725), .C2(new_n727), .ZN(new_n731));
  NOR2_X1   g306(.A1(G25), .A2(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n481), .A2(G131), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n478), .A2(G119), .ZN(new_n734));
  MUX2_X1   g309(.A(G95), .B(G107), .S(G2105), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G2104), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n732), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n610), .A2(new_n612), .A3(G16), .ZN(new_n742));
  OR2_X1    g317(.A1(G16), .A2(G24), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n742), .A2(G1986), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(G1986), .B1(new_n742), .B2(new_n743), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AND3_X1   g322(.A1(new_n731), .A2(new_n747), .A3(KEYINPUT86), .ZN(new_n748));
  AOI21_X1  g323(.A(KEYINPUT86), .B1(new_n731), .B2(new_n747), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n729), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(KEYINPUT36), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(KEYINPUT36), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n731), .A2(new_n747), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT86), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n731), .A2(new_n747), .A3(KEYINPUT86), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n759), .A2(new_n751), .A3(KEYINPUT36), .A4(new_n729), .ZN(new_n760));
  NOR2_X1   g335(.A1(G16), .A2(G19), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n554), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT88), .B(G1341), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(G162), .A2(G29), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G29), .B2(G35), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT29), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n764), .B1(new_n768), .B2(G2090), .ZN(new_n769));
  INV_X1    g344(.A(G29), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n770), .A2(G33), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n467), .A2(G103), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT25), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n498), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n774));
  AND3_X1   g349(.A1(new_n481), .A2(KEYINPUT90), .A3(G139), .ZN(new_n775));
  AOI21_X1  g350(.A(KEYINPUT90), .B1(new_n481), .B2(G139), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n773), .B1(new_n462), .B2(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n771), .B1(new_n777), .B2(G29), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G2072), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n770), .A2(G32), .ZN(new_n780));
  AOI22_X1  g355(.A1(G129), .A2(new_n478), .B1(new_n481), .B2(G141), .ZN(new_n781));
  NAND3_X1  g356(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT26), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n784), .A2(new_n785), .B1(G105), .B2(new_n467), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n781), .A2(KEYINPUT93), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n780), .B1(new_n792), .B2(new_n770), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT27), .B(G1996), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G34), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n770), .B1(new_n796), .B2(G34), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n799), .B2(new_n798), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G29), .B2(G160), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n793), .A2(new_n795), .B1(G2084), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n793), .A2(new_n795), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n779), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n770), .A2(G26), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT28), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n481), .A2(G140), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n478), .A2(G128), .ZN(new_n809));
  MUX2_X1   g384(.A(G104), .B(G116), .S(G2105), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G2104), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(G29), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n813), .A2(KEYINPUT89), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(KEYINPUT89), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n807), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2067), .ZN(new_n817));
  INV_X1    g392(.A(G2090), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n767), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n635), .A2(G16), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G4), .B2(G16), .ZN(new_n821));
  INV_X1    g396(.A(G1348), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(G164), .A2(G29), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G27), .B2(G29), .ZN(new_n825));
  INV_X1    g400(.A(G2078), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n821), .A2(new_n822), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n825), .A2(new_n826), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n823), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(G171), .A2(new_n707), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G5), .B2(new_n707), .ZN(new_n832));
  INV_X1    g407(.A(G1961), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n802), .A2(G2084), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n833), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n646), .A2(new_n770), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT31), .B(G11), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT94), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT30), .B(G28), .Z(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(G29), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n830), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n769), .A2(new_n805), .A3(new_n819), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(G16), .A2(G21), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G168), .B2(G16), .ZN(new_n847));
  INV_X1    g422(.A(G1966), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n707), .A2(G20), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT23), .Z(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G299), .B2(G16), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(G1956), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n845), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n754), .A2(new_n760), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(G311));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n856), .B(new_n858), .ZN(G150));
  AOI22_X1  g434(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n510), .ZN(new_n861));
  INV_X1    g436(.A(G93), .ZN(new_n862));
  INV_X1    g437(.A(G55), .ZN(new_n863));
  OAI22_X1  g438(.A1(new_n513), .A2(new_n862), .B1(new_n515), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G860), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT37), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n553), .B(new_n865), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n626), .A2(new_n636), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(KEYINPUT96), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n875), .B(new_n866), .C1(new_n873), .C2(new_n872), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(KEYINPUT96), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n868), .B1(new_n876), .B2(new_n877), .ZN(G145));
  AOI22_X1  g453(.A1(G130), .A2(new_n478), .B1(new_n481), .B2(G142), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n880), .A2(KEYINPUT97), .ZN(new_n881));
  OAI22_X1  g456(.A1(new_n880), .A2(KEYINPUT97), .B1(G118), .B2(new_n462), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n737), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n651), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n791), .B(new_n812), .Z(new_n886));
  OR2_X1    g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n777), .B(new_n502), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n887), .B2(new_n888), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n646), .B(G160), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G162), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n894), .A2(G37), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n890), .B2(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(KEYINPUT98), .B(KEYINPUT40), .Z(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(G395));
  AND3_X1   g477(.A1(new_n610), .A2(new_n612), .A3(G288), .ZN(new_n903));
  AOI21_X1  g478(.A(G288), .B1(new_n610), .B2(new_n612), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(G166), .B1(new_n595), .B2(new_n601), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n719), .A2(new_n720), .A3(G303), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT101), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n910));
  INV_X1    g485(.A(G288), .ZN(new_n911));
  NAND2_X1  g486(.A1(G290), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n610), .A2(new_n612), .A3(G288), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n719), .A2(new_n720), .A3(G303), .ZN(new_n915));
  AOI21_X1  g490(.A(G303), .B1(new_n719), .B2(new_n720), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n910), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  OAI22_X1  g493(.A1(new_n909), .A2(new_n918), .B1(new_n917), .B2(new_n914), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n569), .A2(new_n626), .A3(new_n578), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT100), .ZN(new_n921));
  NAND2_X1  g496(.A1(G299), .A2(new_n635), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n569), .A2(new_n626), .A3(new_n924), .A4(new_n578), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n921), .A2(new_n922), .A3(new_n923), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n920), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n928), .B2(new_n923), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n639), .A2(KEYINPUT99), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT99), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n626), .B2(G559), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n865), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(new_n553), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n869), .A2(new_n932), .A3(new_n930), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n929), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n928), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(KEYINPUT42), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT42), .B1(new_n938), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n919), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n938), .A2(new_n940), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT101), .B1(new_n905), .B2(new_n908), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n914), .A2(new_n917), .A3(new_n910), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n948), .A2(new_n949), .B1(new_n908), .B2(new_n905), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n941), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n629), .B1(new_n944), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n934), .A2(G868), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(G295));
  NAND2_X1  g529(.A1(new_n944), .A2(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(G868), .ZN(new_n956));
  INV_X1    g531(.A(new_n953), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT102), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n952), .A2(new_n959), .A3(new_n953), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n958), .A2(new_n960), .ZN(G331));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n532), .A2(new_n533), .A3(G301), .ZN(new_n963));
  AOI21_X1  g538(.A(G301), .B1(new_n532), .B2(new_n533), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n935), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(G168), .A2(G171), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n532), .A2(new_n533), .A3(G301), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n869), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n968), .A3(new_n927), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n965), .A2(new_n968), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n970), .B(new_n926), .C1(new_n923), .C2(new_n928), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n919), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n965), .A2(new_n968), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n969), .B1(new_n973), .B2(new_n929), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n950), .ZN(new_n975));
  INV_X1    g550(.A(G37), .ZN(new_n976));
  XNOR2_X1  g551(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n972), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n978), .A2(KEYINPUT44), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n969), .A2(KEYINPUT106), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n965), .A2(new_n968), .A3(new_n981), .A4(new_n927), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n626), .B1(new_n569), .B2(new_n578), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(KEYINPUT100), .B2(new_n920), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT41), .A4(new_n925), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT41), .A4(new_n925), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT105), .ZN(new_n989));
  INV_X1    g564(.A(new_n920), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n923), .B1(new_n990), .B2(new_n984), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n927), .A2(KEYINPUT104), .A3(new_n923), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n987), .A2(new_n989), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n970), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n919), .B1(new_n983), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n976), .B1(new_n974), .B2(new_n950), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT43), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n962), .B1(new_n979), .B2(new_n999), .ZN(new_n1000));
  AND4_X1   g575(.A1(new_n962), .A2(new_n999), .A3(KEYINPUT44), .A4(new_n978), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n977), .B1(new_n997), .B2(new_n998), .ZN(new_n1002));
  INV_X1    g577(.A(new_n977), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n972), .A2(new_n975), .A3(new_n976), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  OAI22_X1  g580(.A1(new_n1000), .A2(new_n1001), .B1(KEYINPUT44), .B2(new_n1005), .ZN(G397));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n502), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1384), .B1(new_n495), .B2(new_n501), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT108), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT45), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G40), .ZN(new_n1014));
  AOI211_X1 g589(.A(new_n1014), .B(new_n469), .C1(new_n475), .C2(G2105), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  XOR2_X1   g592(.A(new_n737), .B(new_n740), .Z(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT109), .ZN(new_n1019));
  INV_X1    g594(.A(G1996), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n812), .B(G2067), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n791), .B2(G1996), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(G290), .B(G1986), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1017), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1008), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1028), .A2(new_n826), .A3(new_n1015), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT124), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n473), .A2(new_n474), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT67), .B1(new_n498), .B2(G125), .ZN(new_n1033));
  OAI21_X1  g608(.A(G2105), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n469), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(G40), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n1008), .B2(new_n1027), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT124), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n826), .A4(new_n1029), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1031), .A2(KEYINPUT53), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT50), .B1(new_n502), .B2(new_n1007), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n1042), .B(G1384), .C1(new_n495), .C2(new_n501), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1015), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT119), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(new_n1015), .C1(new_n1041), .C2(new_n1043), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n833), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1029), .A2(KEYINPUT110), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1011), .A2(new_n1051), .A3(KEYINPUT45), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1037), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1049), .B1(new_n1053), .B2(G2078), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1040), .A2(new_n1048), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G171), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT125), .B1(new_n1013), .B2(new_n1036), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1011), .A2(KEYINPUT108), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1009), .B(G1384), .C1(new_n495), .C2(new_n501), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1027), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT125), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1015), .ZN(new_n1062));
  AND4_X1   g637(.A1(KEYINPUT53), .A2(new_n1050), .A3(new_n826), .A4(new_n1052), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1057), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1064), .A2(G301), .A3(new_n1048), .A4(new_n1054), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1056), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G288), .A2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT112), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n1072));
  INV_X1    g647(.A(G8), .ZN(new_n1073));
  AOI211_X1 g648(.A(new_n1072), .B(new_n1073), .C1(new_n1015), .C2(new_n1011), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1011), .A2(G40), .A3(G160), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT111), .B1(new_n1075), .B2(G8), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1071), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(KEYINPUT113), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n1008), .B2(new_n1036), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1072), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1075), .A2(KEYINPUT111), .A3(G8), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(new_n1071), .A3(new_n1079), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n911), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1081), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n1092));
  INV_X1    g667(.A(G1981), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n600), .B2(new_n587), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n1095));
  INV_X1    g670(.A(G86), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1095), .B1(new_n513), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g672(.A(G1981), .B(new_n1097), .C1(new_n598), .C2(new_n599), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1092), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n594), .A2(G1981), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n600), .A2(new_n1093), .A3(new_n587), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1101), .A3(KEYINPUT49), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1090), .B1(new_n1091), .B2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1085), .A2(KEYINPUT114), .A3(new_n1102), .A4(new_n1099), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(G303), .A2(G8), .ZN(new_n1107));
  XOR2_X1   g682(.A(new_n1107), .B(KEYINPUT55), .Z(new_n1108));
  INV_X1    g683(.A(G1971), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1053), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n818), .B(new_n1015), .C1(new_n1041), .C2(new_n1043), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1108), .B(G8), .C1(new_n1110), .C2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1107), .B(KEYINPUT55), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1008), .A2(new_n1042), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1036), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1053), .A2(new_n1109), .B1(new_n1117), .B2(new_n818), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1114), .B1(new_n1118), .B2(new_n1073), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1089), .A2(new_n1106), .A3(new_n1113), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1057), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1048), .A2(new_n1054), .ZN(new_n1123));
  OAI21_X1  g698(.A(G171), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1040), .A2(G301), .A3(new_n1048), .A4(new_n1054), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(KEYINPUT54), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT51), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1037), .A2(new_n1029), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n848), .ZN(new_n1129));
  INV_X1    g704(.A(G2084), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1117), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1131), .A3(G168), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1073), .A2(KEYINPUT123), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1127), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1127), .A3(new_n1133), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(G8), .A3(G286), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1068), .A2(new_n1121), .A3(new_n1126), .A4(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(KEYINPUT116), .B(G1956), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1044), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT56), .B(G2072), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1037), .A2(new_n1050), .A3(new_n1052), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1146));
  NAND2_X1  g721(.A1(G299), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1146), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n569), .A2(new_n578), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1145), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1045), .A2(new_n822), .A3(new_n1047), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1075), .A2(G2067), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1152), .B1(new_n1155), .B2(new_n626), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1142), .A2(new_n1144), .A3(new_n1150), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT118), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT118), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1142), .A2(new_n1144), .A3(new_n1150), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1156), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT61), .B1(new_n1161), .B2(new_n1152), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1037), .A2(new_n1050), .A3(new_n1020), .A4(new_n1052), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT58), .B(G1341), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT121), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1075), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1171));
  OAI211_X1 g746(.A(KEYINPUT59), .B(new_n554), .C1(new_n1167), .C2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1152), .A2(KEYINPUT61), .A3(new_n1157), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1175), .A2(KEYINPUT120), .A3(new_n1020), .A4(new_n1037), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1176), .A2(new_n1166), .A3(new_n1170), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT59), .B1(new_n1177), .B2(new_n554), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1163), .A2(new_n1174), .A3(new_n1178), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1153), .A2(KEYINPUT60), .A3(new_n626), .A4(new_n1154), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(KEYINPUT122), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1153), .A2(KEYINPUT60), .A3(new_n1154), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n635), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1180), .A2(KEYINPUT122), .ZN(new_n1185));
  OAI22_X1  g760(.A1(new_n1184), .A2(new_n1185), .B1(KEYINPUT60), .B2(new_n1155), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1140), .B1(new_n1162), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT63), .ZN(new_n1189));
  NOR2_X1   g764(.A1(G286), .A2(new_n1073), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1137), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1189), .B1(new_n1120), .B2(new_n1191), .ZN(new_n1192));
  XOR2_X1   g767(.A(new_n1070), .B(KEYINPUT112), .Z(new_n1193));
  AOI21_X1  g768(.A(new_n1193), .B1(new_n1084), .B2(new_n1083), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1087), .B1(new_n1194), .B2(new_n1079), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1195), .A2(new_n1081), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT115), .B1(new_n1196), .B2(new_n1119), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1118), .A2(new_n1073), .A3(new_n1114), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1198), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1089), .A2(new_n1106), .A3(KEYINPUT115), .A4(new_n1119), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1192), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1106), .A2(new_n1069), .A3(new_n911), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n1101), .ZN(new_n1204));
  AOI22_X1  g779(.A1(new_n1204), .A2(new_n1085), .B1(new_n1198), .B2(new_n1196), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1206));
  OAI21_X1  g781(.A(KEYINPUT62), .B1(new_n1206), .B2(new_n1134), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT62), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1135), .A2(new_n1208), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1056), .ZN(new_n1210));
  NAND4_X1  g785(.A1(new_n1207), .A2(new_n1209), .A3(new_n1121), .A4(new_n1210), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1202), .A2(new_n1205), .A3(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1026), .B1(new_n1188), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n1214));
  OAI211_X1 g789(.A(new_n1017), .B(new_n1020), .C1(new_n1214), .C2(KEYINPUT46), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1214), .A2(KEYINPUT46), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n1215), .B(new_n1216), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1017), .B1(new_n791), .B2(new_n1022), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1218), .B(KEYINPUT127), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n1220), .B(KEYINPUT47), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n738), .A2(new_n740), .ZN(new_n1223));
  OAI22_X1  g798(.A1(new_n1222), .A2(new_n1223), .B1(G2067), .B2(new_n812), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1224), .A2(new_n1017), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1024), .A2(new_n1017), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT48), .ZN(new_n1227));
  OR3_X1    g802(.A1(new_n1016), .A2(G1986), .A3(G290), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1226), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g804(.A(new_n1228), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1230), .A2(KEYINPUT48), .ZN(new_n1231));
  OAI21_X1  g806(.A(new_n1225), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1221), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1213), .A2(new_n1233), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g809(.A1(G401), .A2(new_n460), .ZN(new_n1236));
  NAND3_X1  g810(.A1(new_n1236), .A2(new_n687), .A3(new_n705), .ZN(new_n1237));
  AOI211_X1 g811(.A(new_n1237), .B(new_n1005), .C1(new_n896), .C2(new_n895), .ZN(G308));
  AOI21_X1  g812(.A(new_n1237), .B1(new_n895), .B2(new_n896), .ZN(new_n1239));
  NAND3_X1  g813(.A1(new_n1239), .A2(new_n1002), .A3(new_n1004), .ZN(G225));
endmodule


