//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  NAND2_X1  g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT96), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT14), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n206), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n212), .A2(KEYINPUT95), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT95), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n209), .A2(new_n211), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n203), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT17), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n221), .A2(G1gat), .ZN(new_n222));
  AOI21_X1  g021(.A(G8gat), .B1(new_n222), .B2(KEYINPUT97), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n223), .B(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n219), .A2(KEYINPUT17), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n220), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n227), .ZN(new_n231));
  INV_X1    g030(.A(new_n219), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT98), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n237), .B1(new_n227), .B2(new_n219), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n230), .B(KEYINPUT13), .Z(new_n240));
  NAND3_X1  g039(.A1(new_n231), .A2(new_n237), .A3(new_n232), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n234), .A2(new_n235), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n236), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT94), .ZN(new_n246));
  XNOR2_X1  g045(.A(G169gat), .B(G197gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT12), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n244), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n236), .A2(new_n251), .A3(new_n242), .A4(new_n243), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G78gat), .B(G106gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT31), .B(G50gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G22gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT22), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT74), .B(G218gat), .ZN(new_n263));
  INV_X1    g062(.A(G211gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G197gat), .B(G204gat), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n261), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n266), .A3(new_n261), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(G155gat), .A2(G162gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274));
  INV_X1    g073(.A(G141gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(G148gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT77), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n273), .A2(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G148gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G141gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n275), .A2(G148gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT77), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n279), .A2(G141gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n272), .B1(new_n276), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n274), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(new_n271), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n278), .A2(new_n282), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT3), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT29), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n270), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G228gat), .A2(G233gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293));
  INV_X1    g092(.A(new_n269), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(new_n267), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n288), .ZN(new_n296));
  INV_X1    g095(.A(G155gat), .ZN(new_n297));
  INV_X1    g096(.A(G162gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n274), .B1(new_n299), .B2(KEYINPUT2), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n277), .A2(new_n279), .A3(G141gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n282), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G141gat), .B(G148gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n286), .B1(new_n303), .B2(KEYINPUT2), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n302), .A2(KEYINPUT78), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT78), .B1(new_n302), .B2(new_n304), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n287), .B1(new_n295), .B2(new_n288), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n291), .B1(new_n310), .B2(new_n290), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n260), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n259), .B1(new_n312), .B2(KEYINPUT85), .ZN(new_n313));
  INV_X1    g112(.A(new_n291), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT77), .ZN(new_n315));
  NOR3_X1   g114(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n301), .B1(new_n316), .B2(new_n285), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT2), .B1(new_n280), .B2(new_n281), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n274), .ZN(new_n319));
  OAI22_X1  g118(.A1(new_n315), .A2(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n296), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n270), .A2(new_n289), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n314), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n314), .B1(new_n270), .B2(new_n289), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n324), .B1(new_n296), .B2(new_n307), .ZN(new_n325));
  OAI21_X1  g124(.A(G22gat), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n311), .A3(new_n260), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT85), .A4(new_n259), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G1gat), .B(G29gat), .Z(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT83), .ZN(new_n333));
  XOR2_X1   g132(.A(G57gat), .B(G85gat), .Z(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT86), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341));
  INV_X1    g140(.A(G134gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G127gat), .ZN(new_n343));
  INV_X1    g142(.A(G127gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G134gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G113gat), .B(G120gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n346), .B1(new_n347), .B2(KEYINPUT1), .ZN(new_n348));
  INV_X1    g147(.A(G120gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G113gat), .ZN(new_n350));
  INV_X1    g149(.A(G113gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G120gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT1), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n348), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n287), .A3(KEYINPUT80), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n302), .A2(new_n304), .A3(new_n348), .A4(new_n356), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n341), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n359), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(KEYINPUT4), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n356), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n320), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n302), .A2(new_n304), .A3(KEYINPUT78), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT3), .A4(new_n370), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n305), .A2(new_n306), .A3(new_n288), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT79), .B1(new_n287), .B2(new_n288), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n366), .B(new_n371), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n340), .B1(new_n365), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT39), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n339), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT87), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT87), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n339), .A2(new_n380), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n368), .A2(new_n370), .A3(new_n366), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(new_n361), .A3(new_n358), .ZN(new_n384));
  INV_X1    g183(.A(new_n340), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT39), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n386), .B2(KEYINPUT39), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n388), .A2(new_n389), .A3(new_n375), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n382), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT40), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT75), .ZN(new_n395));
  INV_X1    g194(.A(G190gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT68), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT68), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G190gat), .ZN(new_n399));
  INV_X1    g198(.A(G183gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT27), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT27), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(G183gat), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n397), .A2(new_n399), .A3(new_n401), .A4(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT28), .B1(new_n404), .B2(KEYINPUT69), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT26), .ZN(new_n408));
  INV_X1    g207(.A(G169gat), .ZN(new_n409));
  INV_X1    g208(.A(G176gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n412));
  AND3_X1   g211(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n411), .B(new_n412), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT70), .ZN(new_n416));
  NAND2_X1  g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n415), .B2(new_n417), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n406), .B(new_n407), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT64), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT24), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n400), .A2(new_n396), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n423), .A2(new_n424), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(G169gat), .A2(G176gat), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT65), .B1(new_n429), .B2(KEYINPUT23), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT65), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT23), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n431), .B(new_n432), .C1(G169gat), .C2(G176gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT66), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n437), .A2(new_n438), .B1(KEYINPUT23), .B2(new_n429), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n428), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT25), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n429), .A2(KEYINPUT23), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n414), .B2(new_n413), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT67), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n446), .A2(new_n421), .A3(new_n426), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n441), .B1(new_n430), .B2(new_n433), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n443), .B(new_n449), .C1(new_n414), .C2(new_n413), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n445), .A2(new_n447), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n442), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT29), .B1(new_n420), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G226gat), .ZN(new_n454));
  INV_X1    g253(.A(G233gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n395), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n456), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n415), .A2(new_n417), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT70), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n407), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(new_n405), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n462), .A2(new_n464), .B1(new_n442), .B2(new_n451), .ZN(new_n465));
  OAI211_X1 g264(.A(KEYINPUT75), .B(new_n458), .C1(new_n465), .C2(KEYINPUT29), .ZN(new_n466));
  INV_X1    g265(.A(new_n270), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n420), .A2(new_n452), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n468), .B2(new_n456), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n457), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n456), .B1(new_n468), .B2(new_n293), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n465), .A2(new_n458), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G8gat), .B(G36gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(G64gat), .B(G92gat), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n475), .B(new_n476), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n470), .A2(new_n473), .A3(new_n477), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT76), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n481), .B2(new_n480), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n483), .A3(new_n480), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT81), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n358), .A2(new_n361), .A3(new_n341), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n385), .B1(new_n363), .B2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n373), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n368), .A2(new_n370), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(new_n288), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n371), .A2(new_n366), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n384), .A2(new_n385), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n488), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n373), .B1(new_n307), .B2(KEYINPUT3), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n371), .A2(new_n366), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n489), .B(new_n490), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n384), .B2(new_n385), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(KEYINPUT81), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n500), .A2(new_n501), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT80), .B1(new_n357), .B2(new_n287), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n359), .A2(new_n360), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT4), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n364), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n385), .A2(KEYINPUT5), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT84), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n512), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n362), .A2(new_n364), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT84), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n374), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n339), .B1(new_n506), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n487), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n382), .A2(KEYINPUT40), .A3(new_n391), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n394), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n478), .B1(new_n474), .B2(KEYINPUT37), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(KEYINPUT38), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT90), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n457), .A2(new_n466), .ZN(new_n528));
  INV_X1    g327(.A(new_n472), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n270), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n471), .A2(new_n472), .ZN(new_n531));
  OAI22_X1  g330(.A1(new_n530), .A2(KEYINPUT89), .B1(new_n467), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(KEYINPUT89), .B2(new_n530), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT37), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n527), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n531), .A2(new_n467), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n528), .A2(new_n529), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n467), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n539), .B2(new_n538), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(KEYINPUT90), .A3(KEYINPUT37), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n526), .B1(new_n535), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n502), .A2(KEYINPUT81), .A3(new_n504), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT81), .B1(new_n502), .B2(new_n504), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n519), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n337), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(KEYINPUT6), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT6), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n544), .A2(new_n545), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n516), .A2(new_n517), .A3(new_n374), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n517), .B1(new_n516), .B2(new_n374), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n337), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n549), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n548), .B1(new_n554), .B2(new_n520), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n534), .B1(new_n470), .B2(new_n473), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT38), .B1(new_n524), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n481), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n331), .B(new_n523), .C1(new_n543), .C2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n366), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n357), .A2(KEYINPUT71), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n468), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G227gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(new_n455), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n420), .A2(new_n452), .A3(new_n562), .A4(new_n366), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT33), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G15gat), .B(G43gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT72), .ZN(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G99gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT73), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n565), .A2(new_n568), .ZN(new_n579));
  INV_X1    g378(.A(new_n567), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT34), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT34), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n578), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n569), .A2(KEYINPUT32), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n576), .B1(new_n569), .B2(new_n570), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n583), .B1(new_n579), .B2(new_n580), .ZN(new_n589));
  AOI211_X1 g388(.A(KEYINPUT34), .B(new_n567), .C1(new_n565), .C2(new_n568), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n585), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n587), .B1(new_n585), .B2(new_n591), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT36), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n594), .A2(KEYINPUT36), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n477), .B1(new_n470), .B2(new_n473), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n470), .A2(new_n473), .A3(new_n477), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(KEYINPUT30), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n481), .A2(new_n483), .A3(new_n480), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n601), .B2(new_n484), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n546), .A2(new_n547), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n506), .A2(new_n519), .A3(new_n337), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n549), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n602), .B1(new_n605), .B2(new_n548), .ZN(new_n606));
  OAI22_X1  g405(.A1(new_n596), .A2(new_n597), .B1(new_n331), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n561), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT91), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n592), .B2(new_n593), .ZN(new_n611));
  INV_X1    g410(.A(new_n591), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n586), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n585), .A2(new_n587), .A3(new_n591), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(KEYINPUT91), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT35), .B1(new_n329), .B2(new_n330), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n555), .A2(new_n487), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT35), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n614), .A2(new_n331), .A3(new_n615), .ZN(new_n623));
  AOI211_X1 g422(.A(KEYINPUT92), .B(new_n622), .C1(new_n606), .C2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT92), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n337), .B1(new_n506), .B2(new_n519), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n548), .B1(new_n554), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n594), .A2(new_n627), .A3(new_n331), .A4(new_n487), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n625), .B1(new_n628), .B2(KEYINPUT35), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n621), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n256), .B1(new_n609), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G85gat), .A2(G92gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT7), .ZN(new_n633));
  NAND2_X1  g432(.A1(G99gat), .A2(G106gat), .ZN(new_n634));
  INV_X1    g433(.A(G85gat), .ZN(new_n635));
  INV_X1    g434(.A(G92gat), .ZN(new_n636));
  AOI22_X1  g435(.A1(KEYINPUT8), .A2(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G99gat), .B(G106gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n220), .A2(new_n228), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G190gat), .B(G218gat), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n640), .ZN(new_n644));
  AND2_X1   g443(.A1(G232gat), .A2(G233gat), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n232), .A2(new_n644), .B1(KEYINPUT41), .B2(new_n645), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n641), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n643), .B1(new_n641), .B2(new_n646), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n645), .A2(KEYINPUT41), .ZN(new_n649));
  XNOR2_X1  g448(.A(G134gat), .B(G162gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  OR3_X1    g451(.A1(new_n647), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n652), .B1(new_n647), .B2(new_n648), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(G71gat), .B(G78gat), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G57gat), .B(G64gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT99), .Z(new_n660));
  AOI21_X1  g459(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n658), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n661), .B(KEYINPUT100), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT101), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n657), .A2(new_n659), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT102), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n666), .A2(new_n668), .A3(new_n672), .A4(new_n669), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n664), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT103), .B(KEYINPUT21), .Z(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(G231gat), .A2(G233gat), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G127gat), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n231), .B1(new_n674), .B2(KEYINPUT21), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n679), .A2(new_n344), .A3(new_n680), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n682), .B2(new_n685), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(new_n297), .ZN(new_n690));
  XNOR2_X1  g489(.A(G183gat), .B(G211gat), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n690), .B(new_n691), .Z(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n687), .A2(new_n688), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n687), .B2(new_n688), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n656), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697));
  XNOR2_X1  g496(.A(G120gat), .B(G148gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(G176gat), .B(G204gat), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n698), .B(new_n699), .Z(new_n700));
  NAND2_X1  g499(.A1(G230gat), .A2(G233gat), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n674), .A2(new_n644), .ZN(new_n703));
  AOI211_X1 g502(.A(new_n640), .B(new_n664), .C1(new_n671), .C2(new_n673), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT104), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n707), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n671), .A2(new_n673), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n640), .B1(new_n711), .B2(new_n664), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT10), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n674), .A2(new_n644), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n704), .A2(KEYINPUT10), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n702), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n700), .B1(new_n710), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n700), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n709), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n697), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n721), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n720), .B1(new_n709), .B2(new_n717), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(KEYINPUT105), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n631), .A2(new_n696), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n627), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n731), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g531(.A1(new_n730), .A2(new_n487), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT16), .B(G8gat), .Z(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(KEYINPUT42), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT107), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n733), .A2(KEYINPUT106), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(KEYINPUT106), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n737), .A2(G8gat), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n734), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n737), .B2(new_n738), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n736), .B(new_n739), .C1(new_n741), .C2(KEYINPUT42), .ZN(G1325gat));
  NOR2_X1   g541(.A1(new_n596), .A2(new_n597), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G15gat), .B1(new_n730), .B2(new_n744), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n617), .A2(G15gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n730), .B2(new_n746), .ZN(G1326gat));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n331), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT108), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT43), .B(G22gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1327gat));
  AND2_X1   g550(.A1(new_n609), .A2(new_n630), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n694), .A2(new_n695), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n728), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n255), .ZN(new_n755));
  OR3_X1    g554(.A1(new_n752), .A2(new_n655), .A3(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n756), .A2(G29gat), .A3(new_n627), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT45), .Z(new_n758));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n533), .A2(new_n527), .A3(new_n534), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT90), .B1(new_n541), .B2(KEYINPUT37), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n525), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n559), .ZN(new_n763));
  INV_X1    g562(.A(new_n331), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT40), .B1(new_n382), .B2(new_n391), .ZN(new_n765));
  AOI211_X1 g564(.A(new_n393), .B(new_n390), .C1(new_n379), .C2(new_n381), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n764), .B1(new_n767), .B2(new_n521), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n607), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n630), .A2(KEYINPUT109), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n627), .A2(new_n487), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n614), .A2(new_n331), .A3(new_n615), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT35), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT92), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n628), .A2(new_n625), .A3(KEYINPUT35), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n777), .A3(new_n621), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n769), .B1(new_n770), .B2(new_n778), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n653), .A2(KEYINPUT110), .A3(new_n654), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT110), .B1(new_n653), .B2(new_n654), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(KEYINPUT44), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n759), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n777), .B1(new_n776), .B2(new_n621), .ZN(new_n786));
  AOI211_X1 g585(.A(KEYINPUT109), .B(new_n620), .C1(new_n774), .C2(new_n775), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n609), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(KEYINPUT111), .A3(new_n783), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT44), .B1(new_n752), .B2(new_n655), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n785), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n755), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G29gat), .B1(new_n793), .B2(new_n627), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n758), .A2(new_n794), .ZN(G1328gat));
  OAI21_X1  g594(.A(G36gat), .B1(new_n793), .B2(new_n487), .ZN(new_n796));
  AOI21_X1  g595(.A(G36gat), .B1(KEYINPUT112), .B2(KEYINPUT46), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n656), .A2(new_n602), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n631), .A2(new_n754), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(G1329gat));
  NAND3_X1  g601(.A1(new_n791), .A2(new_n743), .A3(new_n792), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT113), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n791), .A2(new_n805), .A3(new_n743), .A4(new_n792), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(G43gat), .A3(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n756), .A2(G43gat), .A3(new_n617), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n803), .A2(G43gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n809), .B1(new_n812), .B2(new_n808), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1330gat));
  NAND2_X1  g613(.A1(new_n764), .A2(G50gat), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n756), .A2(new_n331), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n793), .A2(new_n815), .B1(G50gat), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g617(.A1(new_n256), .A2(new_n788), .A3(new_n696), .A4(new_n728), .ZN(new_n819));
  INV_X1    g618(.A(new_n627), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n602), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n824));
  XOR2_X1   g623(.A(KEYINPUT49), .B(G64gat), .Z(new_n825));
  OAI21_X1  g624(.A(new_n824), .B1(new_n823), .B2(new_n825), .ZN(G1333gat));
  INV_X1    g625(.A(G71gat), .ZN(new_n827));
  INV_X1    g626(.A(new_n617), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n819), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n819), .A2(new_n743), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(new_n827), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n831), .B(new_n832), .ZN(G1334gat));
  NAND2_X1  g632(.A1(new_n819), .A2(new_n764), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(G78gat), .ZN(G1335gat));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n729), .A2(new_n255), .A3(new_n753), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n791), .A2(new_n820), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G85gat), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n841));
  INV_X1    g640(.A(new_n753), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n256), .A3(new_n656), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n841), .B1(new_n779), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n843), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n788), .A2(new_n845), .A3(KEYINPUT51), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n728), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n820), .A2(new_n635), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n836), .B1(new_n840), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n839), .B(KEYINPUT114), .C1(new_n848), .C2(new_n849), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1336gat));
  NAND3_X1  g652(.A1(new_n791), .A2(new_n602), .A3(new_n837), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n791), .A2(KEYINPUT116), .A3(new_n602), .A4(new_n837), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(G92gat), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n848), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n487), .A2(G92gat), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT52), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n854), .A2(G92gat), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n844), .A2(KEYINPUT115), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n844), .A2(new_n846), .A3(KEYINPUT115), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n728), .A2(new_n860), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT52), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n862), .A2(new_n868), .ZN(G1337gat));
  AND3_X1   g668(.A1(new_n791), .A2(new_n743), .A3(new_n837), .ZN(new_n870));
  XOR2_X1   g669(.A(KEYINPUT117), .B(G99gat), .Z(new_n871));
  NAND2_X1  g670(.A1(new_n828), .A2(new_n871), .ZN(new_n872));
  OAI22_X1  g671(.A1(new_n870), .A2(new_n871), .B1(new_n848), .B2(new_n872), .ZN(G1338gat));
  NAND3_X1  g672(.A1(new_n791), .A2(new_n764), .A3(new_n837), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT118), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n791), .A2(new_n876), .A3(new_n764), .A4(new_n837), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(G106gat), .A3(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n729), .A2(G106gat), .A3(new_n331), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n847), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n874), .A2(G106gat), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n864), .A2(new_n865), .A3(new_n879), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT53), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(G1339gat));
  INV_X1    g684(.A(new_n782), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n240), .B1(new_n239), .B2(new_n241), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n230), .B1(new_n229), .B2(new_n233), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n250), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n254), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n722), .A2(new_n726), .A3(new_n891), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n715), .A2(new_n702), .A3(new_n716), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n894));
  OR3_X1    g693(.A1(new_n893), .A2(new_n717), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n700), .B1(new_n717), .B2(new_n894), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(KEYINPUT55), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT55), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n893), .A2(new_n717), .A3(new_n894), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n717), .A2(new_n894), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n720), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n897), .A2(new_n902), .A3(new_n255), .A4(new_n724), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n886), .B1(new_n892), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n897), .A2(new_n724), .ZN(new_n905));
  AOI21_X1  g704(.A(KEYINPUT55), .B1(new_n895), .B2(new_n896), .ZN(new_n906));
  NOR4_X1   g705(.A1(new_n905), .A2(new_n782), .A3(new_n906), .A4(new_n890), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n842), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n729), .A2(new_n696), .A3(new_n256), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n627), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n910), .A2(new_n487), .A3(new_n623), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n351), .A3(new_n255), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n764), .B1(new_n908), .B2(new_n909), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n627), .A2(new_n602), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n828), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G113gat), .B1(new_n915), .B2(new_n256), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT119), .Z(G1340gat));
  AOI21_X1  g717(.A(G120gat), .B1(new_n911), .B2(new_n728), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n915), .A2(new_n349), .A3(new_n729), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT120), .ZN(G1341gat));
  NAND3_X1  g721(.A1(new_n911), .A2(new_n344), .A3(new_n753), .ZN(new_n923));
  OAI21_X1  g722(.A(G127gat), .B1(new_n915), .B2(new_n842), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1342gat));
  NAND3_X1  g724(.A1(new_n911), .A2(new_n342), .A3(new_n656), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n926), .A2(KEYINPUT56), .ZN(new_n927));
  OAI21_X1  g726(.A(G134gat), .B1(new_n915), .B2(new_n655), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(KEYINPUT56), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(G1343gat));
  NOR2_X1   g729(.A1(new_n743), .A2(new_n331), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n910), .A2(new_n487), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n275), .B1(new_n932), .B2(new_n256), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n908), .A2(new_n909), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT57), .B1(new_n934), .B2(new_n764), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT57), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n656), .B1(new_n892), .B2(new_n903), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n842), .B1(new_n937), .B2(new_n907), .ZN(new_n938));
  AOI211_X1 g737(.A(new_n936), .B(new_n331), .C1(new_n938), .C2(new_n909), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n744), .B(new_n914), .C1(new_n935), .C2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n255), .A2(G141gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n933), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT121), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g743(.A(KEYINPUT59), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n945), .B(G148gat), .C1(new_n940), .C2(new_n729), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n744), .A2(new_n728), .A3(new_n914), .ZN(new_n948));
  NOR4_X1   g747(.A1(new_n905), .A2(new_n906), .A3(new_n655), .A4(new_n890), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n842), .B1(new_n937), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n331), .B1(new_n950), .B2(new_n909), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT122), .B1(new_n951), .B2(KEYINPUT57), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n934), .A2(KEYINPUT57), .A3(new_n764), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n951), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n948), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G148gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n947), .B1(new_n957), .B2(KEYINPUT59), .ZN(new_n958));
  AOI211_X1 g757(.A(KEYINPUT123), .B(new_n945), .C1(new_n956), .C2(G148gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n946), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n932), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n279), .A3(new_n728), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1345gat));
  OAI21_X1  g762(.A(G155gat), .B1(new_n940), .B2(new_n842), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n961), .A2(new_n297), .A3(new_n753), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1346gat));
  OR3_X1    g765(.A1(new_n940), .A2(new_n298), .A3(new_n782), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n298), .B1(new_n932), .B2(new_n655), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n967), .A2(new_n968), .ZN(G1347gat));
  AOI21_X1  g768(.A(new_n820), .B1(new_n908), .B2(new_n909), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(new_n602), .A3(new_n623), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n971), .A2(new_n409), .A3(new_n255), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n820), .A2(new_n487), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n913), .A2(new_n828), .A3(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT124), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n976), .A2(new_n255), .A3(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT125), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n978), .A2(new_n979), .A3(G169gat), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n978), .B2(G169gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n972), .B1(new_n980), .B2(new_n981), .ZN(G1348gat));
  NAND3_X1  g781(.A1(new_n971), .A2(new_n410), .A3(new_n728), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n976), .A2(new_n728), .A3(new_n977), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n984), .B2(new_n410), .ZN(G1349gat));
  NAND3_X1  g784(.A1(new_n976), .A2(new_n753), .A3(new_n977), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n753), .A2(new_n401), .A3(new_n403), .ZN(new_n987));
  AOI22_X1  g786(.A1(new_n986), .A2(G183gat), .B1(new_n971), .B2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n988), .A2(new_n989), .A3(KEYINPUT60), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n989), .A2(KEYINPUT60), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n989), .A2(KEYINPUT60), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n990), .A2(new_n993), .ZN(G1350gat));
  NAND4_X1  g793(.A1(new_n971), .A2(new_n397), .A3(new_n399), .A4(new_n886), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n976), .A2(new_n656), .A3(new_n977), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n996), .A2(new_n997), .A3(G190gat), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n997), .B1(new_n996), .B2(G190gat), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(G1351gat));
  AND3_X1   g799(.A1(new_n970), .A2(new_n602), .A3(new_n931), .ZN(new_n1001));
  AOI21_X1  g800(.A(G197gat), .B1(new_n1001), .B2(new_n255), .ZN(new_n1002));
  NOR3_X1   g801(.A1(new_n743), .A2(new_n820), .A3(new_n487), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1003), .B1(new_n954), .B2(new_n955), .ZN(new_n1004));
  INV_X1    g803(.A(new_n1004), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n255), .A2(G197gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(G1352gat));
  INV_X1    g806(.A(G204gat), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1001), .A2(new_n1008), .A3(new_n728), .ZN(new_n1009));
  XOR2_X1   g808(.A(new_n1009), .B(KEYINPUT62), .Z(new_n1010));
  OAI21_X1  g809(.A(G204gat), .B1(new_n1004), .B2(new_n729), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1010), .A2(new_n1011), .ZN(G1353gat));
  OAI21_X1  g811(.A(G211gat), .B1(new_n1004), .B2(new_n842), .ZN(new_n1013));
  OR2_X1    g812(.A1(new_n1013), .A2(KEYINPUT63), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(KEYINPUT63), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1001), .A2(new_n264), .A3(new_n753), .ZN(new_n1016));
  XOR2_X1   g815(.A(new_n1016), .B(KEYINPUT127), .Z(new_n1017));
  NAND3_X1  g816(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(G1354gat));
  AOI21_X1  g817(.A(G218gat), .B1(new_n1001), .B2(new_n886), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n655), .A2(new_n263), .ZN(new_n1020));
  AOI21_X1  g819(.A(new_n1019), .B1(new_n1005), .B2(new_n1020), .ZN(G1355gat));
endmodule


