

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U559 ( .A1(n742), .A2(n741), .ZN(n743) );
  BUF_X4 U560 ( .A(n892), .Z(n523) );
  XNOR2_X1 U561 ( .A(n526), .B(KEYINPUT65), .ZN(n892) );
  XNOR2_X1 U562 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n529) );
  NOR2_X1 U563 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U564 ( .A1(n524), .A2(n819), .ZN(n820) );
  NAND2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  AND2_X1 U566 ( .A1(n830), .A2(n818), .ZN(n524) );
  XNOR2_X2 U567 ( .A(n529), .B(n528), .ZN(n896) );
  INV_X1 U568 ( .A(KEYINPUT27), .ZN(n692) );
  XNOR2_X1 U569 ( .A(n693), .B(n692), .ZN(n694) );
  INV_X1 U570 ( .A(KEYINPUT100), .ZN(n696) );
  INV_X1 U571 ( .A(KEYINPUT29), .ZN(n722) );
  INV_X1 U572 ( .A(KEYINPUT12), .ZN(n564) );
  XNOR2_X1 U573 ( .A(n564), .B(KEYINPUT77), .ZN(n565) );
  XNOR2_X1 U574 ( .A(n566), .B(n565), .ZN(n568) );
  NOR2_X1 U575 ( .A1(G651), .A2(G543), .ZN(n659) );
  NOR2_X1 U576 ( .A1(G2104), .A2(n536), .ZN(n893) );
  XNOR2_X1 U577 ( .A(KEYINPUT68), .B(n532), .ZN(n533) );
  XOR2_X1 U578 ( .A(KEYINPUT79), .B(n577), .Z(n961) );
  INV_X1 U579 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U580 ( .A1(G125), .A2(n893), .ZN(n525) );
  XNOR2_X1 U581 ( .A(n525), .B(KEYINPUT64), .ZN(n535) );
  NAND2_X1 U582 ( .A1(n523), .A2(G113), .ZN(n527) );
  XNOR2_X1 U583 ( .A(n527), .B(KEYINPUT66), .ZN(n531) );
  NOR2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  NAND2_X1 U585 ( .A1(G137), .A2(n896), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U587 ( .A(n533), .ZN(n534) );
  NAND2_X1 U588 ( .A1(n535), .A2(n534), .ZN(n539) );
  AND2_X1 U589 ( .A1(n536), .A2(G2104), .ZN(n897) );
  NAND2_X1 U590 ( .A1(G101), .A2(n897), .ZN(n537) );
  XNOR2_X1 U591 ( .A(KEYINPUT23), .B(n537), .ZN(n538) );
  NOR2_X2 U592 ( .A1(n539), .A2(n538), .ZN(G160) );
  AND2_X1 U593 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U594 ( .A(G57), .ZN(G237) );
  INV_X1 U595 ( .A(G132), .ZN(G219) );
  NAND2_X1 U596 ( .A1(G138), .A2(n896), .ZN(n541) );
  NAND2_X1 U597 ( .A1(G102), .A2(n897), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U599 ( .A(KEYINPUT92), .B(n542), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G114), .A2(n523), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G126), .A2(n893), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n546), .A2(n545), .ZN(G164) );
  NAND2_X1 U604 ( .A1(G89), .A2(n659), .ZN(n547) );
  XNOR2_X1 U605 ( .A(n547), .B(KEYINPUT84), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n548), .B(KEYINPUT4), .ZN(n550) );
  XOR2_X1 U607 ( .A(G543), .B(KEYINPUT0), .Z(n644) );
  INV_X1 U608 ( .A(G651), .ZN(n552) );
  NOR2_X1 U609 ( .A1(n644), .A2(n552), .ZN(n660) );
  NAND2_X1 U610 ( .A1(G76), .A2(n660), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U612 ( .A(n551), .B(KEYINPUT5), .ZN(n560) );
  NOR2_X1 U613 ( .A1(G543), .A2(n552), .ZN(n554) );
  XNOR2_X1 U614 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n553) );
  XNOR2_X1 U615 ( .A(n554), .B(n553), .ZN(n655) );
  NAND2_X1 U616 ( .A1(n655), .A2(G63), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT85), .B(n555), .Z(n557) );
  NOR2_X2 U618 ( .A1(G651), .A2(n644), .ZN(n654) );
  NAND2_X1 U619 ( .A1(n654), .A2(G51), .ZN(n556) );
  NAND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT6), .B(n558), .Z(n559) );
  NAND2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U623 ( .A(n561), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U627 ( .A(G223), .ZN(n839) );
  NAND2_X1 U628 ( .A1(n839), .A2(G567), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U630 ( .A1(G81), .A2(n659), .ZN(n566) );
  NAND2_X1 U631 ( .A1(G68), .A2(n660), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT13), .B(n569), .ZN(n576) );
  XOR2_X1 U634 ( .A(KEYINPUT76), .B(KEYINPUT14), .Z(n571) );
  NAND2_X1 U635 ( .A1(G56), .A2(n655), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G43), .A2(n654), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT78), .B(n572), .Z(n573) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  INV_X1 U641 ( .A(G860), .ZN(n626) );
  NOR2_X1 U642 ( .A1(n961), .A2(n626), .ZN(n578) );
  XOR2_X1 U643 ( .A(KEYINPUT80), .B(n578), .Z(G153) );
  NAND2_X1 U644 ( .A1(G52), .A2(n654), .ZN(n587) );
  NAND2_X1 U645 ( .A1(n655), .A2(G64), .ZN(n579) );
  XNOR2_X1 U646 ( .A(KEYINPUT71), .B(n579), .ZN(n585) );
  NAND2_X1 U647 ( .A1(G90), .A2(n659), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G77), .A2(n660), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U650 ( .A(KEYINPUT9), .B(n582), .Z(n583) );
  XNOR2_X1 U651 ( .A(KEYINPUT72), .B(n583), .ZN(n584) );
  NOR2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n588), .B(KEYINPUT73), .ZN(G171) );
  XNOR2_X1 U655 ( .A(G171), .B(KEYINPUT81), .ZN(G301) );
  NAND2_X1 U656 ( .A1(G868), .A2(G301), .ZN(n589) );
  XNOR2_X1 U657 ( .A(n589), .B(KEYINPUT82), .ZN(n599) );
  INV_X1 U658 ( .A(G868), .ZN(n612) );
  NAND2_X1 U659 ( .A1(G79), .A2(n660), .ZN(n596) );
  NAND2_X1 U660 ( .A1(G66), .A2(n655), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G92), .A2(n659), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G54), .A2(n654), .ZN(n592) );
  XNOR2_X1 U664 ( .A(KEYINPUT83), .B(n592), .ZN(n593) );
  NOR2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n597), .B(KEYINPUT15), .ZN(n960) );
  INV_X1 U668 ( .A(n960), .ZN(n710) );
  NAND2_X1 U669 ( .A1(n612), .A2(n710), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U671 ( .A1(G91), .A2(n659), .ZN(n601) );
  NAND2_X1 U672 ( .A1(G78), .A2(n660), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n655), .A2(G65), .ZN(n602) );
  XOR2_X1 U675 ( .A(KEYINPUT74), .B(n602), .Z(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n654), .A2(G53), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(G299) );
  NOR2_X1 U679 ( .A1(G286), .A2(n612), .ZN(n608) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n626), .A2(G559), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n609), .A2(n960), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  OR2_X1 U685 ( .A1(G559), .A2(n710), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n611), .A2(G868), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n961), .A2(n612), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U689 ( .A1(G135), .A2(n896), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G111), .A2(n523), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n893), .A2(G123), .ZN(n617) );
  XOR2_X1 U693 ( .A(KEYINPUT18), .B(n617), .Z(n618) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n897), .A2(G99), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n937) );
  XOR2_X1 U697 ( .A(G2096), .B(KEYINPUT86), .Z(n622) );
  XNOR2_X1 U698 ( .A(n937), .B(n622), .ZN(n624) );
  INV_X1 U699 ( .A(G2100), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(G156) );
  NAND2_X1 U701 ( .A1(G559), .A2(n960), .ZN(n625) );
  XOR2_X1 U702 ( .A(n961), .B(n625), .Z(n670) );
  NAND2_X1 U703 ( .A1(n626), .A2(n670), .ZN(n633) );
  NAND2_X1 U704 ( .A1(G93), .A2(n659), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G80), .A2(n660), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U707 ( .A1(G67), .A2(n655), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G55), .A2(n654), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n674) );
  XOR2_X1 U711 ( .A(n633), .B(n674), .Z(G145) );
  NAND2_X1 U712 ( .A1(G61), .A2(n655), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G86), .A2(n659), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n660), .A2(G73), .ZN(n636) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n654), .A2(G48), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U720 ( .A1(G49), .A2(n654), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U723 ( .A1(n655), .A2(n643), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n644), .A2(G87), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(G288) );
  NAND2_X1 U726 ( .A1(G88), .A2(n659), .ZN(n648) );
  NAND2_X1 U727 ( .A1(G75), .A2(n660), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G62), .A2(n655), .ZN(n649) );
  XNOR2_X1 U730 ( .A(KEYINPUT87), .B(n649), .ZN(n650) );
  NOR2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n654), .A2(G50), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(G303) );
  INV_X1 U734 ( .A(G303), .ZN(G166) );
  NAND2_X1 U735 ( .A1(n654), .A2(G47), .ZN(n657) );
  NAND2_X1 U736 ( .A1(n655), .A2(G60), .ZN(n656) );
  NAND2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U738 ( .A(KEYINPUT70), .B(n658), .Z(n664) );
  NAND2_X1 U739 ( .A1(G85), .A2(n659), .ZN(n662) );
  NAND2_X1 U740 ( .A1(G72), .A2(n660), .ZN(n661) );
  AND2_X1 U741 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U742 ( .A1(n664), .A2(n663), .ZN(G290) );
  XNOR2_X1 U743 ( .A(G288), .B(KEYINPUT19), .ZN(n666) );
  INV_X1 U744 ( .A(G299), .ZN(n717) );
  XNOR2_X1 U745 ( .A(n717), .B(G166), .ZN(n665) );
  XNOR2_X1 U746 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U747 ( .A(n674), .B(n667), .Z(n668) );
  XNOR2_X1 U748 ( .A(G305), .B(n668), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n669), .B(G290), .ZN(n907) );
  XNOR2_X1 U750 ( .A(n907), .B(n670), .ZN(n671) );
  XNOR2_X1 U751 ( .A(n671), .B(KEYINPUT88), .ZN(n672) );
  NAND2_X1 U752 ( .A1(n672), .A2(G868), .ZN(n673) );
  XOR2_X1 U753 ( .A(KEYINPUT89), .B(n673), .Z(n676) );
  OR2_X1 U754 ( .A1(n674), .A2(G868), .ZN(n675) );
  NAND2_X1 U755 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U757 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n678), .ZN(n680) );
  XNOR2_X1 U759 ( .A(KEYINPUT90), .B(KEYINPUT21), .ZN(n679) );
  XNOR2_X1 U760 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U761 ( .A1(G2072), .A2(n681), .ZN(G158) );
  XNOR2_X1 U762 ( .A(KEYINPUT75), .B(G82), .ZN(G220) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U764 ( .A1(G219), .A2(G220), .ZN(n682) );
  XNOR2_X1 U765 ( .A(KEYINPUT22), .B(n682), .ZN(n683) );
  NAND2_X1 U766 ( .A1(n683), .A2(G96), .ZN(n684) );
  NOR2_X1 U767 ( .A1(n684), .A2(G218), .ZN(n685) );
  XNOR2_X1 U768 ( .A(n685), .B(KEYINPUT91), .ZN(n845) );
  NAND2_X1 U769 ( .A1(n845), .A2(G2106), .ZN(n689) );
  NAND2_X1 U770 ( .A1(G120), .A2(G69), .ZN(n686) );
  NOR2_X1 U771 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U772 ( .A1(G108), .A2(n687), .ZN(n846) );
  NAND2_X1 U773 ( .A1(n846), .A2(G567), .ZN(n688) );
  NAND2_X1 U774 ( .A1(n689), .A2(n688), .ZN(n847) );
  NAND2_X1 U775 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U776 ( .A1(n847), .A2(n690), .ZN(n844) );
  NAND2_X1 U777 ( .A1(n844), .A2(G36), .ZN(G176) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n786) );
  INV_X1 U779 ( .A(n786), .ZN(n691) );
  NOR2_X1 U780 ( .A1(G164), .A2(G1384), .ZN(n787) );
  NAND2_X1 U781 ( .A1(n691), .A2(n787), .ZN(n702) );
  BUF_X2 U782 ( .A(n702), .Z(n732) );
  NAND2_X1 U783 ( .A1(G1956), .A2(n732), .ZN(n695) );
  INV_X1 U784 ( .A(n702), .ZN(n724) );
  NAND2_X1 U785 ( .A1(n724), .A2(G2072), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n697) );
  XNOR2_X1 U787 ( .A(n697), .B(n696), .ZN(n716) );
  NOR2_X1 U788 ( .A1(n717), .A2(n716), .ZN(n699) );
  XNOR2_X1 U789 ( .A(KEYINPUT101), .B(KEYINPUT28), .ZN(n698) );
  XNOR2_X1 U790 ( .A(n699), .B(n698), .ZN(n721) );
  NOR2_X1 U791 ( .A1(n724), .A2(G1348), .ZN(n701) );
  NOR2_X1 U792 ( .A1(G2067), .A2(n732), .ZN(n700) );
  NOR2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n711) );
  NAND2_X1 U794 ( .A1(n710), .A2(n711), .ZN(n709) );
  INV_X1 U795 ( .A(G1996), .ZN(n1015) );
  NOR2_X1 U796 ( .A1(n702), .A2(n1015), .ZN(n704) );
  INV_X1 U797 ( .A(KEYINPUT26), .ZN(n703) );
  XNOR2_X1 U798 ( .A(n704), .B(n703), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n732), .A2(G1341), .ZN(n705) );
  NAND2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U801 ( .A1(n961), .A2(n707), .ZN(n708) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n713) );
  OR2_X1 U803 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n715) );
  INV_X1 U805 ( .A(KEYINPUT102), .ZN(n714) );
  XNOR2_X1 U806 ( .A(n715), .B(n714), .ZN(n719) );
  NAND2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U809 ( .A1(n721), .A2(n720), .ZN(n723) );
  XNOR2_X1 U810 ( .A(n723), .B(n722), .ZN(n730) );
  NOR2_X1 U811 ( .A1(n724), .A2(G1961), .ZN(n725) );
  XOR2_X1 U812 ( .A(KEYINPUT98), .B(n725), .Z(n728) );
  XOR2_X1 U813 ( .A(G2078), .B(KEYINPUT25), .Z(n1018) );
  NOR2_X1 U814 ( .A1(n1018), .A2(n732), .ZN(n726) );
  XNOR2_X1 U815 ( .A(KEYINPUT99), .B(n726), .ZN(n727) );
  NAND2_X1 U816 ( .A1(n728), .A2(n727), .ZN(n737) );
  NAND2_X1 U817 ( .A1(G171), .A2(n737), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U819 ( .A(KEYINPUT103), .B(n731), .ZN(n742) );
  NAND2_X1 U820 ( .A1(G8), .A2(n732), .ZN(n781) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n781), .ZN(n755) );
  NOR2_X1 U822 ( .A1(G2084), .A2(n732), .ZN(n756) );
  NOR2_X1 U823 ( .A1(n755), .A2(n756), .ZN(n733) );
  XNOR2_X1 U824 ( .A(KEYINPUT104), .B(n733), .ZN(n734) );
  NAND2_X1 U825 ( .A1(n734), .A2(G8), .ZN(n735) );
  XNOR2_X1 U826 ( .A(KEYINPUT30), .B(n735), .ZN(n736) );
  NOR2_X1 U827 ( .A1(G168), .A2(n736), .ZN(n739) );
  NOR2_X1 U828 ( .A1(G171), .A2(n737), .ZN(n738) );
  NOR2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U830 ( .A(n740), .B(KEYINPUT31), .ZN(n741) );
  XNOR2_X1 U831 ( .A(n743), .B(KEYINPUT105), .ZN(n753) );
  NAND2_X1 U832 ( .A1(n753), .A2(G286), .ZN(n750) );
  INV_X1 U833 ( .A(G8), .ZN(n748) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n781), .ZN(n745) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n732), .ZN(n744) );
  NOR2_X1 U836 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U837 ( .A1(n746), .A2(G303), .ZN(n747) );
  OR2_X1 U838 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n752) );
  INV_X1 U840 ( .A(KEYINPUT32), .ZN(n751) );
  XNOR2_X1 U841 ( .A(n752), .B(n751), .ZN(n773) );
  INV_X1 U842 ( .A(n773), .ZN(n760) );
  INV_X1 U843 ( .A(n753), .ZN(n754) );
  NOR2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n758) );
  NAND2_X1 U845 ( .A1(G8), .A2(n756), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n774) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n965) );
  NAND2_X1 U848 ( .A1(n774), .A2(n965), .ZN(n759) );
  NOR2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n767) );
  INV_X1 U850 ( .A(n965), .ZN(n762) );
  NOR2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n768) );
  NOR2_X1 U852 ( .A1(G1971), .A2(G303), .ZN(n761) );
  NOR2_X1 U853 ( .A1(n768), .A2(n761), .ZN(n969) );
  OR2_X1 U854 ( .A1(n762), .A2(n969), .ZN(n763) );
  OR2_X1 U855 ( .A1(n781), .A2(n763), .ZN(n765) );
  INV_X1 U856 ( .A(KEYINPUT33), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n771) );
  NAND2_X1 U859 ( .A1(n768), .A2(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U860 ( .A1(n769), .A2(n781), .ZN(n770) );
  NOR2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U862 ( .A(G1981), .B(G305), .Z(n957) );
  AND2_X1 U863 ( .A1(n772), .A2(n957), .ZN(n785) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n777) );
  NOR2_X1 U865 ( .A1(G2090), .A2(G303), .ZN(n775) );
  NAND2_X1 U866 ( .A1(G8), .A2(n775), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U868 ( .A1(n778), .A2(n781), .ZN(n783) );
  NOR2_X1 U869 ( .A1(G1981), .A2(G305), .ZN(n779) );
  XOR2_X1 U870 ( .A(n779), .B(KEYINPUT24), .Z(n780) );
  OR2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n821) );
  NOR2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n834) );
  NAND2_X1 U875 ( .A1(G140), .A2(n896), .ZN(n789) );
  NAND2_X1 U876 ( .A1(G104), .A2(n897), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n791) );
  XOR2_X1 U878 ( .A(KEYINPUT93), .B(KEYINPUT34), .Z(n790) );
  XNOR2_X1 U879 ( .A(n791), .B(n790), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G116), .A2(n523), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G128), .A2(n893), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U883 ( .A(KEYINPUT35), .B(n794), .Z(n795) );
  NOR2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U885 ( .A(n797), .B(KEYINPUT36), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n798), .B(KEYINPUT94), .ZN(n889) );
  XNOR2_X1 U887 ( .A(KEYINPUT37), .B(G2067), .ZN(n832) );
  NOR2_X1 U888 ( .A1(n889), .A2(n832), .ZN(n945) );
  NAND2_X1 U889 ( .A1(n834), .A2(n945), .ZN(n830) );
  NAND2_X1 U890 ( .A1(G107), .A2(n523), .ZN(n800) );
  NAND2_X1 U891 ( .A1(G119), .A2(n893), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U893 ( .A(n801), .B(KEYINPUT95), .ZN(n806) );
  NAND2_X1 U894 ( .A1(G131), .A2(n896), .ZN(n803) );
  NAND2_X1 U895 ( .A1(G95), .A2(n897), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n804) );
  XOR2_X1 U897 ( .A(KEYINPUT96), .B(n804), .Z(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U899 ( .A(n807), .B(KEYINPUT97), .Z(n888) );
  AND2_X1 U900 ( .A1(n888), .A2(G1991), .ZN(n816) );
  NAND2_X1 U901 ( .A1(G141), .A2(n896), .ZN(n809) );
  NAND2_X1 U902 ( .A1(G117), .A2(n523), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n897), .A2(G105), .ZN(n810) );
  XOR2_X1 U905 ( .A(KEYINPUT38), .B(n810), .Z(n811) );
  NOR2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n893), .A2(G129), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n882) );
  AND2_X1 U909 ( .A1(G1996), .A2(n882), .ZN(n815) );
  NOR2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n947) );
  INV_X1 U911 ( .A(n834), .ZN(n817) );
  NOR2_X1 U912 ( .A1(n947), .A2(n817), .ZN(n826) );
  INV_X1 U913 ( .A(n826), .ZN(n818) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n971) );
  NAND2_X1 U915 ( .A1(n971), .A2(n834), .ZN(n819) );
  INV_X1 U916 ( .A(n822), .ZN(n837) );
  XOR2_X1 U917 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n823) );
  XNOR2_X1 U918 ( .A(KEYINPUT106), .B(n823), .ZN(n829) );
  NOR2_X1 U919 ( .A1(G1996), .A2(n882), .ZN(n935) );
  NOR2_X1 U920 ( .A1(G1991), .A2(n888), .ZN(n940) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n824) );
  NOR2_X1 U922 ( .A1(n940), .A2(n824), .ZN(n825) );
  NOR2_X1 U923 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U924 ( .A1(n935), .A2(n827), .ZN(n828) );
  XNOR2_X1 U925 ( .A(n829), .B(n828), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n889), .A2(n832), .ZN(n949) );
  NAND2_X1 U928 ( .A1(n833), .A2(n949), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U931 ( .A(KEYINPUT40), .B(n838), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n839), .ZN(G217) );
  NAND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n841) );
  INV_X1 U934 ( .A(G661), .ZN(n840) );
  NOR2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U936 ( .A(n842), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U938 ( .A1(n844), .A2(n843), .ZN(G188) );
  XOR2_X1 U939 ( .A(G96), .B(KEYINPUT110), .Z(G221) );
  XNOR2_X1 U940 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  NOR2_X1 U943 ( .A1(n846), .A2(n845), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  INV_X1 U945 ( .A(n847), .ZN(G319) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n849) );
  XNOR2_X1 U947 ( .A(G2072), .B(G2678), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U949 ( .A(n850), .B(KEYINPUT112), .Z(n852) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2090), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U952 ( .A(KEYINPUT42), .B(G2100), .Z(n854) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(G227) );
  XOR2_X1 U956 ( .A(G1976), .B(G1961), .Z(n858) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1966), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U959 ( .A(G1971), .B(G1956), .Z(n860) );
  XNOR2_X1 U960 ( .A(G1996), .B(G1991), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U962 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U963 ( .A(G2474), .B(KEYINPUT113), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n866) );
  XOR2_X1 U965 ( .A(G1981), .B(KEYINPUT41), .Z(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(G229) );
  NAND2_X1 U967 ( .A1(G124), .A2(n893), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n523), .A2(G112), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G136), .A2(n896), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G100), .A2(n897), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U974 ( .A1(n873), .A2(n872), .ZN(G162) );
  XOR2_X1 U975 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n884) );
  NAND2_X1 U976 ( .A1(G115), .A2(n523), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G127), .A2(n893), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n876), .B(KEYINPUT47), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G139), .A2(n896), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n881) );
  NAND2_X1 U982 ( .A1(n897), .A2(G103), .ZN(n879) );
  XOR2_X1 U983 ( .A(KEYINPUT114), .B(n879), .Z(n880) );
  NOR2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n929) );
  XOR2_X1 U985 ( .A(n882), .B(n929), .Z(n883) );
  XNOR2_X1 U986 ( .A(n884), .B(n883), .ZN(n887) );
  XOR2_X1 U987 ( .A(G164), .B(G162), .Z(n885) );
  XNOR2_X1 U988 ( .A(n937), .B(n885), .ZN(n886) );
  XOR2_X1 U989 ( .A(n887), .B(n886), .Z(n891) );
  XOR2_X1 U990 ( .A(n889), .B(n888), .Z(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n905) );
  NAND2_X1 U992 ( .A1(G118), .A2(n523), .ZN(n895) );
  NAND2_X1 U993 ( .A1(G130), .A2(n893), .ZN(n894) );
  NAND2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n902) );
  NAND2_X1 U995 ( .A1(G142), .A2(n896), .ZN(n899) );
  NAND2_X1 U996 ( .A1(G106), .A2(n897), .ZN(n898) );
  NAND2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(KEYINPUT45), .B(n900), .Z(n901) );
  NOR2_X1 U999 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(G160), .B(n903), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n906), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(n961), .B(n907), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(G171), .B(n960), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(G286), .B(n910), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n911), .ZN(G397) );
  XOR2_X1 U1008 ( .A(KEYINPUT108), .B(G2446), .Z(n913) );
  XNOR2_X1 U1009 ( .A(G2443), .B(G2454), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1011 ( .A(n914), .B(G2451), .Z(n916) );
  XNOR2_X1 U1012 ( .A(G1348), .B(G1341), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(n916), .B(n915), .ZN(n920) );
  XOR2_X1 U1014 ( .A(G2435), .B(G2427), .Z(n918) );
  XNOR2_X1 U1015 ( .A(G2430), .B(G2438), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1017 ( .A(n920), .B(n919), .Z(n921) );
  NAND2_X1 U1018 ( .A1(G14), .A2(n921), .ZN(n928) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n928), .ZN(n925) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n922) );
  XOR2_X1 U1021 ( .A(KEYINPUT49), .B(n922), .Z(n923) );
  XNOR2_X1 U1022 ( .A(n923), .B(KEYINPUT115), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G108), .ZN(G238) );
  INV_X1 U1028 ( .A(n928), .ZN(G401) );
  XNOR2_X1 U1029 ( .A(G164), .B(G2078), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G2072), .B(n929), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(n930), .B(KEYINPUT118), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(n933), .B(KEYINPUT50), .ZN(n952) );
  XOR2_X1 U1034 ( .A(G2090), .B(G162), .Z(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1036 ( .A(KEYINPUT51), .B(n936), .Z(n943) );
  XNOR2_X1 U1037 ( .A(G160), .B(G2084), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(n941), .B(KEYINPUT116), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(n948), .B(KEYINPUT117), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(n953), .ZN(n955) );
  INV_X1 U1048 ( .A(KEYINPUT55), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n956), .A2(G29), .ZN(n1035) );
  XNOR2_X1 U1051 ( .A(G16), .B(KEYINPUT56), .ZN(n980) );
  XNOR2_X1 U1052 ( .A(G1966), .B(G168), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(n959), .B(KEYINPUT57), .ZN(n978) );
  XOR2_X1 U1055 ( .A(G1348), .B(n960), .Z(n963) );
  XNOR2_X1 U1056 ( .A(n961), .B(G1341), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n974) );
  NAND2_X1 U1058 ( .A1(G1971), .A2(G303), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G1956), .B(G299), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1064 ( .A(KEYINPUT121), .B(n972), .Z(n973) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n976) );
  XOR2_X1 U1066 ( .A(G171), .B(G1961), .Z(n975) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n1008) );
  INV_X1 U1070 ( .A(G16), .ZN(n1006) );
  XNOR2_X1 U1071 ( .A(G1348), .B(KEYINPUT59), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(n981), .B(G4), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(G1956), .B(G20), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(G19), .B(G1341), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1077 ( .A(KEYINPUT123), .B(G1981), .Z(n986) );
  XNOR2_X1 U1078 ( .A(G6), .B(n986), .ZN(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(KEYINPUT124), .B(n989), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n990), .B(KEYINPUT60), .ZN(n1000) );
  XNOR2_X1 U1082 ( .A(G1961), .B(KEYINPUT122), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n991), .B(G5), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(G1971), .B(G22), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(G23), .B(G1976), .ZN(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n995) );
  XOR2_X1 U1087 ( .A(G1986), .B(G24), .Z(n994) );
  NAND2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(KEYINPUT58), .B(n996), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(KEYINPUT125), .B(G1966), .Z(n1001) );
  XNOR2_X1 U1093 ( .A(G21), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(KEYINPUT61), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1098 ( .A(KEYINPUT126), .B(n1009), .Z(n1010) );
  NAND2_X1 U1099 ( .A1(G11), .A2(n1010), .ZN(n1033) );
  XOR2_X1 U1100 ( .A(G2072), .B(G33), .Z(n1011) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(G28), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(G25), .B(G1991), .Z(n1012) );
  XNOR2_X1 U1103 ( .A(KEYINPUT119), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1022) );
  XOR2_X1 U1105 ( .A(G2067), .B(G26), .Z(n1017) );
  XNOR2_X1 U1106 ( .A(n1015), .B(G32), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(G27), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(n1023), .B(KEYINPUT53), .ZN(n1026) );
  XOR2_X1 U1112 ( .A(G2084), .B(G34), .Z(n1024) );
  XNOR2_X1 U1113 ( .A(KEYINPUT54), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(G35), .B(G2090), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1117 ( .A(KEYINPUT55), .B(n1029), .Z(n1030) );
  NOR2_X1 U1118 ( .A1(G29), .A2(n1030), .ZN(n1031) );
  XNOR2_X1 U1119 ( .A(n1031), .B(KEYINPUT120), .ZN(n1032) );
  NOR2_X1 U1120 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1122 ( .A(n1036), .B(KEYINPUT127), .ZN(n1037) );
  XNOR2_X1 U1123 ( .A(KEYINPUT62), .B(n1037), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

