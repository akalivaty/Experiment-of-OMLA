

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U547 ( .A1(G8), .A2(n655), .ZN(n692) );
  BUF_X1 U548 ( .A(n702), .Z(n703) );
  BUF_X2 U549 ( .A(n609), .Z(n655) );
  AND2_X1 U550 ( .A1(n734), .A2(n747), .ZN(n514) );
  OR2_X1 U551 ( .A1(n962), .A2(n626), .ZN(n625) );
  XNOR2_X1 U552 ( .A(n639), .B(KEYINPUT29), .ZN(n640) );
  NOR2_X1 U553 ( .A1(n653), .A2(n652), .ZN(n654) );
  OR2_X1 U554 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U555 ( .A1(G2105), .A2(G2104), .ZN(n515) );
  NAND2_X1 U556 ( .A1(G160), .A2(G40), .ZN(n720) );
  NOR2_X1 U557 ( .A1(n739), .A2(n514), .ZN(n735) );
  NOR2_X1 U558 ( .A1(G651), .A2(n578), .ZN(n783) );
  AND2_X1 U559 ( .A1(n537), .A2(n536), .ZN(G164) );
  XOR2_X1 U560 ( .A(KEYINPUT17), .B(n515), .Z(n516) );
  XNOR2_X1 U561 ( .A(n516), .B(KEYINPUT66), .ZN(n702) );
  NAND2_X1 U562 ( .A1(n702), .A2(G137), .ZN(n526) );
  AND2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n867) );
  NAND2_X1 U564 ( .A1(G113), .A2(n867), .ZN(n517) );
  XOR2_X1 U565 ( .A(KEYINPUT65), .B(n517), .Z(n524) );
  INV_X1 U566 ( .A(KEYINPUT23), .ZN(n519) );
  INV_X1 U567 ( .A(G2104), .ZN(n520) );
  NOR2_X4 U568 ( .A1(G2105), .A2(n520), .ZN(n864) );
  NAND2_X1 U569 ( .A1(G101), .A2(n864), .ZN(n518) );
  XNOR2_X1 U570 ( .A(n519), .B(n518), .ZN(n522) );
  AND2_X1 U571 ( .A1(n520), .A2(G2105), .ZN(n868) );
  NAND2_X1 U572 ( .A1(n868), .A2(G125), .ZN(n521) );
  AND2_X1 U573 ( .A1(n522), .A2(n521), .ZN(n523) );
  AND2_X1 U574 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n528) );
  INV_X1 U576 ( .A(KEYINPUT64), .ZN(n527) );
  XNOR2_X2 U577 ( .A(n528), .B(n527), .ZN(G160) );
  NAND2_X1 U578 ( .A1(n702), .A2(G138), .ZN(n529) );
  XNOR2_X1 U579 ( .A(n529), .B(KEYINPUT88), .ZN(n531) );
  NAND2_X1 U580 ( .A1(G102), .A2(n864), .ZN(n530) );
  NAND2_X1 U581 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U582 ( .A(n532), .B(KEYINPUT89), .ZN(n537) );
  NAND2_X1 U583 ( .A1(G126), .A2(n868), .ZN(n535) );
  NAND2_X1 U584 ( .A1(G114), .A2(n867), .ZN(n533) );
  XOR2_X1 U585 ( .A(KEYINPUT87), .B(n533), .Z(n534) );
  AND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U587 ( .A1(G651), .A2(G543), .ZN(n775) );
  NAND2_X1 U588 ( .A1(n775), .A2(G91), .ZN(n539) );
  XOR2_X1 U589 ( .A(KEYINPUT0), .B(G543), .Z(n578) );
  XNOR2_X1 U590 ( .A(KEYINPUT67), .B(G651), .ZN(n540) );
  NOR2_X1 U591 ( .A1(n578), .A2(n540), .ZN(n776) );
  NAND2_X1 U592 ( .A1(G78), .A2(n776), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n539), .A2(n538), .ZN(n546) );
  NOR2_X1 U594 ( .A1(G543), .A2(n540), .ZN(n542) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(KEYINPUT68), .Z(n541) );
  XNOR2_X1 U596 ( .A(n542), .B(n541), .ZN(n780) );
  NAND2_X1 U597 ( .A1(G65), .A2(n780), .ZN(n544) );
  NAND2_X1 U598 ( .A1(G53), .A2(n783), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U600 ( .A1(n546), .A2(n545), .ZN(G299) );
  NAND2_X1 U601 ( .A1(n775), .A2(G90), .ZN(n547) );
  XOR2_X1 U602 ( .A(KEYINPUT71), .B(n547), .Z(n549) );
  NAND2_X1 U603 ( .A1(G77), .A2(n776), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U605 ( .A(n550), .B(KEYINPUT9), .ZN(n552) );
  NAND2_X1 U606 ( .A1(G64), .A2(n780), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n783), .A2(G52), .ZN(n553) );
  XOR2_X1 U609 ( .A(KEYINPUT70), .B(n553), .Z(n554) );
  NOR2_X1 U610 ( .A1(n555), .A2(n554), .ZN(G171) );
  INV_X1 U611 ( .A(G171), .ZN(G301) );
  NAND2_X1 U612 ( .A1(G89), .A2(n775), .ZN(n556) );
  XOR2_X1 U613 ( .A(KEYINPUT4), .B(n556), .Z(n557) );
  XNOR2_X1 U614 ( .A(n557), .B(KEYINPUT77), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G76), .A2(n776), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U617 ( .A(n560), .B(KEYINPUT5), .ZN(n565) );
  NAND2_X1 U618 ( .A1(G63), .A2(n780), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G51), .A2(n783), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U621 ( .A(KEYINPUT6), .B(n563), .Z(n564) );
  NAND2_X1 U622 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U623 ( .A(n566), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U624 ( .A1(n775), .A2(G88), .ZN(n568) );
  NAND2_X1 U625 ( .A1(G75), .A2(n776), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U627 ( .A1(G62), .A2(n780), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G50), .A2(n783), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U630 ( .A1(n572), .A2(n571), .ZN(G166) );
  XOR2_X1 U631 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(n573) );
  XNOR2_X1 U633 ( .A(KEYINPUT78), .B(n573), .ZN(G286) );
  NAND2_X1 U634 ( .A1(G49), .A2(n783), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G74), .A2(G651), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT83), .B(n576), .Z(n577) );
  NOR2_X1 U638 ( .A1(n780), .A2(n577), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n578), .A2(G87), .ZN(n579) );
  NAND2_X1 U640 ( .A1(n580), .A2(n579), .ZN(G288) );
  XOR2_X1 U641 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n582) );
  NAND2_X1 U642 ( .A1(G73), .A2(n776), .ZN(n581) );
  XNOR2_X1 U643 ( .A(n582), .B(n581), .ZN(n586) );
  NAND2_X1 U644 ( .A1(G61), .A2(n780), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G86), .A2(n775), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U647 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U648 ( .A1(n783), .A2(G48), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n588), .A2(n587), .ZN(G305) );
  NAND2_X1 U650 ( .A1(n775), .A2(G85), .ZN(n590) );
  NAND2_X1 U651 ( .A1(G72), .A2(n776), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U653 ( .A1(G47), .A2(n783), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT69), .B(n591), .ZN(n592) );
  NOR2_X1 U655 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U656 ( .A1(n780), .A2(G60), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n595), .A2(n594), .ZN(G290) );
  NAND2_X1 U658 ( .A1(n783), .A2(G54), .ZN(n597) );
  NAND2_X1 U659 ( .A1(G79), .A2(n776), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n597), .A2(n596), .ZN(n602) );
  NAND2_X1 U661 ( .A1(G66), .A2(n780), .ZN(n599) );
  NAND2_X1 U662 ( .A1(G92), .A2(n775), .ZN(n598) );
  NAND2_X1 U663 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U664 ( .A(KEYINPUT75), .B(n600), .Z(n601) );
  NOR2_X1 U665 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U666 ( .A(KEYINPUT15), .B(n603), .Z(n962) );
  NOR2_X1 U667 ( .A1(G164), .A2(G1384), .ZN(n721) );
  INV_X1 U668 ( .A(KEYINPUT94), .ZN(n604) );
  XNOR2_X1 U669 ( .A(n604), .B(n720), .ZN(n605) );
  NAND2_X1 U670 ( .A1(n721), .A2(n605), .ZN(n609) );
  INV_X1 U671 ( .A(n609), .ZN(n642) );
  NAND2_X1 U672 ( .A1(n642), .A2(G2067), .ZN(n607) );
  NAND2_X1 U673 ( .A1(G1348), .A2(n609), .ZN(n606) );
  NAND2_X1 U674 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U675 ( .A(KEYINPUT95), .B(n608), .ZN(n626) );
  INV_X1 U676 ( .A(G1996), .ZN(n938) );
  NOR2_X1 U677 ( .A1(n655), .A2(n938), .ZN(n610) );
  XOR2_X1 U678 ( .A(n610), .B(KEYINPUT26), .Z(n623) );
  AND2_X1 U679 ( .A1(n655), .A2(G1341), .ZN(n621) );
  NAND2_X1 U680 ( .A1(n780), .A2(G56), .ZN(n611) );
  XOR2_X1 U681 ( .A(KEYINPUT14), .B(n611), .Z(n617) );
  NAND2_X1 U682 ( .A1(n775), .A2(G81), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n612), .B(KEYINPUT12), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G68), .A2(n776), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U686 ( .A(KEYINPUT13), .B(n615), .Z(n616) );
  NOR2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n618), .B(KEYINPUT74), .ZN(n620) );
  NAND2_X1 U689 ( .A1(G43), .A2(n783), .ZN(n619) );
  NAND2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n968) );
  NOR2_X1 U691 ( .A1(n621), .A2(n968), .ZN(n622) );
  AND2_X1 U692 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U694 ( .A1(n626), .A2(n962), .ZN(n627) );
  NAND2_X1 U695 ( .A1(n628), .A2(n627), .ZN(n633) );
  NAND2_X1 U696 ( .A1(n642), .A2(G2072), .ZN(n629) );
  XOR2_X1 U697 ( .A(KEYINPUT27), .B(n629), .Z(n631) );
  NAND2_X1 U698 ( .A1(G1956), .A2(n655), .ZN(n630) );
  NAND2_X1 U699 ( .A1(n631), .A2(n630), .ZN(n635) );
  NOR2_X1 U700 ( .A1(n635), .A2(G299), .ZN(n632) );
  NOR2_X1 U701 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n634), .B(KEYINPUT96), .ZN(n638) );
  NAND2_X1 U703 ( .A1(G299), .A2(n635), .ZN(n636) );
  XOR2_X1 U704 ( .A(n636), .B(KEYINPUT28), .Z(n637) );
  NOR2_X1 U705 ( .A1(n638), .A2(n637), .ZN(n641) );
  INV_X1 U706 ( .A(KEYINPUT97), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n641), .B(n640), .ZN(n646) );
  NAND2_X1 U708 ( .A1(G1961), .A2(n655), .ZN(n644) );
  XOR2_X1 U709 ( .A(G2078), .B(KEYINPUT25), .Z(n940) );
  NAND2_X1 U710 ( .A1(n642), .A2(n940), .ZN(n643) );
  NAND2_X1 U711 ( .A1(n644), .A2(n643), .ZN(n647) );
  OR2_X1 U712 ( .A1(n647), .A2(G301), .ZN(n645) );
  NAND2_X1 U713 ( .A1(n646), .A2(n645), .ZN(n668) );
  NAND2_X1 U714 ( .A1(G301), .A2(n647), .ZN(n648) );
  XOR2_X1 U715 ( .A(KEYINPUT98), .B(n648), .Z(n653) );
  NOR2_X1 U716 ( .A1(G1966), .A2(n692), .ZN(n670) );
  NOR2_X1 U717 ( .A1(G2084), .A2(n655), .ZN(n669) );
  NOR2_X1 U718 ( .A1(n670), .A2(n669), .ZN(n649) );
  NAND2_X1 U719 ( .A1(G8), .A2(n649), .ZN(n650) );
  XNOR2_X1 U720 ( .A(KEYINPUT30), .B(n650), .ZN(n651) );
  NOR2_X1 U721 ( .A1(G168), .A2(n651), .ZN(n652) );
  XOR2_X1 U722 ( .A(KEYINPUT31), .B(n654), .Z(n667) );
  NOR2_X1 U723 ( .A1(G1971), .A2(n692), .ZN(n657) );
  NOR2_X1 U724 ( .A1(G2090), .A2(n655), .ZN(n656) );
  NOR2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n658), .A2(G303), .ZN(n660) );
  AND2_X1 U727 ( .A1(n667), .A2(n660), .ZN(n659) );
  NAND2_X1 U728 ( .A1(n668), .A2(n659), .ZN(n664) );
  INV_X1 U729 ( .A(n660), .ZN(n661) );
  OR2_X1 U730 ( .A1(n661), .A2(G286), .ZN(n662) );
  AND2_X1 U731 ( .A1(G8), .A2(n662), .ZN(n663) );
  NAND2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n666) );
  XOR2_X1 U733 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n665) );
  XNOR2_X1 U734 ( .A(n666), .B(n665), .ZN(n675) );
  AND2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n673) );
  AND2_X1 U736 ( .A1(G8), .A2(n669), .ZN(n671) );
  OR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n688) );
  NOR2_X1 U739 ( .A1(G1976), .A2(G288), .ZN(n680) );
  NOR2_X1 U740 ( .A1(G303), .A2(G1971), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n680), .A2(n676), .ZN(n978) );
  NAND2_X1 U742 ( .A1(n688), .A2(n978), .ZN(n677) );
  XNOR2_X1 U743 ( .A(n677), .B(KEYINPUT100), .ZN(n678) );
  NAND2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n972) );
  NAND2_X1 U745 ( .A1(n678), .A2(n972), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n679), .B(KEYINPUT101), .ZN(n685) );
  XOR2_X1 U747 ( .A(G1981), .B(G305), .Z(n963) );
  INV_X1 U748 ( .A(n963), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n680), .A2(KEYINPUT33), .ZN(n681) );
  NOR2_X1 U750 ( .A1(n681), .A2(n692), .ZN(n682) );
  OR2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n695) );
  NOR2_X1 U752 ( .A1(n692), .A2(n695), .ZN(n684) );
  AND2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n700) );
  NOR2_X1 U754 ( .A1(G2090), .A2(G303), .ZN(n686) );
  NAND2_X1 U755 ( .A1(G8), .A2(n686), .ZN(n687) );
  NAND2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U757 ( .A1(n689), .A2(n692), .ZN(n694) );
  NOR2_X1 U758 ( .A1(G1981), .A2(G305), .ZN(n690) );
  XOR2_X1 U759 ( .A(n690), .B(KEYINPUT24), .Z(n691) );
  OR2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n698) );
  INV_X1 U762 ( .A(n695), .ZN(n696) );
  AND2_X1 U763 ( .A1(n696), .A2(KEYINPUT33), .ZN(n697) );
  OR2_X1 U764 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n701) );
  INV_X1 U766 ( .A(n701), .ZN(n736) );
  NAND2_X1 U767 ( .A1(G131), .A2(n703), .ZN(n706) );
  NAND2_X1 U768 ( .A1(G119), .A2(n868), .ZN(n704) );
  XOR2_X1 U769 ( .A(KEYINPUT93), .B(n704), .Z(n705) );
  NAND2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n710) );
  NAND2_X1 U771 ( .A1(G95), .A2(n864), .ZN(n708) );
  NAND2_X1 U772 ( .A1(G107), .A2(n867), .ZN(n707) );
  NAND2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n709) );
  OR2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n875) );
  AND2_X1 U775 ( .A1(n875), .A2(G1991), .ZN(n719) );
  NAND2_X1 U776 ( .A1(n868), .A2(G129), .ZN(n712) );
  NAND2_X1 U777 ( .A1(G141), .A2(n703), .ZN(n711) );
  NAND2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U779 ( .A1(n864), .A2(G105), .ZN(n713) );
  XOR2_X1 U780 ( .A(KEYINPUT38), .B(n713), .Z(n714) );
  NOR2_X1 U781 ( .A1(n715), .A2(n714), .ZN(n717) );
  NAND2_X1 U782 ( .A1(n867), .A2(G117), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n876) );
  AND2_X1 U784 ( .A1(n876), .A2(G1996), .ZN(n718) );
  NOR2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n911) );
  NOR2_X1 U786 ( .A1(n721), .A2(n720), .ZN(n747) );
  INV_X1 U787 ( .A(n747), .ZN(n722) );
  NOR2_X1 U788 ( .A1(n911), .A2(n722), .ZN(n739) );
  XOR2_X1 U789 ( .A(G1986), .B(G290), .Z(n974) );
  NAND2_X1 U790 ( .A1(n867), .A2(G116), .ZN(n723) );
  XNOR2_X1 U791 ( .A(n723), .B(KEYINPUT92), .ZN(n725) );
  NAND2_X1 U792 ( .A1(G128), .A2(n868), .ZN(n724) );
  NAND2_X1 U793 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U794 ( .A(n726), .B(KEYINPUT35), .ZN(n732) );
  XNOR2_X1 U795 ( .A(KEYINPUT91), .B(KEYINPUT34), .ZN(n730) );
  NAND2_X1 U796 ( .A1(n864), .A2(G104), .ZN(n728) );
  NAND2_X1 U797 ( .A1(G140), .A2(n703), .ZN(n727) );
  NAND2_X1 U798 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U799 ( .A(n730), .B(n729), .ZN(n731) );
  NAND2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U801 ( .A(KEYINPUT36), .B(n733), .ZN(n863) );
  XOR2_X1 U802 ( .A(G2067), .B(KEYINPUT37), .Z(n744) );
  NAND2_X1 U803 ( .A1(n863), .A2(n744), .ZN(n919) );
  NAND2_X1 U804 ( .A1(n974), .A2(n919), .ZN(n734) );
  NAND2_X1 U805 ( .A1(n736), .A2(n735), .ZN(n750) );
  NOR2_X1 U806 ( .A1(G1996), .A2(n876), .ZN(n908) );
  NOR2_X1 U807 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U808 ( .A1(G1991), .A2(n875), .ZN(n914) );
  NOR2_X1 U809 ( .A1(n737), .A2(n914), .ZN(n738) );
  NOR2_X1 U810 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U811 ( .A(n740), .B(KEYINPUT102), .ZN(n741) );
  NOR2_X1 U812 ( .A1(n908), .A2(n741), .ZN(n742) );
  XNOR2_X1 U813 ( .A(n742), .B(KEYINPUT39), .ZN(n743) );
  NAND2_X1 U814 ( .A1(n743), .A2(n919), .ZN(n746) );
  NOR2_X1 U815 ( .A1(n863), .A2(n744), .ZN(n745) );
  XNOR2_X1 U816 ( .A(KEYINPUT103), .B(n745), .ZN(n924) );
  NAND2_X1 U817 ( .A1(n746), .A2(n924), .ZN(n748) );
  NAND2_X1 U818 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U819 ( .A1(n750), .A2(n749), .ZN(n752) );
  XNOR2_X1 U820 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n751) );
  XNOR2_X1 U821 ( .A(n752), .B(n751), .ZN(G329) );
  AND2_X1 U822 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U823 ( .A(G57), .ZN(G237) );
  INV_X1 U824 ( .A(G82), .ZN(G220) );
  NAND2_X1 U825 ( .A1(G7), .A2(G661), .ZN(n753) );
  XNOR2_X1 U826 ( .A(n753), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U827 ( .A(G223), .B(KEYINPUT73), .ZN(n816) );
  NAND2_X1 U828 ( .A1(n816), .A2(G567), .ZN(n754) );
  XOR2_X1 U829 ( .A(KEYINPUT11), .B(n754), .Z(G234) );
  INV_X1 U830 ( .A(G860), .ZN(n788) );
  OR2_X1 U831 ( .A1(n968), .A2(n788), .ZN(G153) );
  INV_X1 U832 ( .A(G868), .ZN(n800) );
  NOR2_X1 U833 ( .A1(G301), .A2(n800), .ZN(n756) );
  AND2_X1 U834 ( .A1(n800), .A2(n962), .ZN(n755) );
  NOR2_X1 U835 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U836 ( .A(KEYINPUT76), .B(n757), .ZN(G284) );
  NAND2_X1 U837 ( .A1(G868), .A2(G286), .ZN(n759) );
  NAND2_X1 U838 ( .A1(G299), .A2(n800), .ZN(n758) );
  NAND2_X1 U839 ( .A1(n759), .A2(n758), .ZN(G297) );
  NAND2_X1 U840 ( .A1(n788), .A2(G559), .ZN(n760) );
  NAND2_X1 U841 ( .A1(n760), .A2(n962), .ZN(n761) );
  XNOR2_X1 U842 ( .A(n761), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U843 ( .A1(G868), .A2(n968), .ZN(n764) );
  NAND2_X1 U844 ( .A1(G868), .A2(n962), .ZN(n762) );
  NOR2_X1 U845 ( .A1(G559), .A2(n762), .ZN(n763) );
  NOR2_X1 U846 ( .A1(n764), .A2(n763), .ZN(G282) );
  NAND2_X1 U847 ( .A1(G123), .A2(n868), .ZN(n765) );
  XNOR2_X1 U848 ( .A(n765), .B(KEYINPUT18), .ZN(n768) );
  NAND2_X1 U849 ( .A1(n703), .A2(G135), .ZN(n766) );
  XOR2_X1 U850 ( .A(KEYINPUT79), .B(n766), .Z(n767) );
  NAND2_X1 U851 ( .A1(n768), .A2(n767), .ZN(n772) );
  NAND2_X1 U852 ( .A1(G99), .A2(n864), .ZN(n770) );
  NAND2_X1 U853 ( .A1(G111), .A2(n867), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U855 ( .A1(n772), .A2(n771), .ZN(n913) );
  XNOR2_X1 U856 ( .A(n913), .B(G2096), .ZN(n774) );
  INV_X1 U857 ( .A(G2100), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n774), .A2(n773), .ZN(G156) );
  NAND2_X1 U859 ( .A1(n775), .A2(G93), .ZN(n778) );
  NAND2_X1 U860 ( .A1(G80), .A2(n776), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U862 ( .A(n779), .B(KEYINPUT81), .ZN(n782) );
  NAND2_X1 U863 ( .A1(G67), .A2(n780), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U865 ( .A1(n783), .A2(G55), .ZN(n784) );
  XOR2_X1 U866 ( .A(KEYINPUT82), .B(n784), .Z(n785) );
  OR2_X1 U867 ( .A1(n786), .A2(n785), .ZN(n799) );
  XNOR2_X1 U868 ( .A(n799), .B(KEYINPUT80), .ZN(n790) );
  NAND2_X1 U869 ( .A1(G559), .A2(n962), .ZN(n787) );
  XOR2_X1 U870 ( .A(n968), .B(n787), .Z(n797) );
  NAND2_X1 U871 ( .A1(n797), .A2(n788), .ZN(n789) );
  XNOR2_X1 U872 ( .A(n790), .B(n789), .ZN(G145) );
  XOR2_X1 U873 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n792) );
  XOR2_X1 U874 ( .A(G166), .B(n799), .Z(n791) );
  XNOR2_X1 U875 ( .A(n792), .B(n791), .ZN(n793) );
  XNOR2_X1 U876 ( .A(n793), .B(G299), .ZN(n794) );
  XNOR2_X1 U877 ( .A(n794), .B(G305), .ZN(n795) );
  XNOR2_X1 U878 ( .A(n795), .B(G288), .ZN(n796) );
  XNOR2_X1 U879 ( .A(n796), .B(G290), .ZN(n886) );
  XNOR2_X1 U880 ( .A(n797), .B(n886), .ZN(n798) );
  NAND2_X1 U881 ( .A1(n798), .A2(G868), .ZN(n802) );
  NAND2_X1 U882 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U883 ( .A1(n802), .A2(n801), .ZN(G295) );
  NAND2_X1 U884 ( .A1(G2078), .A2(G2084), .ZN(n803) );
  XOR2_X1 U885 ( .A(KEYINPUT20), .B(n803), .Z(n804) );
  NAND2_X1 U886 ( .A1(G2090), .A2(n804), .ZN(n805) );
  XNOR2_X1 U887 ( .A(KEYINPUT21), .B(n805), .ZN(n806) );
  NAND2_X1 U888 ( .A1(n806), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U889 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U890 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  NAND2_X1 U891 ( .A1(G483), .A2(G661), .ZN(n814) );
  NOR2_X1 U892 ( .A1(G219), .A2(G220), .ZN(n807) );
  XOR2_X1 U893 ( .A(KEYINPUT22), .B(n807), .Z(n808) );
  NOR2_X1 U894 ( .A1(G218), .A2(n808), .ZN(n809) );
  NAND2_X1 U895 ( .A1(G96), .A2(n809), .ZN(n821) );
  NAND2_X1 U896 ( .A1(n821), .A2(G2106), .ZN(n813) );
  NAND2_X1 U897 ( .A1(G69), .A2(G120), .ZN(n810) );
  NOR2_X1 U898 ( .A1(G237), .A2(n810), .ZN(n811) );
  NAND2_X1 U899 ( .A1(G108), .A2(n811), .ZN(n820) );
  NAND2_X1 U900 ( .A1(n820), .A2(G567), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n813), .A2(n812), .ZN(n823) );
  NOR2_X1 U902 ( .A1(n814), .A2(n823), .ZN(n815) );
  XNOR2_X1 U903 ( .A(n815), .B(KEYINPUT86), .ZN(n819) );
  NAND2_X1 U904 ( .A1(G36), .A2(n819), .ZN(G176) );
  NAND2_X1 U905 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U906 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U907 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U908 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(G188) );
  INV_X1 U911 ( .A(G120), .ZN(G236) );
  INV_X1 U912 ( .A(G96), .ZN(G221) );
  INV_X1 U913 ( .A(G69), .ZN(G235) );
  NOR2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U915 ( .A(n822), .B(KEYINPUT106), .ZN(G325) );
  INV_X1 U916 ( .A(G325), .ZN(G261) );
  INV_X1 U917 ( .A(n823), .ZN(G319) );
  XOR2_X1 U918 ( .A(KEYINPUT107), .B(G2084), .Z(n825) );
  XNOR2_X1 U919 ( .A(G2067), .B(G2078), .ZN(n824) );
  XNOR2_X1 U920 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U921 ( .A(n826), .B(G2100), .Z(n828) );
  XNOR2_X1 U922 ( .A(G2072), .B(G2090), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U924 ( .A(G2096), .B(KEYINPUT43), .Z(n830) );
  XNOR2_X1 U925 ( .A(KEYINPUT42), .B(G2678), .ZN(n829) );
  XNOR2_X1 U926 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U927 ( .A(n832), .B(n831), .Z(G227) );
  XOR2_X1 U928 ( .A(G1991), .B(G1981), .Z(n834) );
  XNOR2_X1 U929 ( .A(G1966), .B(G1996), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n844) );
  XOR2_X1 U931 ( .A(G2474), .B(KEYINPUT110), .Z(n836) );
  XNOR2_X1 U932 ( .A(G1956), .B(KEYINPUT41), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U934 ( .A(G1986), .B(G1976), .Z(n838) );
  XNOR2_X1 U935 ( .A(G1961), .B(G1971), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U937 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U938 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(G229) );
  NAND2_X1 U941 ( .A1(G124), .A2(n868), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n845), .B(KEYINPUT44), .ZN(n847) );
  NAND2_X1 U943 ( .A1(n864), .A2(G100), .ZN(n846) );
  NAND2_X1 U944 ( .A1(n847), .A2(n846), .ZN(n851) );
  NAND2_X1 U945 ( .A1(n867), .A2(G112), .ZN(n849) );
  NAND2_X1 U946 ( .A1(G136), .A2(n703), .ZN(n848) );
  NAND2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U948 ( .A1(n851), .A2(n850), .ZN(G162) );
  NAND2_X1 U949 ( .A1(G118), .A2(n867), .ZN(n853) );
  NAND2_X1 U950 ( .A1(G130), .A2(n868), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n858) );
  NAND2_X1 U952 ( .A1(n864), .A2(G106), .ZN(n855) );
  NAND2_X1 U953 ( .A1(G142), .A2(n703), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n856), .B(KEYINPUT45), .Z(n857) );
  NOR2_X1 U956 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n859), .B(G160), .ZN(n882) );
  XOR2_X1 U958 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n861) );
  XNOR2_X1 U959 ( .A(n913), .B(G162), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n880) );
  NAND2_X1 U962 ( .A1(n864), .A2(G103), .ZN(n866) );
  NAND2_X1 U963 ( .A1(G139), .A2(n703), .ZN(n865) );
  NAND2_X1 U964 ( .A1(n866), .A2(n865), .ZN(n873) );
  NAND2_X1 U965 ( .A1(G115), .A2(n867), .ZN(n870) );
  NAND2_X1 U966 ( .A1(G127), .A2(n868), .ZN(n869) );
  NAND2_X1 U967 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U968 ( .A(KEYINPUT47), .B(n871), .Z(n872) );
  NOR2_X1 U969 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U970 ( .A(KEYINPUT111), .B(n874), .Z(n926) );
  XNOR2_X1 U971 ( .A(n926), .B(n875), .ZN(n878) );
  XOR2_X1 U972 ( .A(G164), .B(n876), .Z(n877) );
  XNOR2_X1 U973 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U974 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U975 ( .A(n882), .B(n881), .Z(n883) );
  NOR2_X1 U976 ( .A1(G37), .A2(n883), .ZN(G395) );
  XNOR2_X1 U977 ( .A(G286), .B(KEYINPUT112), .ZN(n885) );
  XNOR2_X1 U978 ( .A(n962), .B(G171), .ZN(n884) );
  XNOR2_X1 U979 ( .A(n885), .B(n884), .ZN(n888) );
  XNOR2_X1 U980 ( .A(n968), .B(n886), .ZN(n887) );
  XNOR2_X1 U981 ( .A(n888), .B(n887), .ZN(n889) );
  NOR2_X1 U982 ( .A1(G37), .A2(n889), .ZN(n890) );
  XOR2_X1 U983 ( .A(KEYINPUT113), .B(n890), .Z(G397) );
  XOR2_X1 U984 ( .A(G2454), .B(G2435), .Z(n892) );
  XNOR2_X1 U985 ( .A(G2438), .B(G2427), .ZN(n891) );
  XNOR2_X1 U986 ( .A(n892), .B(n891), .ZN(n899) );
  XOR2_X1 U987 ( .A(KEYINPUT105), .B(G2446), .Z(n894) );
  XNOR2_X1 U988 ( .A(G2443), .B(G2430), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U990 ( .A(n895), .B(G2451), .Z(n897) );
  XNOR2_X1 U991 ( .A(G1341), .B(G1348), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n900) );
  NAND2_X1 U994 ( .A1(n900), .A2(G14), .ZN(n906) );
  NAND2_X1 U995 ( .A1(G319), .A2(n906), .ZN(n903) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n901) );
  XNOR2_X1 U997 ( .A(KEYINPUT49), .B(n901), .ZN(n902) );
  NOR2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n905) );
  NOR2_X1 U999 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1001 ( .A(G225), .ZN(G308) );
  INV_X1 U1002 ( .A(G108), .ZN(G238) );
  INV_X1 U1003 ( .A(n906), .ZN(G401) );
  XOR2_X1 U1004 ( .A(G2090), .B(G162), .Z(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n909), .B(KEYINPUT51), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n910), .B(KEYINPUT117), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n923) );
  NOR2_X1 U1009 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1010 ( .A(KEYINPUT114), .B(n915), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(G160), .B(G2084), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1013 ( .A(KEYINPUT115), .B(n918), .ZN(n920) );
  NAND2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(KEYINPUT116), .B(n921), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(n923), .A2(n922), .ZN(n925) );
  NAND2_X1 U1017 ( .A1(n925), .A2(n924), .ZN(n932) );
  XOR2_X1 U1018 ( .A(G2072), .B(n926), .Z(n928) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n927) );
  NOR2_X1 U1020 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1021 ( .A(KEYINPUT118), .B(n929), .Z(n930) );
  XNOR2_X1 U1022 ( .A(KEYINPUT50), .B(n930), .ZN(n931) );
  NOR2_X1 U1023 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1024 ( .A(KEYINPUT52), .B(n933), .Z(n934) );
  NOR2_X1 U1025 ( .A1(KEYINPUT55), .A2(n934), .ZN(n935) );
  XNOR2_X1 U1026 ( .A(KEYINPUT119), .B(n935), .ZN(n936) );
  NAND2_X1 U1027 ( .A1(n936), .A2(G29), .ZN(n1015) );
  XNOR2_X1 U1028 ( .A(G25), .B(G1991), .ZN(n937) );
  XNOR2_X1 U1029 ( .A(n937), .B(KEYINPUT121), .ZN(n949) );
  XNOR2_X1 U1030 ( .A(G32), .B(n938), .ZN(n939) );
  NAND2_X1 U1031 ( .A1(n939), .A2(G28), .ZN(n947) );
  XOR2_X1 U1032 ( .A(n940), .B(G27), .Z(n945) );
  XNOR2_X1 U1033 ( .A(G2072), .B(G33), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(G26), .B(G2067), .ZN(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(n943), .B(KEYINPUT122), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1038 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1039 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(n950), .B(KEYINPUT53), .ZN(n953) );
  XOR2_X1 U1041 ( .A(G2084), .B(G34), .Z(n951) );
  XNOR2_X1 U1042 ( .A(KEYINPUT54), .B(n951), .ZN(n952) );
  NAND2_X1 U1043 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1044 ( .A(KEYINPUT120), .B(G2090), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(G35), .B(n954), .ZN(n955) );
  NOR2_X1 U1046 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(KEYINPUT55), .B(n957), .ZN(n959) );
  INV_X1 U1048 ( .A(G29), .ZN(n958) );
  NAND2_X1 U1049 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1050 ( .A1(n960), .A2(G11), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(n961), .B(KEYINPUT123), .ZN(n986) );
  XNOR2_X1 U1052 ( .A(KEYINPUT56), .B(G16), .ZN(n984) );
  XNOR2_X1 U1053 ( .A(n962), .B(G1348), .ZN(n967) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n964) );
  NAND2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(n965), .B(KEYINPUT57), .ZN(n966) );
  NAND2_X1 U1057 ( .A1(n967), .A2(n966), .ZN(n970) );
  XNOR2_X1 U1058 ( .A(G1341), .B(n968), .ZN(n969) );
  NOR2_X1 U1059 ( .A1(n970), .A2(n969), .ZN(n982) );
  XOR2_X1 U1060 ( .A(G1956), .B(G299), .Z(n971) );
  NAND2_X1 U1061 ( .A1(n972), .A2(n971), .ZN(n980) );
  NAND2_X1 U1062 ( .A1(G303), .A2(G1971), .ZN(n973) );
  NAND2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1064 ( .A(G1961), .B(G301), .ZN(n975) );
  NOR2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1066 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1067 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1068 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1069 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1070 ( .A1(n986), .A2(n985), .ZN(n1012) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G21), .ZN(n988) );
  XNOR2_X1 U1072 ( .A(G5), .B(G1961), .ZN(n987) );
  NOR2_X1 U1073 ( .A1(n988), .A2(n987), .ZN(n998) );
  XOR2_X1 U1074 ( .A(G1348), .B(KEYINPUT59), .Z(n989) );
  XNOR2_X1 U1075 ( .A(G4), .B(n989), .ZN(n991) );
  XNOR2_X1 U1076 ( .A(G20), .B(G1956), .ZN(n990) );
  NOR2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n995) );
  XNOR2_X1 U1078 ( .A(G1341), .B(G19), .ZN(n993) );
  XNOR2_X1 U1079 ( .A(G1981), .B(G6), .ZN(n992) );
  NOR2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1082 ( .A(KEYINPUT60), .B(n996), .Z(n997) );
  NAND2_X1 U1083 ( .A1(n998), .A2(n997), .ZN(n1006) );
  XNOR2_X1 U1084 ( .A(G1971), .B(G22), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(G23), .B(G1976), .ZN(n999) );
  NOR2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XNOR2_X1 U1087 ( .A(G1986), .B(KEYINPUT125), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(n1001), .B(G24), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(KEYINPUT58), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1091 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1092 ( .A(KEYINPUT61), .B(n1007), .Z(n1009) );
  XNOR2_X1 U1093 ( .A(G16), .B(KEYINPUT124), .ZN(n1008) );
  NOR2_X1 U1094 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(n1010), .B(KEYINPUT126), .ZN(n1011) );
  NOR2_X1 U1096 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1097 ( .A(KEYINPUT127), .B(n1013), .Z(n1014) );
  NAND2_X1 U1098 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1099 ( .A(KEYINPUT62), .B(n1016), .Z(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

