//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n626, new_n629, new_n631, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(new_n455), .B(KEYINPUT65), .Z(G261));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT66), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n465), .B(KEYINPUT67), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT3), .B1(new_n469), .B2(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n472), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n467), .B1(new_n462), .B2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n470), .A2(new_n473), .A3(KEYINPUT69), .ZN(new_n481));
  AOI21_X1  g056(.A(KEYINPUT69), .B1(new_n470), .B2(new_n473), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n462), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n480), .B1(new_n484), .B2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n481), .A2(new_n482), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(new_n462), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND3_X1  g065(.A1(new_n463), .A2(G138), .A3(new_n462), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n470), .A2(new_n473), .A3(G126), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n462), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n491), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(G102), .A2(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT4), .A2(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n474), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(new_n462), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT6), .B1(new_n506), .B2(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n507), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n510), .A2(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n510), .A2(new_n511), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n518), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT7), .Z(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n516), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n523), .B1(new_n529), .B2(G89), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n514), .B1(new_n513), .B2(G651), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n506), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT73), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n512), .A2(new_n515), .A3(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n533), .A2(G51), .A3(G543), .A4(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n536), .A2(KEYINPUT74), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(KEYINPUT74), .B1(new_n536), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n530), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g117(.A(KEYINPUT75), .B(new_n530), .C1(new_n538), .C2(new_n539), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n506), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n524), .B1(new_n516), .B2(KEYINPUT73), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n547), .A2(G52), .A3(new_n535), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT76), .B(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n529), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n546), .A2(new_n548), .A3(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND2_X1  g127(.A1(new_n547), .A2(new_n535), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n528), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  INV_X1    g134(.A(new_n529), .ZN(new_n560));
  INV_X1    g135(.A(G81), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(G188));
  NOR2_X1   g144(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n553), .B2(new_n571), .ZN(new_n572));
  XOR2_X1   g147(.A(KEYINPUT77), .B(KEYINPUT9), .Z(new_n573));
  NAND4_X1  g148(.A1(new_n547), .A2(G53), .A3(new_n535), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n528), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(G91), .A2(new_n529), .B1(new_n577), .B2(G651), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n572), .A2(new_n574), .A3(new_n578), .ZN(G299));
  INV_X1    g154(.A(G168), .ZN(G286));
  OAI21_X1  g155(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n507), .A2(G87), .A3(new_n512), .A4(new_n515), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n533), .A2(G49), .A3(G543), .A4(new_n535), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(KEYINPUT78), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n547), .A2(new_n586), .A3(G49), .A4(new_n535), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n528), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(G48), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n528), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n531), .A2(new_n532), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT79), .ZN(G305));
  NAND3_X1  g174(.A1(new_n525), .A2(new_n527), .A3(G60), .ZN(new_n600));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n529), .A2(G85), .B1(new_n602), .B2(G651), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n533), .A2(G47), .A3(G543), .A4(new_n535), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n596), .A2(G92), .A3(new_n507), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(KEYINPUT80), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n529), .A2(new_n609), .A3(G92), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n553), .A2(KEYINPUT81), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n547), .A2(new_n615), .A3(new_n535), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n614), .A2(G54), .A3(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(new_n506), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n608), .A2(KEYINPUT10), .A3(new_n610), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n613), .A2(new_n617), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n606), .B1(new_n622), .B2(G868), .ZN(G284));
  OAI21_X1  g198(.A(new_n606), .B1(new_n622), .B2(G868), .ZN(G321));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(G299), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G168), .B2(new_n625), .ZN(G297));
  OAI21_X1  g202(.A(new_n626), .B1(G168), .B2(new_n625), .ZN(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n622), .B1(new_n629), .B2(G860), .ZN(G148));
  OAI221_X1 g205(.A(new_n559), .B1(new_n560), .B2(new_n561), .C1(new_n553), .C2(new_n554), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n625), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n621), .A2(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n625), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g210(.A1(new_n469), .A2(G2105), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n463), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2100), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n487), .A2(G123), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n484), .A2(G135), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n462), .A2(G111), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(G2096), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n640), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT82), .Z(G156));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT84), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT15), .B(G2435), .Z(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2443), .B(G2446), .Z(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT17), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XOR2_X1   g245(.A(G2067), .B(G2678), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT86), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n671), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n670), .B1(new_n668), .B2(new_n671), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n674), .B1(KEYINPUT85), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(KEYINPUT85), .B2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(new_n670), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n679), .A2(new_n668), .A3(new_n671), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT18), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n673), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2096), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT87), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n690), .A2(new_n691), .A3(KEYINPUT89), .ZN(new_n692));
  OAI21_X1  g267(.A(KEYINPUT89), .B1(new_n690), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1971), .B(G1976), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT19), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n688), .A2(new_n695), .A3(new_n689), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT88), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n688), .A2(new_n689), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(new_n695), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n696), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1991), .ZN(new_n704));
  INV_X1    g279(.A(G1996), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n703), .A2(G1991), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n703), .A2(G1991), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n709), .A2(G1996), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n706), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n708), .B1(new_n706), .B2(new_n711), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n686), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n714), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n716), .A2(new_n685), .A3(new_n712), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n717), .ZN(G229));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G6), .ZN(new_n720));
  INV_X1    g295(.A(G305), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT32), .B(G1981), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G288), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G16), .B2(G23), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT33), .B(G1976), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n719), .A2(G22), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G166), .B2(new_n719), .ZN(new_n731));
  INV_X1    g306(.A(G1971), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n727), .A2(new_n728), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n724), .A2(new_n729), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT34), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT34), .ZN(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G24), .ZN(new_n738));
  XNOR2_X1  g313(.A(G290), .B(KEYINPUT93), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1986), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G25), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(KEYINPUT90), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(KEYINPUT90), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n487), .A2(G119), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n487), .A2(KEYINPUT91), .A3(G119), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G107), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n484), .B2(G131), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n748), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n744), .B(new_n745), .C1(new_n754), .C2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT35), .B(G1991), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT92), .Z(new_n757));
  AND2_X1   g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n755), .A2(new_n757), .ZN(new_n759));
  NOR4_X1   g334(.A1(new_n741), .A2(new_n758), .A3(new_n759), .A4(KEYINPUT94), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n736), .A2(new_n737), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NOR2_X1   g339(.A1(G16), .A2(G21), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G168), .B2(G16), .ZN(new_n766));
  INV_X1    g341(.A(G1966), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n742), .A2(G35), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G162), .B2(new_n742), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT29), .Z(new_n771));
  INV_X1    g346(.A(G2090), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n742), .A2(G32), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n487), .A2(G129), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n484), .A2(G141), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT26), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n779), .A2(new_n780), .B1(G105), .B2(new_n636), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n775), .A2(new_n776), .A3(new_n781), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT99), .Z(new_n783));
  OAI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(new_n742), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT27), .B(G1996), .Z(new_n785));
  AOI22_X1  g360(.A1(new_n771), .A2(new_n772), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n742), .A2(G33), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n636), .A2(G103), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT25), .Z(new_n789));
  AOI22_X1  g364(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n790));
  INV_X1    g365(.A(G139), .ZN(new_n791));
  OAI221_X1 g366(.A(new_n789), .B1(new_n462), .B2(new_n790), .C1(new_n483), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT97), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n787), .B1(new_n793), .B2(new_n742), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT98), .B(G2072), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n773), .A2(new_n786), .A3(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT23), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n719), .A2(G20), .ZN(new_n799));
  AOI211_X1 g374(.A(new_n798), .B(new_n799), .C1(G299), .C2(G16), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n798), .B2(new_n799), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT101), .B(G1956), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n785), .B2(new_n784), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n719), .A2(G4), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n622), .B2(new_n719), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT95), .B(G1348), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT24), .ZN(new_n809));
  INV_X1    g384(.A(G34), .ZN(new_n810));
  AOI21_X1  g385(.A(G29), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n809), .B2(new_n810), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G160), .B2(new_n742), .ZN(new_n813));
  INV_X1    g388(.A(G2084), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT31), .B(G11), .Z(new_n816));
  XOR2_X1   g391(.A(KEYINPUT100), .B(KEYINPUT30), .Z(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(G28), .ZN(new_n818));
  AOI21_X1  g393(.A(G29), .B1(new_n817), .B2(G28), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n815), .B(new_n820), .C1(new_n742), .C2(new_n645), .ZN(new_n821));
  NAND2_X1  g396(.A1(G164), .A2(G29), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G27), .B2(G29), .ZN(new_n823));
  INV_X1    g398(.A(G2078), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n821), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n719), .A2(G19), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n563), .B2(new_n719), .ZN(new_n829));
  INV_X1    g404(.A(G1341), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(G5), .A2(G16), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G171), .B2(G16), .ZN(new_n833));
  INV_X1    g408(.A(G1961), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n808), .A2(new_n827), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n742), .A2(G26), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n838));
  INV_X1    g413(.A(G116), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(G2105), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n487), .B2(G128), .ZN(new_n841));
  INV_X1    g416(.A(G140), .ZN(new_n842));
  OR3_X1    g417(.A1(new_n483), .A2(KEYINPUT96), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT96), .B1(new_n483), .B2(new_n842), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n837), .B1(new_n845), .B2(G29), .ZN(new_n846));
  MUX2_X1   g421(.A(new_n837), .B(new_n846), .S(KEYINPUT28), .Z(new_n847));
  INV_X1    g422(.A(G2067), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NOR4_X1   g424(.A1(new_n797), .A2(new_n804), .A3(new_n836), .A4(new_n849), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n763), .A2(new_n764), .A3(new_n768), .A4(new_n850), .ZN(G150));
  INV_X1    g426(.A(G150), .ZN(G311));
  NAND2_X1  g427(.A1(new_n622), .A2(G559), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n533), .A2(G55), .A3(G543), .A4(new_n535), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n529), .A2(G93), .ZN(new_n855));
  NAND2_X1  g430(.A1(G80), .A2(G543), .ZN(new_n856));
  INV_X1    g431(.A(G67), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n528), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(G651), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n854), .A2(new_n855), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT103), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n860), .A2(KEYINPUT103), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n631), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n854), .A2(new_n855), .A3(new_n859), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n631), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n563), .A2(KEYINPUT102), .A3(new_n860), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n853), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n872));
  AOI21_X1  g447(.A(G860), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n872), .B2(new_n871), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n862), .A2(new_n863), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G860), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT37), .Z(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT104), .ZN(G145));
  NAND2_X1  g454(.A1(new_n476), .A2(new_n462), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n464), .A2(new_n466), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n462), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n845), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n645), .A2(new_n489), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n489), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT105), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n887), .A2(KEYINPUT105), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n887), .A2(KEYINPUT105), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n888), .A3(new_n883), .ZN(new_n893));
  INV_X1    g468(.A(new_n782), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n793), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(new_n783), .B2(new_n793), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n891), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n891), .B2(new_n893), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n484), .A2(G142), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n462), .A2(G118), .ZN(new_n901));
  OAI21_X1  g476(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n903), .B1(G130), .B2(new_n487), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(G164), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n754), .B(new_n638), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n898), .A2(new_n899), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n908), .B1(new_n898), .B2(new_n899), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g488(.A(KEYINPUT111), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n602), .A2(G651), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n507), .A2(G85), .A3(new_n512), .A4(new_n515), .ZN(new_n917));
  AND4_X1   g492(.A1(new_n915), .A2(new_n604), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n603), .B2(new_n604), .ZN(new_n919));
  OAI21_X1  g494(.A(G288), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n604), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(new_n917), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT108), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n603), .A2(new_n915), .A3(new_n604), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n923), .A2(new_n587), .A3(new_n585), .A4(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n920), .A2(new_n925), .A3(G305), .ZN(new_n926));
  AOI21_X1  g501(.A(G305), .B1(new_n920), .B2(new_n925), .ZN(new_n927));
  NOR3_X1   g502(.A1(new_n926), .A2(new_n927), .A3(G303), .ZN(new_n928));
  NOR3_X1   g503(.A1(G288), .A2(new_n918), .A3(new_n919), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n923), .A2(new_n924), .B1(new_n587), .B2(new_n585), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n721), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n920), .A2(new_n925), .A3(G305), .ZN(new_n932));
  AOI21_X1  g507(.A(G166), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n928), .A2(new_n933), .A3(KEYINPUT42), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n928), .B2(new_n933), .ZN(new_n936));
  OAI21_X1  g511(.A(G303), .B1(new_n926), .B2(new_n927), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n931), .A2(G166), .A3(new_n932), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(KEYINPUT109), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n934), .B1(new_n940), .B2(KEYINPUT42), .ZN(new_n941));
  INV_X1    g516(.A(G299), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT106), .B1(new_n621), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n620), .A2(new_n619), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT10), .B1(new_n608), .B2(new_n610), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n946), .A2(new_n947), .A3(G299), .A4(new_n617), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n621), .A2(new_n942), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT41), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n621), .A2(KEYINPUT107), .A3(new_n942), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n953), .A2(new_n954), .B1(new_n943), .B2(new_n948), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n951), .B1(new_n955), .B2(KEYINPUT41), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n869), .A2(new_n633), .ZN(new_n957));
  INV_X1    g532(.A(new_n944), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n958), .A2(new_n629), .A3(new_n617), .A4(new_n613), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(new_n864), .A3(new_n867), .A4(new_n868), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n956), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n949), .A2(new_n950), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT110), .B1(new_n941), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n961), .A2(new_n964), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n962), .B2(new_n956), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n936), .B2(new_n939), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n969), .B(new_n970), .C1(new_n972), .C2(new_n934), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n941), .A2(new_n966), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n967), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G868), .ZN(new_n976));
  INV_X1    g551(.A(new_n875), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(G868), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n914), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  AOI211_X1 g555(.A(KEYINPUT111), .B(new_n978), .C1(new_n975), .C2(G868), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(G295));
  NAND2_X1  g557(.A1(new_n976), .A2(new_n979), .ZN(G331));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n985));
  AOI21_X1  g560(.A(G301), .B1(new_n542), .B2(new_n543), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n542), .A2(new_n543), .A3(G301), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n988), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n990), .A2(new_n869), .A3(new_n986), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n964), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT112), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n989), .A2(new_n991), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n956), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n996), .B(new_n964), .C1(new_n989), .C2(new_n991), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n993), .A2(new_n995), .A3(new_n940), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n910), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n992), .A2(KEYINPUT112), .B1(new_n994), .B2(new_n956), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n940), .B1(new_n1000), .B2(new_n997), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n984), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n964), .B1(new_n994), .B2(KEYINPUT41), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n869), .B1(new_n990), .B2(new_n986), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n987), .A2(new_n985), .A3(new_n988), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(new_n1005), .A3(KEYINPUT41), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(new_n955), .ZN(new_n1007));
  OR3_X1    g582(.A1(new_n1003), .A2(new_n940), .A3(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1008), .A2(KEYINPUT43), .A3(new_n998), .A4(new_n910), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT44), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT43), .B1(new_n999), .B2(new_n1001), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1008), .A2(new_n984), .A3(new_n998), .A4(new_n910), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1011), .A2(new_n1016), .ZN(G397));
  AOI21_X1  g592(.A(G1384), .B1(new_n499), .B2(new_n503), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(KEYINPUT45), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G160), .A2(G40), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n705), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n845), .B(new_n848), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1023), .B(new_n1024), .C1(new_n705), .C2(new_n894), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n754), .B(new_n756), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1022), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1022), .ZN(new_n1028));
  XOR2_X1   g603(.A(G290), .B(G1986), .Z(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT113), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n598), .B(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n592), .A2(KEYINPUT116), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G1981), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1032), .B(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G40), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n882), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n1018), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G8), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1039), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n725), .A2(G1976), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n725), .B2(G1976), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1041), .B(new_n1045), .C1(KEYINPUT52), .C2(new_n1042), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1040), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1018), .A2(KEYINPUT45), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1037), .B1(new_n1018), .B2(KEYINPUT45), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n767), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1384), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n504), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT50), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1018), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1058), .A3(new_n1037), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1053), .B1(G2084), .B2(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1060), .A2(G8), .A3(G168), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT45), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1021), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1018), .A2(new_n1064), .A3(KEYINPUT45), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n1018), .B2(KEYINPUT45), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1058), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1037), .B1(new_n1018), .B2(new_n1057), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1067), .A2(new_n732), .B1(new_n1070), .B2(new_n772), .ZN(new_n1071));
  INV_X1    g646(.A(G8), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G303), .A2(G8), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1075), .B(new_n1076), .C1(KEYINPUT120), .C2(new_n1072), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1071), .A2(new_n1072), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1072), .A2(KEYINPUT120), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1050), .A2(KEYINPUT114), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1018), .A2(new_n1064), .A3(KEYINPUT45), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1052), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1084), .A2(G1971), .B1(G2090), .B2(new_n1059), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1081), .B1(new_n1085), .B2(G8), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1049), .B(new_n1061), .C1(new_n1078), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT121), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1077), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1085), .A2(new_n1081), .A3(G8), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n1049), .A4(new_n1061), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1088), .A2(new_n1089), .A3(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1049), .B1(new_n1096), .B2(new_n1079), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT122), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1061), .A2(KEYINPUT63), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1096), .B2(new_n1079), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1049), .B(new_n1101), .C1(new_n1096), .C2(new_n1079), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1095), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1049), .A2(new_n1096), .A3(new_n1079), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1039), .B(KEYINPUT117), .Z(new_n1106));
  NOR2_X1   g681(.A1(G288), .A2(G1976), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT118), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1040), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n598), .A2(G1981), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1106), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1105), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT119), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1104), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1092), .A2(new_n1049), .ZN(new_n1115));
  XNOR2_X1  g690(.A(G299), .B(KEYINPUT57), .ZN(new_n1116));
  XOR2_X1   g691(.A(new_n1116), .B(KEYINPUT123), .Z(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT56), .B(G2072), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1063), .B(new_n1118), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(G1956), .B2(new_n1070), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1116), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1119), .B(new_n1121), .C1(G1956), .C2(new_n1070), .ZN(new_n1122));
  INV_X1    g697(.A(G1348), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1059), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1038), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n848), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n621), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1117), .A2(new_n1120), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n621), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1126), .B(new_n1130), .C1(new_n1070), .C2(G1348), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n622), .A2(KEYINPUT60), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1124), .A2(KEYINPUT60), .A3(new_n1126), .A4(new_n622), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT124), .B(KEYINPUT58), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(new_n830), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1084), .A2(new_n705), .B1(new_n1038), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1136), .B1(new_n1139), .B2(new_n631), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1122), .A2(KEYINPUT61), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1038), .A2(new_n1138), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1067), .B2(G1996), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(KEYINPUT59), .A3(new_n563), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1135), .A2(new_n1140), .A3(new_n1141), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1120), .A2(new_n1116), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT61), .B1(new_n1146), .B2(new_n1122), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1128), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT51), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1149), .B(G8), .C1(new_n1060), .C2(G286), .ZN(new_n1150));
  NOR2_X1   g725(.A1(G168), .A2(new_n1072), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1060), .A2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1149), .B(new_n1151), .C1(new_n1060), .C2(G8), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1067), .B2(G2078), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1059), .A2(new_n834), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n880), .A2(KEYINPUT126), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n880), .A2(KEYINPUT126), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n824), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1162));
  NOR4_X1   g737(.A1(new_n1160), .A2(new_n1161), .A3(new_n467), .A4(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1020), .B(new_n1163), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1158), .A2(new_n1159), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1156), .B1(new_n1165), .B2(G171), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1063), .A2(KEYINPUT53), .A3(new_n824), .A4(new_n1050), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1158), .A2(G301), .A3(new_n1159), .A4(new_n1167), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1153), .A2(new_n1155), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(KEYINPUT125), .B(KEYINPUT54), .Z(new_n1170));
  AND2_X1   g745(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1171));
  AOI21_X1  g746(.A(G301), .B1(new_n1171), .B2(new_n1167), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1165), .A2(G171), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1170), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1148), .A2(new_n1169), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1176));
  OR3_X1    g751(.A1(new_n1176), .A2(new_n1154), .A3(KEYINPUT62), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT62), .B1(new_n1176), .B2(new_n1154), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(new_n1178), .A3(new_n1172), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1115), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1031), .B1(new_n1114), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1028), .B1(new_n1024), .B2(new_n894), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT46), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1182), .B1(KEYINPUT127), .B2(new_n1183), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1028), .A2(G1996), .B1(KEYINPUT127), .B2(new_n1183), .ZN(new_n1185));
  OR4_X1    g760(.A1(KEYINPUT127), .A2(new_n1028), .A3(new_n1183), .A4(G1996), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT47), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1028), .A2(G1986), .A3(G290), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT48), .Z(new_n1190));
  OR2_X1    g765(.A1(new_n754), .A2(new_n756), .ZN(new_n1191));
  OAI22_X1  g766(.A1(new_n1025), .A2(new_n1191), .B1(G2067), .B2(new_n845), .ZN(new_n1192));
  AOI22_X1  g767(.A1(new_n1190), .A2(new_n1027), .B1(new_n1022), .B2(new_n1192), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1188), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1181), .A2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g770(.A(G319), .ZN(new_n1197));
  OR3_X1    g771(.A1(G401), .A2(new_n1197), .A3(G227), .ZN(new_n1198));
  NOR2_X1   g772(.A1(G229), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n1199), .A2(new_n1014), .A3(new_n912), .ZN(G225));
  INV_X1    g774(.A(G225), .ZN(G308));
endmodule


