//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n190), .B2(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n192), .A2(new_n189), .A3(KEYINPUT75), .A4(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G140), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n190), .A2(new_n196), .A3(KEYINPUT16), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT74), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT74), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT16), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(new_n198), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n194), .A2(new_n198), .A3(new_n201), .A4(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT87), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  INV_X1    g023(.A(G237), .ZN(new_n210));
  INV_X1    g024(.A(G953), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G143), .A4(G214), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(G143), .ZN(new_n213));
  INV_X1    g027(.A(G214), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n214), .A2(G237), .A3(G953), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n209), .B(new_n212), .C1(new_n213), .C2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT84), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n212), .B1(new_n213), .B2(new_n215), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT64), .A2(G143), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT64), .A2(G143), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n210), .A2(new_n211), .A3(G214), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT84), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n224), .A2(new_n225), .A3(new_n209), .A4(new_n212), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n217), .A2(new_n219), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT17), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n204), .A2(KEYINPUT87), .A3(new_n205), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n218), .A2(KEYINPUT17), .A3(G131), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n208), .A2(new_n229), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G113), .B(G122), .ZN(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n233), .B(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n199), .A2(new_n203), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT76), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(new_n203), .B2(new_n199), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT18), .A2(G131), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n218), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n232), .A2(new_n235), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n235), .B1(new_n232), .B2(new_n242), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n187), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G475), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT20), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n232), .A2(new_n235), .A3(new_n242), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n217), .A2(new_n226), .A3(new_n219), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT85), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT85), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n217), .A2(new_n226), .A3(new_n219), .A4(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT86), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n199), .A2(new_n253), .A3(KEYINPUT19), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT19), .B1(new_n199), .B2(new_n253), .ZN(new_n255));
  OR2_X1    g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n203), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n250), .A2(new_n205), .A3(new_n252), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n242), .ZN(new_n259));
  INV_X1    g073(.A(new_n235), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n248), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(G475), .A2(G902), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n247), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n263), .ZN(new_n265));
  AOI211_X1 g079(.A(KEYINPUT20), .B(new_n265), .C1(new_n248), .C2(new_n261), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n246), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G478), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT15), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(KEYINPUT89), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(KEYINPUT89), .B2(new_n269), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G122), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G116), .ZN(new_n274));
  INV_X1    g088(.A(G116), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G122), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT88), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT88), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n274), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G107), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n275), .A2(KEYINPUT14), .A3(G122), .ZN(new_n284));
  OAI211_X1 g098(.A(G107), .B(new_n284), .C1(new_n277), .C2(KEYINPUT14), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT65), .B(G128), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G143), .ZN(new_n287));
  INV_X1    g101(.A(G134), .ZN(new_n288));
  OR2_X1    g102(.A1(KEYINPUT64), .A2(G143), .ZN(new_n289));
  NAND2_X1  g103(.A1(KEYINPUT64), .A2(G143), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(G128), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n288), .B1(new_n287), .B2(new_n291), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n283), .B(new_n285), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT9), .B(G234), .ZN(new_n296));
  INV_X1    g110(.A(G217), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n296), .A2(new_n297), .A3(G953), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n281), .A2(new_n282), .ZN(new_n300));
  AOI21_X1  g114(.A(G107), .B1(new_n278), .B2(new_n280), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n292), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT13), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n291), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n222), .A2(KEYINPUT13), .A3(G128), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n287), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G134), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n295), .B(new_n299), .C1(new_n302), .C2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n307), .B(new_n292), .C1(new_n300), .C2(new_n301), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n299), .B1(new_n311), .B2(new_n295), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT90), .B1(new_n313), .B2(new_n187), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n295), .B1(new_n302), .B2(new_n308), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n298), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n187), .A3(new_n309), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT90), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n272), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n272), .B1(new_n317), .B2(new_n318), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n211), .A2(G952), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(G234), .B2(G237), .ZN(new_n325));
  AOI211_X1 g139(.A(new_n187), .B(new_n211), .C1(G234), .C2(G237), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT21), .B(G898), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n267), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G214), .B1(G237), .B2(G902), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n234), .A2(G107), .ZN(new_n331));
  INV_X1    g145(.A(G101), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n234), .A2(G107), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT3), .B1(new_n335), .B2(KEYINPUT77), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n282), .A2(KEYINPUT77), .A3(KEYINPUT3), .A4(G104), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n334), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n282), .A2(G104), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n332), .B1(new_n340), .B2(new_n331), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(KEYINPUT78), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n282), .A2(KEYINPUT77), .A3(G104), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n333), .B1(new_n347), .B2(new_n337), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n344), .B1(new_n348), .B2(new_n341), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G113), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n275), .A2(G119), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT5), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT66), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n275), .B2(G119), .ZN(new_n356));
  INV_X1    g170(.A(G119), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT66), .A3(G116), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n275), .A2(G119), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n354), .B1(new_n360), .B2(new_n353), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n351), .A2(KEYINPUT2), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT2), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G113), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n365), .A2(new_n356), .A3(new_n358), .A4(new_n359), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n350), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n282), .A2(G104), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(new_n347), .B2(new_n337), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n339), .B(KEYINPUT4), .C1(new_n371), .C2(new_n332), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n362), .A2(new_n364), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n360), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n366), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT67), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n331), .B1(new_n336), .B2(new_n338), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G101), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n374), .A2(new_n366), .A3(KEYINPUT67), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n372), .A2(new_n377), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n369), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G110), .B(G122), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n369), .A2(new_n382), .A3(new_n384), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(KEYINPUT6), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT6), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n383), .A2(new_n389), .A3(new_n385), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n203), .A2(G143), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n222), .B2(G146), .ZN(new_n393));
  INV_X1    g207(.A(G128), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(KEYINPUT1), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n203), .B1(new_n220), .B2(new_n221), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n203), .A2(G143), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(KEYINPUT65), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT65), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G128), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n391), .A2(KEYINPUT1), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n393), .A2(new_n395), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n195), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n289), .A2(G146), .A3(new_n290), .ZN(new_n408));
  AND2_X1   g222(.A1(KEYINPUT0), .A2(G128), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n391), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n397), .B1(new_n213), .B2(new_n203), .ZN(new_n411));
  NOR2_X1   g225(.A1(KEYINPUT0), .A2(G128), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n410), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G125), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n407), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G224), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(G953), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n417), .B(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n388), .A2(new_n390), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n384), .B(KEYINPUT8), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n348), .A2(new_n341), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n368), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n367), .B1(new_n343), .B2(new_n349), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(KEYINPUT82), .A2(KEYINPUT7), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n407), .A2(new_n416), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT7), .B1(new_n418), .B2(G953), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n429), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n407), .A2(new_n416), .A3(new_n431), .A4(new_n427), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n387), .A2(new_n426), .A3(new_n430), .A4(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n433), .A2(new_n187), .ZN(new_n434));
  OAI21_X1  g248(.A(G210), .B1(G237), .B2(G902), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n421), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n435), .B1(new_n421), .B2(new_n434), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n330), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(KEYINPUT83), .B(new_n330), .C1(new_n436), .C2(new_n437), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n329), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT28), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n377), .A2(new_n381), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n288), .B2(G137), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n288), .A2(G137), .ZN(new_n447));
  INV_X1    g261(.A(G137), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT11), .A3(G134), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G131), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n446), .A2(new_n449), .A3(new_n209), .A4(new_n447), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n399), .A2(new_n413), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n410), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n448), .A2(G134), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n288), .A2(G137), .ZN(new_n457));
  OAI21_X1  g271(.A(G131), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n408), .A2(new_n391), .A3(new_n395), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n396), .A2(new_n398), .B1(new_n403), .B2(new_n404), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n444), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n393), .A2(new_n409), .B1(new_n399), .B2(new_n413), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT1), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n467), .B1(G143), .B2(new_n203), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n286), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n460), .B1(new_n411), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n466), .A2(new_n453), .B1(new_n470), .B2(new_n459), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n377), .A2(new_n381), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n443), .B1(new_n465), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n210), .A2(new_n211), .A3(G210), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT26), .B(G101), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT28), .B1(new_n471), .B2(new_n472), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n474), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(G902), .B1(new_n481), .B2(KEYINPUT29), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n444), .A2(new_n464), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n471), .A2(new_n472), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT28), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n479), .ZN(new_n486));
  INV_X1    g300(.A(new_n480), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT68), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n451), .A2(new_n452), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(new_n415), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n452), .A2(new_n458), .ZN(new_n492));
  AOI21_X1  g306(.A(G146), .B1(new_n289), .B2(new_n290), .ZN(new_n493));
  OAI22_X1  g307(.A1(new_n493), .A2(new_n397), .B1(new_n468), .B2(new_n286), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n494), .B2(new_n460), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n489), .B(KEYINPUT30), .C1(new_n491), .C2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT68), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n489), .A2(KEYINPUT30), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n455), .A2(new_n463), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n472), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n479), .B1(new_n501), .B2(new_n483), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT29), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n488), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n482), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT71), .B1(new_n505), .B2(G472), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT71), .ZN(new_n507));
  INV_X1    g321(.A(G472), .ZN(new_n508));
  AOI211_X1 g322(.A(new_n507), .B(new_n508), .C1(new_n482), .C2(new_n504), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  AOI211_X1 g324(.A(KEYINPUT68), .B(new_n497), .C1(new_n455), .C2(new_n463), .ZN(new_n511));
  AND4_X1   g325(.A1(new_n463), .A2(new_n455), .A3(new_n498), .A4(new_n499), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n444), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT31), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n486), .A4(new_n473), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n479), .B1(new_n474), .B2(new_n480), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n496), .A2(new_n500), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n483), .B1(new_n518), .B2(new_n444), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n514), .B1(new_n519), .B2(new_n486), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n508), .B(new_n187), .C1(new_n517), .C2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT32), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(KEYINPUT70), .A3(new_n522), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n513), .A2(new_n486), .A3(new_n473), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT31), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n516), .A3(new_n515), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n529), .A2(KEYINPUT32), .A3(new_n508), .A4(new_n187), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n510), .A2(new_n525), .A3(new_n526), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n297), .B1(G234), .B2(new_n187), .ZN(new_n532));
  INV_X1    g346(.A(G110), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n286), .A2(KEYINPUT23), .A3(G119), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n357), .A2(G128), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT23), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT73), .B1(new_n357), .B2(G128), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT73), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(new_n394), .A3(G119), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n533), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n400), .A2(new_n402), .A3(G119), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT72), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n542), .A2(new_n543), .A3(new_n535), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n543), .B1(new_n542), .B2(new_n535), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT24), .B(G110), .Z(new_n547));
  AOI21_X1  g361(.A(new_n541), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n206), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n542), .A2(new_n535), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT72), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n542), .A2(new_n543), .A3(new_n535), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n534), .A2(new_n540), .A3(new_n533), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n205), .B(new_n238), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT22), .B(G137), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n211), .A2(G221), .A3(G234), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n549), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n549), .B2(new_n555), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT25), .B1(new_n561), .B2(new_n187), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT25), .ZN(new_n563));
  NOR4_X1   g377(.A1(new_n559), .A2(new_n560), .A3(new_n563), .A4(G902), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n532), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n532), .A2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(G221), .B1(new_n296), .B2(G902), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G140), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n211), .A2(G227), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n572), .B(new_n573), .Z(new_n574));
  AOI21_X1  g388(.A(new_n394), .B1(new_n396), .B2(KEYINPUT1), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n460), .B1(new_n575), .B2(new_n393), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n423), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n372), .A2(new_n380), .A3(new_n466), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n494), .B2(new_n460), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT79), .B1(new_n350), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT78), .B1(new_n339), .B2(new_n342), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n348), .A2(new_n344), .A3(new_n341), .ZN(new_n585));
  OAI211_X1 g399(.A(KEYINPUT79), .B(new_n582), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n581), .B(new_n490), .C1(new_n583), .C2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n343), .A2(new_n406), .A3(new_n349), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT80), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n343), .A2(new_n406), .A3(KEYINPUT80), .A4(new_n349), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n577), .A3(new_n592), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n593), .A2(KEYINPUT12), .A3(new_n453), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT12), .B1(new_n593), .B2(new_n453), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n588), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n587), .A2(new_n583), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n579), .A2(new_n580), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT81), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT81), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n581), .B(new_n600), .C1(new_n583), .C2(new_n587), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n601), .A3(new_n453), .ZN(new_n602));
  INV_X1    g416(.A(new_n583), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n598), .B1(new_n603), .B2(new_n586), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n574), .B1(new_n604), .B2(new_n490), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n574), .A2(new_n596), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G469), .B1(new_n606), .B2(G902), .ZN(new_n607));
  INV_X1    g421(.A(G469), .ZN(new_n608));
  INV_X1    g422(.A(new_n574), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n602), .B2(new_n588), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n594), .A2(new_n595), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n588), .A2(new_n609), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n608), .B(new_n187), .C1(new_n610), .C2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n571), .B1(new_n607), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n442), .A2(new_n531), .A3(new_n569), .A4(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT91), .B(G101), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G3));
  OAI21_X1  g432(.A(new_n187), .B1(new_n517), .B2(new_n520), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT92), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT92), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n529), .A2(new_n621), .A3(new_n187), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n620), .A2(new_n622), .A3(KEYINPUT93), .A4(G472), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n620), .A2(G472), .A3(new_n622), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT93), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n521), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n623), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n568), .B(new_n571), .C1(new_n607), .C2(new_n614), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n317), .A2(new_n268), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT94), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n313), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n316), .A2(new_n632), .A3(new_n309), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT94), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT95), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n299), .B1(new_n315), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n315), .A2(new_n636), .A3(new_n299), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT33), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n633), .B(new_n635), .C1(new_n637), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n187), .A2(G478), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n630), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n267), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n643), .A2(new_n438), .A3(new_n328), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n629), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT96), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT34), .B(G104), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  XNOR2_X1  g462(.A(new_n317), .B(new_n318), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n321), .B1(new_n649), .B2(new_n272), .ZN(new_n650));
  NOR4_X1   g464(.A1(new_n438), .A2(new_n267), .A3(new_n650), .A4(new_n328), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n629), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT97), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NAND2_X1  g469(.A1(new_n549), .A2(new_n555), .ZN(new_n656));
  INV_X1    g470(.A(new_n558), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(KEYINPUT36), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n566), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n565), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n442), .A2(new_n627), .A3(new_n615), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT98), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  AOI21_X1  g479(.A(new_n235), .B1(new_n258), .B2(new_n242), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n230), .A2(new_n231), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n207), .A2(new_n206), .B1(new_n227), .B2(new_n228), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n667), .A2(new_n668), .B1(new_n239), .B2(new_n241), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n666), .B1(new_n669), .B2(new_n235), .ZN(new_n670));
  OAI21_X1  g484(.A(KEYINPUT20), .B1(new_n670), .B2(new_n265), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n262), .A2(new_n247), .A3(new_n263), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n325), .ZN(new_n674));
  INV_X1    g488(.A(new_n326), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n674), .B1(G900), .B2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n323), .A2(new_n673), .A3(new_n246), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT99), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n671), .A2(new_n672), .B1(G475), .B2(new_n245), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n680), .A3(new_n323), .A4(new_n676), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n330), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n421), .A2(new_n434), .ZN(new_n684));
  INV_X1    g498(.A(new_n435), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n421), .A2(new_n434), .A3(new_n435), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n683), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n688), .A2(new_n661), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n682), .A2(new_n531), .A3(new_n615), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XNOR2_X1  g505(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n676), .B(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n615), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT104), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n486), .B1(new_n465), .B2(new_n473), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n508), .B1(new_n699), .B2(KEYINPUT100), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n700), .B(new_n527), .C1(KEYINPUT100), .C2(new_n699), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n702));
  NAND2_X1  g516(.A1(G472), .A2(G902), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n701), .B2(new_n703), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n525), .A2(new_n706), .A3(new_n526), .A4(new_n530), .ZN(new_n707));
  NOR4_X1   g521(.A1(new_n679), .A2(new_n661), .A3(new_n650), .A4(new_n683), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n436), .A2(new_n437), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT38), .Z(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n708), .A2(new_n709), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n710), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n697), .A2(new_n698), .A3(new_n707), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n213), .ZN(G45));
  AND3_X1   g531(.A1(new_n642), .A2(new_n267), .A3(new_n676), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n531), .A2(new_n615), .A3(new_n689), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  AND3_X1   g534(.A1(new_n488), .A2(new_n502), .A3(new_n503), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n187), .B1(new_n488), .B2(new_n503), .ZN(new_n722));
  OAI21_X1  g536(.A(G472), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n507), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n505), .A2(KEYINPUT71), .A3(G472), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n724), .A2(new_n530), .A3(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n521), .A2(KEYINPUT70), .A3(new_n522), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT70), .B1(new_n521), .B2(new_n522), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n568), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n187), .B1(new_n610), .B2(new_n613), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G469), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n732), .A2(new_n570), .A3(new_n614), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n644), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND4_X1  g550(.A1(new_n531), .A2(new_n733), .A3(new_n569), .A4(new_n651), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  NAND4_X1  g552(.A1(new_n531), .A2(new_n733), .A3(new_n329), .A4(new_n689), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n619), .A2(G472), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n521), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(new_n743), .B2(new_n568), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n569), .A2(new_n742), .A3(KEYINPUT105), .A4(new_n521), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n732), .A2(new_n570), .A3(new_n614), .A4(new_n688), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT106), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n679), .B2(new_n650), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n267), .A2(KEYINPUT106), .A3(new_n323), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n328), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n746), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  INV_X1    g568(.A(new_n743), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n718), .A2(new_n755), .A3(new_n661), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n748), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G125), .ZN(G27));
  NOR3_X1   g573(.A1(new_n436), .A2(new_n437), .A3(new_n683), .ZN(new_n760));
  INV_X1    g574(.A(new_n614), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n596), .A2(new_n574), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n602), .A2(new_n605), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n608), .B1(new_n764), .B2(new_n187), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n570), .B(new_n760), .C1(new_n761), .C2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT107), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n615), .A2(KEYINPUT107), .A3(new_n760), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT42), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n718), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n730), .A2(new_n768), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n615), .A2(KEYINPUT107), .A3(new_n760), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT107), .B1(new_n615), .B2(new_n760), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n724), .A2(new_n530), .A3(new_n725), .A4(new_n523), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n569), .A3(new_n718), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n772), .B1(new_n777), .B2(new_n770), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n209), .ZN(G33));
  NAND4_X1  g593(.A1(new_n730), .A2(new_n768), .A3(new_n682), .A4(new_n769), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n608), .B1(new_n764), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n782), .B2(new_n764), .ZN(new_n784));
  NAND2_X1  g598(.A1(G469), .A2(G902), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT46), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(new_n761), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n785), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n570), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n693), .ZN(new_n790));
  INV_X1    g604(.A(new_n760), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT108), .B1(new_n679), .B2(new_n642), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT43), .Z(new_n793));
  INV_X1    g607(.A(new_n627), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n793), .A2(new_n794), .A3(new_n661), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n791), .B1(new_n795), .B2(KEYINPUT44), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n790), .B(new_n796), .C1(KEYINPUT44), .C2(new_n795), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  XNOR2_X1  g612(.A(new_n789), .B(KEYINPUT47), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n718), .A2(new_n568), .A3(new_n760), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n799), .A2(new_n531), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n189), .ZN(G42));
  AND2_X1   g616(.A1(new_n732), .A2(new_n614), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT110), .Z(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n805), .A2(KEYINPUT49), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(KEYINPUT49), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n679), .A2(new_n642), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n808), .A2(new_n568), .A3(new_n571), .A4(new_n683), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(KEYINPUT109), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(KEYINPUT109), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n810), .A2(new_n811), .A3(new_n707), .A4(new_n712), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n806), .A2(new_n807), .A3(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n793), .A2(new_n325), .A3(new_n746), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n760), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n804), .A2(new_n571), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n815), .B1(new_n799), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n793), .A2(new_n325), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n755), .A2(new_n661), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n733), .A2(new_n760), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n707), .A2(new_n568), .A3(new_n674), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  OR3_X1    g641(.A1(new_n827), .A2(new_n267), .A3(new_n642), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n814), .A2(new_n683), .A3(new_n713), .A4(new_n733), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT50), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n818), .A2(new_n829), .A3(new_n830), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n825), .A3(new_n828), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT51), .B1(new_n835), .B2(new_n817), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n775), .A2(new_n569), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n819), .A2(new_n837), .A3(new_n822), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT48), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n827), .A2(new_n643), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n324), .B(new_n840), .C1(new_n748), .C2(new_n814), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(KEYINPUT119), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n834), .A2(new_n836), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n525), .A2(new_n526), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n724), .A2(new_n530), .A3(new_n725), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n689), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n615), .A2(new_n678), .A3(new_n681), .ZN(new_n849));
  OAI22_X1  g663(.A1(new_n848), .A2(new_n849), .B1(new_n747), .B2(new_n756), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n615), .A2(new_n718), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n438), .B1(new_n750), .B2(new_n751), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n565), .A2(new_n660), .A3(new_n676), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT112), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n565), .A2(new_n857), .A3(new_n660), .A4(new_n676), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n854), .A2(new_n707), .A3(new_n615), .A4(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n859), .A2(new_n615), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(KEYINPUT113), .A3(new_n707), .A4(new_n854), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n853), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT52), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT52), .B1(new_n848), .B2(new_n851), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n850), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n870), .A2(KEYINPUT114), .A3(new_n865), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT114), .B1(new_n870), .B2(new_n865), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n768), .A2(new_n757), .A3(new_n769), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n679), .A2(new_n661), .A3(new_n650), .A4(new_n676), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n531), .A2(new_n615), .A3(new_n760), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n780), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n440), .A2(new_n441), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n679), .A2(new_n323), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n328), .B1(new_n643), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n627), .A2(new_n628), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n662), .A2(new_n616), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT111), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT111), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n662), .A2(new_n616), .A3(new_n882), .A4(new_n885), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n874), .B(new_n878), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n734), .A2(new_n753), .A3(new_n737), .A4(new_n739), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT117), .B1(new_n778), .B2(new_n888), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n734), .A2(new_n753), .A3(new_n737), .A4(new_n739), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n768), .A2(new_n769), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT42), .B1(new_n892), .B2(new_n776), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n890), .A2(new_n891), .A3(new_n893), .A4(new_n772), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n873), .A2(new_n887), .A3(new_n889), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  XOR2_X1   g710(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n897));
  NOR2_X1   g711(.A1(new_n778), .A2(new_n888), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n884), .A2(new_n886), .ZN(new_n899));
  INV_X1    g713(.A(new_n878), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n866), .A2(new_n867), .B1(new_n865), .B2(new_n870), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n895), .A2(new_n896), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT52), .B1(new_n853), .B2(new_n865), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT114), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n862), .A2(new_n864), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n690), .A2(new_n758), .A3(KEYINPUT52), .A4(new_n719), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n870), .A2(new_n865), .A3(KEYINPUT114), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n874), .B1(new_n911), .B2(new_n901), .ZN(new_n912));
  INV_X1    g726(.A(new_n902), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n878), .B1(new_n884), .B2(new_n886), .ZN(new_n914));
  INV_X1    g728(.A(new_n897), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n913), .A2(new_n898), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n896), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT116), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n904), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n845), .B(KEYINPUT120), .C1(new_n919), .C2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(G952), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n211), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n912), .A2(new_n916), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT54), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n895), .A2(new_n896), .A3(new_n903), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(KEYINPUT116), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n920), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT120), .B1(new_n930), .B2(new_n845), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n813), .B1(new_n925), .B2(new_n931), .ZN(G75));
  NOR2_X1   g746(.A1(new_n211), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AND4_X1   g748(.A1(KEYINPUT53), .A2(new_n914), .A3(new_n894), .A4(new_n889), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n907), .A2(new_n908), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n914), .B(new_n898), .C1(new_n905), .C2(new_n936), .ZN(new_n937));
  AOI22_X1  g751(.A1(new_n935), .A2(new_n873), .B1(new_n937), .B2(new_n897), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n187), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT56), .B1(new_n939), .B2(G210), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n388), .A2(new_n390), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n420), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n934), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n940), .B2(new_n943), .ZN(G51));
  NAND2_X1  g759(.A1(new_n895), .A2(new_n903), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT54), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n928), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n785), .B(KEYINPUT57), .Z(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT121), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n610), .A2(new_n613), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n948), .A2(new_n953), .A3(new_n949), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  OR3_X1    g769(.A1(new_n938), .A2(new_n187), .A3(new_n784), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n933), .B1(new_n955), .B2(new_n956), .ZN(G54));
  NAND3_X1  g771(.A1(new_n939), .A2(KEYINPUT58), .A3(G475), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n958), .A2(new_n670), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n670), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n933), .ZN(G60));
  XOR2_X1   g775(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n962));
  NOR2_X1   g776(.A1(new_n268), .A2(new_n187), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n640), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n948), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n934), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n930), .A2(new_n964), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n640), .ZN(G63));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n970));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n970), .B1(new_n946), .B2(new_n973), .ZN(new_n974));
  AOI211_X1 g788(.A(KEYINPUT123), .B(new_n972), .C1(new_n895), .C2(new_n903), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n561), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n933), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n659), .B1(new_n974), .B2(new_n975), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n978), .B(new_n979), .C1(KEYINPUT124), .C2(KEYINPUT61), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT123), .B1(new_n938), .B2(new_n972), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n946), .A2(new_n970), .A3(new_n973), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n977), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n979), .A2(new_n983), .A3(new_n934), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n983), .A2(KEYINPUT124), .A3(new_n934), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n980), .A2(new_n987), .ZN(G66));
  OAI21_X1  g802(.A(G953), .B1(new_n327), .B2(new_n418), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n899), .A2(new_n890), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT125), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n989), .B1(new_n991), .B2(G953), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n941), .B1(G898), .B2(new_n211), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(G69));
  XNOR2_X1  g808(.A(new_n518), .B(new_n256), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n790), .A2(new_n837), .A3(new_n854), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n997), .A2(new_n893), .A3(new_n772), .A4(new_n780), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n801), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT127), .B1(new_n797), .B2(new_n853), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n797), .A2(KEYINPUT127), .A3(new_n853), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n999), .B(new_n211), .C1(new_n1000), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G900), .A2(G953), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n996), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n643), .A2(new_n880), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1006), .A2(KEYINPUT126), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1007), .A2(new_n791), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(KEYINPUT126), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1008), .A2(new_n730), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n797), .B1(new_n696), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT62), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n716), .A2(new_n1012), .A3(new_n853), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n716), .B2(new_n853), .ZN(new_n1014));
  NOR4_X1   g828(.A1(new_n801), .A2(new_n1011), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NOR3_X1   g829(.A1(new_n1015), .A2(G953), .A3(new_n995), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n211), .B1(G227), .B2(G900), .ZN(new_n1017));
  NOR3_X1   g831(.A1(new_n1005), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1019));
  NAND2_X1  g833(.A1(G227), .A2(G900), .ZN(new_n1020));
  AND4_X1   g834(.A1(G953), .A2(new_n1019), .A3(new_n1020), .A4(new_n995), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1018), .A2(new_n1021), .ZN(G72));
  XNOR2_X1  g836(.A(new_n703), .B(KEYINPUT63), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1002), .A2(new_n1000), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1024), .A2(new_n801), .A3(new_n998), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1023), .B1(new_n1025), .B2(new_n991), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n519), .A2(new_n479), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1023), .B1(new_n1015), .B2(new_n991), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n486), .B1(new_n501), .B2(new_n483), .ZN(new_n1029));
  OAI22_X1  g843(.A1(new_n1026), .A2(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1023), .B1(new_n502), .B2(new_n527), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n926), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(new_n934), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1030), .A2(new_n1033), .ZN(G57));
endmodule


