//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n446, new_n448, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n544,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G452), .ZN(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G137), .ZN(new_n461));
  INV_X1    g036(.A(G101), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n459), .A2(G2104), .ZN(new_n463));
  OAI22_X1  g038(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n458), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(new_n467), .ZN(G160));
  NAND2_X1  g043(.A1(new_n458), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G124), .ZN(new_n470));
  NOR2_X1   g045(.A1(G100), .A2(G2105), .ZN(new_n471));
  OAI21_X1  g046(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n472));
  OAI22_X1  g047(.A1(new_n469), .A2(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n460), .B(KEYINPUT69), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G136), .ZN(G162));
  OAI21_X1  g050(.A(G2104), .B1(new_n459), .B2(G114), .ZN(new_n476));
  NOR2_X1   g051(.A1(G102), .A2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(G126), .A2(G2105), .ZN(new_n479));
  AND2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g059(.A(KEYINPUT70), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n478), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G138), .B(new_n459), .C1(new_n480), .C2(new_n481), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n458), .A2(new_n489), .A3(G138), .A4(new_n459), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  INV_X1    g068(.A(G651), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT6), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT6), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G651), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT72), .B(G88), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n495), .A2(new_n497), .A3(G50), .A4(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n500), .A2(new_n502), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n506), .A2(new_n509), .A3(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n498), .A2(new_n503), .ZN(new_n519));
  INV_X1    g094(.A(G89), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n498), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(G51), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n519), .A2(new_n531), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n494), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G171));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n519), .A2(new_n537), .B1(new_n525), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n494), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT74), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G188));
  NAND3_X1  g124(.A1(new_n498), .A2(G53), .A3(G543), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT9), .ZN(new_n551));
  NAND2_X1  g126(.A1(G78), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G65), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n511), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n504), .A2(G91), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n551), .A2(new_n555), .A3(new_n556), .ZN(G299));
  INV_X1    g132(.A(G171), .ZN(G301));
  NAND2_X1  g133(.A1(new_n526), .A2(G49), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n504), .A2(G87), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(G288));
  INV_X1    g137(.A(G61), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n511), .A2(KEYINPUT75), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G73), .A2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT75), .B1(new_n511), .B2(new_n563), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  INV_X1    g143(.A(G86), .ZN(new_n569));
  INV_X1    g144(.A(G48), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n519), .A2(new_n569), .B1(new_n525), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G305));
  INV_X1    g148(.A(G85), .ZN(new_n574));
  INV_X1    g149(.A(G47), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n519), .A2(new_n574), .B1(new_n525), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n494), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n504), .A2(KEYINPUT10), .A3(G92), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT10), .ZN(new_n583));
  INV_X1    g158(.A(G92), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n519), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n526), .A2(G54), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  XOR2_X1   g163(.A(KEYINPUT76), .B(G66), .Z(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n511), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n581), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n581), .B1(new_n593), .B2(G868), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT9), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n550), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n556), .A2(new_n555), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n596), .B1(G868), .B2(new_n600), .ZN(G280));
  XNOR2_X1  g176(.A(G280), .B(KEYINPUT77), .ZN(G297));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n593), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n593), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g183(.A(new_n469), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G123), .ZN(new_n610));
  NOR2_X1   g185(.A1(G99), .A2(G2105), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(new_n459), .B2(G111), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(G135), .B2(new_n474), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT79), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2096), .Z(new_n616));
  NOR2_X1   g191(.A1(new_n480), .A2(new_n481), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n617), .A2(new_n463), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n616), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2451), .B(G2454), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2443), .B(G2446), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n627), .B(new_n628), .Z(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2435), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2438), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n629), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G14), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G401));
  XOR2_X1   g212(.A(G2084), .B(G2090), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2067), .B(G2678), .Z(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(new_n642), .A3(KEYINPUT17), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT18), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n641), .B2(KEYINPUT18), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2096), .B(G2100), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(G227));
  XNOR2_X1  g225(.A(G1971), .B(G1976), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1956), .B(G2474), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1961), .B(G1966), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(KEYINPUT80), .B1(new_n654), .B2(new_n655), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n653), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT81), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n654), .A2(new_n655), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n653), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT82), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n661), .A2(new_n662), .ZN(new_n667));
  OR3_X1    g242(.A1(new_n653), .A2(new_n664), .A3(new_n656), .ZN(new_n668));
  NAND4_X1  g243(.A1(new_n663), .A2(new_n666), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G229));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G23), .ZN(new_n678));
  INV_X1    g253(.A(G288), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT33), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G1976), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n677), .A2(G6), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n571), .B1(G651), .B2(new_n567), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n677), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT32), .B(G1981), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n677), .A2(G22), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G166), .B2(new_n677), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(G1971), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n685), .A2(new_n686), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(G1971), .ZN(new_n692));
  AND3_X1   g267(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n682), .A2(new_n687), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(KEYINPUT34), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT83), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n579), .A2(new_n677), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n677), .B2(G24), .ZN(new_n698));
  INV_X1    g273(.A(G1986), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n694), .A2(KEYINPUT34), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G25), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n474), .A2(G131), .ZN(new_n704));
  INV_X1    g279(.A(G119), .ZN(new_n705));
  NOR2_X1   g280(.A1(G95), .A2(G2105), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(new_n459), .B2(G107), .ZN(new_n707));
  OAI22_X1  g282(.A1(new_n469), .A2(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n703), .B1(new_n709), .B2(new_n702), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT35), .B(G1991), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n699), .B2(new_n698), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n701), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n696), .A2(new_n700), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT36), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n615), .A2(new_n702), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n702), .A2(G33), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n458), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(new_n459), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n474), .B2(G139), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT25), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n719), .B1(new_n727), .B2(new_n702), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n542), .A2(new_n677), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n677), .B2(G19), .ZN(new_n730));
  INV_X1    g305(.A(G1341), .ZN(new_n731));
  OAI22_X1  g306(.A1(new_n728), .A2(G2072), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n718), .B(new_n732), .C1(G2072), .C2(new_n728), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT31), .B(G11), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n730), .A2(new_n731), .ZN(new_n735));
  NOR2_X1   g310(.A1(G5), .A2(G16), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G171), .B2(G16), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G1961), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G28), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(G28), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n740), .A2(new_n741), .A3(new_n702), .ZN(new_n742));
  INV_X1    g317(.A(G2084), .ZN(new_n743));
  AND2_X1   g318(.A1(KEYINPUT24), .A2(G34), .ZN(new_n744));
  NOR2_X1   g319(.A1(KEYINPUT24), .A2(G34), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n744), .A2(new_n745), .A3(G29), .ZN(new_n746));
  INV_X1    g321(.A(G160), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(G29), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n738), .B(new_n742), .C1(new_n743), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n677), .A2(G21), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G168), .B2(new_n677), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n749), .B1(new_n751), .B2(G1966), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n733), .A2(new_n734), .A3(new_n735), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n702), .A2(G27), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G164), .B2(new_n702), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT89), .B(G2078), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n677), .A2(G4), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n593), .B2(new_n677), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1348), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n702), .A2(G26), .ZN(new_n761));
  INV_X1    g336(.A(G128), .ZN(new_n762));
  NOR2_X1   g337(.A1(G104), .A2(G2105), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(new_n459), .B2(G116), .ZN(new_n764));
  OAI22_X1  g339(.A1(new_n469), .A2(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n474), .B2(G140), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n761), .B1(new_n767), .B2(G29), .ZN(new_n768));
  MUX2_X1   g343(.A(new_n761), .B(new_n768), .S(KEYINPUT28), .Z(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n753), .A2(new_n757), .A3(new_n760), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n702), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n702), .ZN(new_n774));
  MUX2_X1   g349(.A(new_n773), .B(new_n774), .S(KEYINPUT90), .Z(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT29), .Z(new_n776));
  INV_X1    g351(.A(G2090), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n772), .B(new_n778), .C1(G1966), .C2(new_n751), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT85), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT86), .B(KEYINPUT26), .ZN(new_n782));
  AND3_X1   g357(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G129), .B2(new_n609), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n474), .A2(KEYINPUT84), .A3(G141), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(KEYINPUT84), .B1(new_n474), .B2(G141), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n781), .B(new_n787), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(KEYINPUT87), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT87), .ZN(new_n793));
  INV_X1    g368(.A(new_n787), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n474), .A2(G141), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT84), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n794), .B1(new_n797), .B2(new_n788), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n793), .B1(new_n798), .B2(new_n781), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n792), .A2(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G32), .B(new_n800), .S(G29), .Z(new_n801));
  XOR2_X1   g376(.A(KEYINPUT27), .B(G1996), .Z(new_n802));
  AOI22_X1  g377(.A1(new_n801), .A2(new_n802), .B1(new_n743), .B2(new_n748), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G1961), .B2(new_n737), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT88), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n776), .A2(new_n777), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT91), .Z(new_n807));
  NOR2_X1   g382(.A1(new_n801), .A2(new_n802), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n779), .A2(new_n805), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n677), .A2(G20), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n600), .B2(new_n677), .ZN(new_n811));
  MUX2_X1   g386(.A(new_n810), .B(new_n811), .S(KEYINPUT23), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT92), .B(G1956), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n717), .A2(new_n809), .A3(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  NAND2_X1  g391(.A1(new_n593), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  INV_X1    g393(.A(G93), .ZN(new_n819));
  INV_X1    g394(.A(G55), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n519), .A2(new_n819), .B1(new_n525), .B2(new_n820), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n494), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(new_n542), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n539), .A2(new_n541), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n821), .A2(new_n823), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT39), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n818), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT93), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n824), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT37), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(G145));
  INV_X1    g411(.A(G37), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n766), .B(new_n492), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n727), .B1(new_n792), .B2(new_n799), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n791), .A2(new_n726), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n791), .A2(KEYINPUT87), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n798), .A2(new_n793), .A3(new_n781), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n726), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n841), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n845), .A2(new_n838), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n850), .B(new_n851), .C1(G118), .C2(new_n459), .ZN(new_n852));
  INV_X1    g427(.A(G130), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(new_n469), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n474), .B2(G142), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n619), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n709), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n842), .A2(new_n847), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(G160), .B(KEYINPUT94), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(G162), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(new_n615), .Z(new_n863));
  NAND3_X1  g438(.A1(new_n840), .A2(new_n839), .A3(new_n841), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n838), .B1(new_n845), .B2(new_n846), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(new_n865), .A3(new_n857), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n860), .B(new_n863), .C1(new_n859), .C2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n858), .B1(new_n842), .B2(new_n847), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n863), .B1(new_n868), .B2(new_n866), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n869), .A2(KEYINPUT96), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n871));
  AOI211_X1 g446(.A(new_n871), .B(new_n863), .C1(new_n868), .C2(new_n866), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n837), .B(new_n867), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT98), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g450(.A(new_n679), .B(new_n684), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n579), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(G290), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n878), .A2(G166), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(G166), .B1(new_n878), .B2(new_n879), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT42), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n605), .B(new_n829), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n586), .A2(new_n591), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT99), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n885), .A2(new_n886), .A3(G299), .A4(new_n587), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT99), .B1(new_n592), .B2(new_n600), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n592), .A2(new_n600), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n884), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n887), .A2(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(KEYINPUT100), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n592), .A2(new_n600), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n892), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n889), .A2(KEYINPUT41), .A3(new_n890), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n889), .A2(new_n894), .A3(new_n896), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(KEYINPUT101), .A3(new_n892), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n891), .B1(new_n904), .B2(new_n884), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n883), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n883), .A2(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(G868), .B2(new_n827), .ZN(G295));
  XNOR2_X1  g485(.A(G295), .B(KEYINPUT102), .ZN(G331));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  AOI21_X1  g487(.A(G301), .B1(new_n825), .B2(new_n828), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n825), .A2(new_n828), .A3(G301), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(G168), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n915), .ZN(new_n917));
  OAI21_X1  g492(.A(G286), .B1(new_n917), .B2(new_n913), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n900), .A2(new_n901), .A3(new_n903), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n889), .A2(new_n890), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n882), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n923), .A2(G37), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n892), .B1(new_n916), .B2(new_n918), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n902), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n882), .B(new_n926), .C1(new_n921), .C2(new_n925), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n912), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n928), .B(KEYINPUT106), .Z(new_n929));
  AND3_X1   g504(.A1(new_n920), .A2(new_n922), .A3(new_n882), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n930), .A2(new_n923), .A3(G37), .ZN(new_n931));
  XOR2_X1   g506(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n929), .A2(KEYINPUT44), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n931), .B2(new_n933), .ZN(new_n937));
  INV_X1    g512(.A(new_n923), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n920), .A2(new_n922), .A3(new_n882), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n837), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(KEYINPUT104), .A3(new_n932), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n938), .A2(new_n837), .A3(new_n933), .A4(new_n927), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n924), .A2(KEYINPUT105), .A3(new_n933), .A4(new_n927), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n937), .A2(new_n941), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n935), .B1(KEYINPUT44), .B2(new_n946), .ZN(G397));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n492), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n952));
  AOI21_X1  g527(.A(G1384), .B1(new_n486), .B2(new_n491), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT107), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G2078), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n465), .A2(new_n466), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(G2105), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n463), .A2(new_n462), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n617), .A2(G2105), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n960), .B2(G137), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n961), .A3(G40), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n953), .B2(KEYINPUT45), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n955), .A2(KEYINPUT53), .A3(new_n956), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n949), .A2(new_n952), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(new_n965), .A3(new_n956), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n958), .A2(G40), .A3(new_n961), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n971), .B(G1384), .C1(new_n486), .C2(new_n491), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n969), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1961), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n964), .A2(new_n968), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(G171), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n963), .A2(new_n965), .A3(KEYINPUT53), .A4(new_n956), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n975), .A2(KEYINPUT120), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT120), .B1(new_n975), .B2(new_n979), .ZN(new_n981));
  INV_X1    g556(.A(new_n968), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n978), .B1(new_n983), .B2(G301), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(KEYINPUT121), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT121), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n975), .A2(new_n979), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT120), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n975), .A2(KEYINPUT120), .A3(new_n979), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n968), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n977), .B1(new_n992), .B2(G171), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n987), .B1(new_n993), .B2(KEYINPUT54), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n995));
  INV_X1    g570(.A(G1981), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n684), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI211_X1 g574(.A(KEYINPUT112), .B(KEYINPUT49), .C1(new_n684), .C2(new_n996), .ZN(new_n1000));
  OAI211_X1 g575(.A(G1981), .B(G305), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n998), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT49), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G305), .A2(G1981), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n997), .A2(new_n998), .A3(new_n995), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n969), .A2(new_n953), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G8), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1001), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n949), .A2(new_n971), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n962), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n777), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n963), .A2(new_n965), .ZN(new_n1015));
  INV_X1    g590(.A(G1971), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G303), .A2(G8), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT111), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n1022));
  NAND4_X1  g597(.A1(G303), .A2(KEYINPUT110), .A3(new_n1022), .A4(G8), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1021), .A2(new_n1026), .A3(new_n1023), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1018), .A2(new_n1028), .A3(G8), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1008), .B1(G1976), .B2(new_n679), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1031), .B(new_n1032), .C1(G1976), .C2(new_n679), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1010), .A2(new_n1030), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1018), .A2(G8), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1037), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1035), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n986), .A2(new_n994), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n983), .A2(G301), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n976), .B(KEYINPUT122), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1043), .B(KEYINPUT54), .C1(new_n1044), .C2(G301), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G286), .A2(G8), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1966), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n492), .A2(KEYINPUT45), .A3(new_n948), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n969), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n953), .A2(KEYINPUT45), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1013), .A2(new_n743), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1015), .A2(KEYINPUT114), .A3(new_n1048), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AOI211_X1 g632(.A(KEYINPUT51), .B(new_n1047), .C1(new_n1057), .C2(G8), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(KEYINPUT118), .A3(G8), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1046), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT118), .B1(new_n1057), .B2(G8), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT51), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT119), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1064), .B(KEYINPUT51), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1058), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1057), .A2(new_n1047), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1042), .B(new_n1045), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT123), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1058), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1065), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1057), .A2(G8), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1075), .A2(new_n1046), .A3(new_n1059), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1064), .B1(new_n1076), .B2(KEYINPUT51), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1071), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n1067), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n1045), .A4(new_n1042), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1013), .A2(G1348), .B1(G2067), .B2(new_n1007), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1082), .A2(new_n593), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n600), .B(KEYINPUT115), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1084), .B(KEYINPUT57), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1015), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  INV_X1    g662(.A(G1956), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1086), .A2(new_n1087), .B1(new_n973), .B2(new_n1088), .ZN(new_n1089));
  OR3_X1    g664(.A1(new_n1085), .A2(KEYINPUT116), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT116), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1083), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1092), .A2(KEYINPUT117), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT117), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1085), .A2(new_n1089), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1996), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  AOI22_X1  g675(.A1(new_n1086), .A2(new_n1099), .B1(new_n1007), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(new_n826), .ZN(new_n1102));
  XOR2_X1   g677(.A(new_n1102), .B(KEYINPUT59), .Z(new_n1103));
  OR3_X1    g678(.A1(new_n1082), .A2(KEYINPUT60), .A3(new_n592), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1082), .A2(new_n593), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT60), .B1(new_n1083), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1098), .A2(new_n1103), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1096), .B(new_n1093), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1094), .B(new_n1095), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1070), .A2(new_n1081), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1010), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(new_n1030), .ZN(new_n1112));
  INV_X1    g687(.A(G1976), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1010), .A2(new_n1113), .A3(new_n679), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1008), .B1(new_n1114), .B2(new_n997), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1073), .A2(G286), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1041), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1111), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1118), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1120), .A2(new_n1030), .A3(new_n1116), .A4(new_n1121), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1112), .B(new_n1115), .C1(new_n1119), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1068), .B1(new_n1125), .B2(new_n1071), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1041), .A2(G171), .A3(new_n992), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1130));
  OAI211_X1 g705(.A(KEYINPUT124), .B(KEYINPUT62), .C1(new_n1066), .C2(new_n1068), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1110), .A2(new_n1123), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n955), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n969), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(G1996), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT108), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(new_n800), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n766), .B(new_n770), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(G1996), .B2(new_n791), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(new_n1135), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n709), .B(new_n711), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT109), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1135), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1144), .B2(new_n1143), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1142), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n579), .A2(new_n699), .ZN(new_n1149));
  NAND2_X1  g724(.A1(G290), .A2(G1986), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1135), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1133), .A2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n704), .A2(new_n711), .A3(new_n708), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1142), .A2(new_n1154), .B1(new_n770), .B2(new_n766), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(new_n1135), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT125), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1146), .B1(new_n791), .B2(new_n1139), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1137), .A2(KEYINPUT46), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1137), .A2(KEYINPUT46), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT47), .Z(new_n1162));
  NOR2_X1   g737(.A1(new_n1135), .A2(new_n1149), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT48), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1148), .A2(new_n1164), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1157), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1153), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n1169));
  INV_X1    g743(.A(G227), .ZN(new_n1170));
  NAND3_X1  g744(.A1(new_n636), .A2(G319), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n873), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n937), .A2(new_n941), .ZN(new_n1175));
  NAND2_X1  g749(.A1(new_n944), .A2(new_n945), .ZN(new_n1176));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g751(.A(new_n675), .B1(new_n1172), .B2(new_n1171), .ZN(new_n1178));
  INV_X1    g752(.A(new_n1178), .ZN(new_n1179));
  AOI21_X1  g753(.A(new_n1169), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  NOR4_X1   g754(.A1(new_n946), .A2(KEYINPUT127), .A3(new_n1178), .A4(new_n1174), .ZN(new_n1181));
  NOR2_X1   g755(.A1(new_n1180), .A2(new_n1181), .ZN(G308));
  NAND2_X1  g756(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1183));
  INV_X1    g757(.A(new_n1174), .ZN(new_n1184));
  NAND3_X1  g758(.A1(new_n1183), .A2(new_n1179), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n1185), .A2(KEYINPUT127), .ZN(new_n1186));
  NAND3_X1  g760(.A1(new_n1177), .A2(new_n1169), .A3(new_n1179), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1187), .ZN(G225));
endmodule


