//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1328, new_n1329, new_n1330, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n213), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n206), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n211), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n233));
  NAND4_X1  g0033(.A1(new_n217), .A2(new_n227), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n226), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n202), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n248), .B(new_n254), .ZN(G351));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT68), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(new_n201), .A3(KEYINPUT8), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n230), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n210), .A2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT16), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G159), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n276));
  AOI211_X1 g0076(.A(new_n271), .B(new_n275), .C1(new_n276), .C2(G20), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT7), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(G20), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT71), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n285));
  OAI211_X1 g0085(.A(KEYINPUT7), .B(new_n211), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n280), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n282), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n290), .A2(KEYINPUT71), .A3(KEYINPUT7), .A4(new_n211), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G68), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n277), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n263), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT72), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n280), .A2(new_n295), .A3(new_n286), .ZN(new_n296));
  OAI211_X1 g0096(.A(KEYINPUT72), .B(new_n278), .C1(new_n279), .C2(G20), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(G68), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n275), .B1(new_n276), .B2(G20), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT16), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n270), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G41), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(G1), .A3(G13), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n288), .A2(new_n289), .A3(G226), .A4(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT73), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n279), .A2(KEYINPUT73), .A3(G226), .A4(G1698), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G1698), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n288), .A2(new_n289), .A3(G223), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G87), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n303), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT67), .ZN(new_n315));
  AND2_X1   g0115(.A1(G33), .A2(G41), .ZN(new_n316));
  OAI21_X1  g0116(.A(G274), .B1(new_n316), .B2(new_n230), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n318), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n320), .A2(new_n303), .A3(KEYINPUT67), .A4(G274), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n303), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G232), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(G169), .B1(new_n314), .B2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n319), .A2(new_n321), .B1(new_n324), .B2(G232), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n312), .B1(new_n306), .B2(new_n307), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n328), .B(G179), .C1(new_n329), .C2(new_n303), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n301), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(KEYINPUT74), .A2(KEYINPUT18), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT17), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n314), .B2(new_n326), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n328), .B(new_n338), .C1(new_n329), .C2(new_n303), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n335), .B1(new_n301), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n298), .A2(new_n299), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n271), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n291), .A2(G68), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n280), .A2(new_n281), .A3(new_n286), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n264), .B1(new_n346), .B2(new_n277), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n343), .A2(new_n347), .B1(new_n269), .B2(new_n267), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n337), .A2(new_n339), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(KEYINPUT17), .A3(new_n349), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n334), .A2(new_n341), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT18), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n301), .A2(new_n352), .A3(new_n331), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n301), .B2(new_n331), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT74), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT75), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n351), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n359));
  INV_X1    g0159(.A(G150), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n211), .A2(G33), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n359), .B1(new_n360), .B2(new_n273), .C1(new_n260), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n263), .ZN(new_n363));
  MUX2_X1   g0163(.A(new_n268), .B(new_n266), .S(G50), .Z(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n322), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(G226), .B2(new_n324), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n279), .A2(G222), .A3(new_n309), .ZN(new_n368));
  INV_X1    g0168(.A(G77), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n279), .A2(G1698), .ZN(new_n370));
  INV_X1    g0170(.A(G223), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n368), .B1(new_n369), .B2(new_n279), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n323), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n365), .B1(new_n374), .B2(G169), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n367), .A2(new_n373), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(G179), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n366), .B1(G244), .B2(new_n324), .ZN(new_n379));
  INV_X1    g0179(.A(G107), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n370), .A2(new_n219), .B1(new_n380), .B2(new_n279), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n290), .A2(new_n238), .A3(G1698), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n323), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G200), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT69), .ZN(new_n386));
  INV_X1    g0186(.A(new_n268), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n263), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n268), .A2(KEYINPUT69), .A3(new_n230), .A4(new_n262), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(G77), .A3(new_n265), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G20), .A2(G77), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT15), .B(G87), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n392), .B1(new_n256), .B2(new_n273), .C1(new_n361), .C2(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n263), .B1(new_n369), .B2(new_n387), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n379), .A2(G190), .A3(new_n383), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n385), .A2(new_n391), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G169), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n384), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G179), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n379), .A2(new_n400), .A3(new_n383), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n395), .A2(new_n391), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n376), .A2(G200), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n338), .B2(new_n376), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT9), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n363), .A2(new_n407), .A3(new_n364), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n363), .B2(new_n364), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT10), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n336), .B1(new_n367), .B2(new_n373), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(G190), .B2(new_n374), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT10), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n413), .B(new_n414), .C1(new_n409), .C2(new_n408), .ZN(new_n415));
  AOI211_X1 g0215(.A(new_n378), .B(new_n404), .C1(new_n411), .C2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n288), .A2(new_n289), .A3(G232), .A4(G1698), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n288), .A2(new_n289), .A3(G226), .A4(new_n309), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G97), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n323), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n324), .A2(G238), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n322), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT13), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT70), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT13), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n421), .A2(new_n322), .A3(new_n426), .A4(new_n422), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n424), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n322), .A2(new_n422), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n429), .A2(KEYINPUT70), .A3(new_n426), .A4(new_n421), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(G200), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n390), .A2(G68), .A3(new_n265), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n211), .A2(G33), .A3(G77), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n272), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n264), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n435), .A2(KEYINPUT11), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n387), .A2(new_n202), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT12), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(KEYINPUT11), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n432), .A2(new_n436), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n338), .B1(new_n423), .B2(KEYINPUT13), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n440), .B1(new_n441), .B2(new_n427), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n428), .A2(G169), .A3(new_n430), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT14), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT14), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n428), .A2(new_n447), .A3(G169), .A4(new_n430), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n424), .A2(G179), .A3(new_n427), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n444), .B1(new_n450), .B2(new_n440), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT74), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n332), .A2(KEYINPUT18), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n452), .B1(new_n453), .B2(new_n353), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n334), .A2(new_n341), .A3(new_n350), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT75), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND4_X1   g0256(.A1(new_n358), .A2(new_n416), .A3(new_n451), .A4(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT81), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n296), .A2(G107), .A3(new_n297), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT6), .ZN(new_n461));
  AND2_X1   g0261(.A1(G97), .A2(G107), .ZN(new_n462));
  NOR2_X1   g0262(.A1(G97), .A2(G107), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n380), .A2(KEYINPUT6), .A3(G97), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n211), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n273), .A2(new_n369), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT76), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT76), .ZN(new_n469));
  INV_X1    g0269(.A(new_n467), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT6), .A2(G97), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G107), .ZN(new_n472));
  XNOR2_X1  g0272(.A(G97), .B(G107), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n461), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n469), .B(new_n470), .C1(new_n474), .C2(new_n211), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n263), .B1(new_n460), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n268), .A2(G97), .ZN(new_n478));
  AOI211_X1 g0278(.A(new_n263), .B(new_n387), .C1(new_n210), .C2(G33), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(G97), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n288), .A2(new_n289), .A3(G244), .A4(new_n309), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  AND2_X1   g0284(.A1(KEYINPUT4), .A2(G244), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n288), .A2(new_n289), .A3(new_n485), .A4(new_n309), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n288), .A2(new_n289), .A3(G250), .A4(G1698), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT77), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT77), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n279), .A2(new_n490), .A3(G250), .A4(G1698), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n323), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT79), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT5), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(G41), .ZN(new_n496));
  INV_X1    g0296(.A(G41), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G274), .ZN(new_n500));
  INV_X1    g0300(.A(new_n230), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(new_n501), .B2(new_n302), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n210), .B(G45), .C1(new_n497), .C2(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT78), .ZN(new_n504));
  INV_X1    g0304(.A(G45), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(G1), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT78), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n495), .A2(G41), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n499), .A2(new_n502), .A3(new_n504), .A4(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n496), .A2(new_n498), .A3(new_n506), .A4(new_n508), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(G257), .A3(new_n303), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n493), .A2(new_n514), .A3(G190), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n477), .A2(new_n480), .A3(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n510), .A2(KEYINPUT80), .A3(new_n512), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT80), .B1(new_n510), .B2(new_n512), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n336), .B1(new_n519), .B2(new_n493), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n459), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n480), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n296), .A2(G107), .A3(new_n297), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(new_n468), .A3(new_n475), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n522), .B1(new_n524), .B2(new_n263), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT80), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n513), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n510), .A2(KEYINPUT80), .A3(new_n512), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n493), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G200), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n525), .A2(new_n530), .A3(KEYINPUT81), .A4(new_n515), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n527), .A2(new_n493), .A3(new_n400), .A4(new_n528), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT82), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n486), .A2(new_n484), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n535), .A2(new_n483), .A3(new_n489), .A4(new_n491), .ZN(new_n536));
  AOI21_X1  g0336(.A(G179), .B1(new_n536), .B2(new_n323), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n519), .A2(KEYINPUT82), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n493), .A2(new_n514), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n477), .A2(new_n480), .B1(new_n398), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n521), .A2(new_n531), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n393), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n479), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n211), .B1(new_n419), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n463), .A2(new_n220), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n288), .A2(new_n289), .A3(new_n211), .A4(G68), .ZN(new_n549));
  INV_X1    g0349(.A(G97), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n545), .B1(new_n361), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(new_n263), .B1(new_n387), .B2(new_n393), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n544), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n288), .A2(new_n289), .A3(G238), .A4(new_n309), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G116), .ZN(new_n556));
  AND2_X1   g0356(.A1(G244), .A2(G1698), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n288), .A2(new_n289), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n323), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n221), .B1(new_n505), .B2(G1), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n210), .A2(new_n500), .A3(G45), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT83), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n303), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n303), .A2(new_n561), .A3(new_n562), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT83), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n560), .A2(new_n400), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n279), .A2(new_n557), .B1(G33), .B2(G116), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n303), .B1(new_n568), .B2(new_n555), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n564), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n398), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n554), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(G200), .B1(new_n569), .B2(new_n570), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n560), .A2(G190), .A3(new_n564), .A4(new_n566), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n210), .A2(G33), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n264), .A2(G87), .A3(new_n268), .A4(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n573), .A2(new_n574), .A3(new_n553), .A4(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n542), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n496), .A2(new_n498), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n303), .B1(new_n581), .B2(new_n503), .ZN(new_n582));
  INV_X1    g0382(.A(G270), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT84), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(G303), .B1(new_n283), .B2(new_n285), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n288), .A2(new_n289), .A3(G264), .A4(G1698), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n288), .A2(new_n289), .A3(G257), .A4(new_n309), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n323), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT84), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n511), .A2(new_n590), .A3(G270), .A4(new_n303), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n584), .A2(new_n589), .A3(new_n510), .A4(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(G116), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n210), .B2(G33), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n388), .A2(new_n389), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n387), .A2(new_n593), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n484), .B(new_n211), .C1(G33), .C2(new_n550), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT85), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT20), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n598), .A2(new_n599), .B1(new_n593), .B2(G20), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n597), .A2(new_n600), .A3(new_n263), .ZN(new_n601));
  NAND2_X1  g0401(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n595), .B(new_n596), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n592), .A2(new_n605), .A3(G169), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n592), .A2(new_n400), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n580), .A2(new_n606), .B1(new_n607), .B2(new_n605), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n592), .A2(new_n605), .A3(KEYINPUT21), .A4(G169), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT86), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n595), .A2(new_n596), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n601), .B(new_n602), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n398), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n614), .A2(KEYINPUT86), .A3(KEYINPUT21), .A4(new_n592), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n608), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n511), .A2(new_n303), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n288), .A2(new_n289), .A3(G257), .A4(G1698), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n288), .A2(new_n289), .A3(G250), .A4(new_n309), .ZN(new_n619));
  NAND2_X1  g0419(.A1(G33), .A2(G294), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n617), .A2(G264), .B1(new_n621), .B2(new_n323), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n622), .A2(new_n400), .A3(new_n510), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n323), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n511), .A2(G264), .A3(new_n303), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n510), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n398), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT23), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(new_n380), .A3(G20), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT88), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n556), .A2(new_n628), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n211), .ZN(new_n633));
  NAND2_X1  g0433(.A1(KEYINPUT23), .A2(G107), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n628), .A2(new_n380), .A3(KEYINPUT88), .A4(G20), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n631), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n288), .A2(new_n289), .A3(new_n211), .A4(G87), .ZN(new_n637));
  XNOR2_X1  g0437(.A(KEYINPUT87), .B(KEYINPUT22), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT24), .ZN(new_n641));
  NOR2_X1   g0441(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(new_n642), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(new_n279), .A3(new_n211), .A4(G87), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n629), .A2(new_n630), .B1(KEYINPUT23), .B2(G107), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n211), .A2(KEYINPUT23), .A3(G107), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n649), .A2(KEYINPUT88), .B1(new_n632), .B2(new_n211), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n647), .A2(new_n643), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT24), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n264), .B1(new_n644), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT25), .ZN(new_n654));
  AOI211_X1 g0454(.A(G107), .B(new_n268), .C1(KEYINPUT89), .C2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(KEYINPUT89), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n479), .A2(G107), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n623), .B(new_n627), .C1(new_n653), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n626), .A2(new_n336), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n624), .A2(new_n338), .A3(new_n510), .A4(new_n625), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n641), .B1(new_n640), .B2(new_n643), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n651), .A2(KEYINPUT24), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n263), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n657), .A2(new_n658), .B1(G107), .B2(new_n479), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n665), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n592), .A2(new_n338), .ZN(new_n672));
  INV_X1    g0472(.A(new_n605), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n592), .A2(G200), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n616), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n458), .A2(new_n579), .A3(new_n678), .ZN(G372));
  NOR2_X1   g0479(.A1(new_n354), .A2(new_n355), .ZN(new_n680));
  INV_X1    g0480(.A(new_n403), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n450), .A2(new_n440), .B1(new_n681), .B2(new_n443), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n341), .A2(new_n350), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n411), .A2(new_n415), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n378), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n539), .A2(new_n578), .A3(new_n541), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT26), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT90), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n560), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n559), .A2(KEYINPUT90), .A3(new_n323), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n566), .A2(KEYINPUT91), .A3(new_n564), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT91), .B1(new_n566), .B2(new_n564), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n690), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n398), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n554), .A2(new_n567), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(G200), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n552), .A2(new_n263), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n393), .A2(new_n387), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n576), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n569), .A2(new_n570), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(G190), .B2(new_n702), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n696), .A2(new_n695), .B1(new_n698), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT26), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n539), .A4(new_n541), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n688), .A2(new_n697), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT92), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT92), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n688), .A2(new_n706), .A3(new_n709), .A4(new_n697), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n521), .A2(new_n531), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n608), .A2(new_n662), .A3(new_n611), .A4(new_n615), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n698), .A2(new_n703), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n670), .A2(new_n697), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n539), .A2(new_n541), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n711), .A2(new_n712), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n708), .A2(new_n710), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n686), .B1(new_n458), .B2(new_n718), .ZN(G369));
  NAND3_X1  g0519(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT93), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n720), .B(KEYINPUT93), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT27), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n723), .A2(new_n726), .A3(G213), .ZN(new_n727));
  XNOR2_X1  g0527(.A(KEYINPUT94), .B(G343), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT95), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(new_n653), .B2(new_n661), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT96), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n623), .A2(new_n627), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n734), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(KEYINPUT96), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n662), .A2(new_n670), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n735), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n607), .A2(new_n605), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n606), .A2(new_n580), .ZN(new_n743));
  AND4_X1   g0543(.A1(new_n742), .A2(new_n611), .A3(new_n615), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n731), .A2(new_n605), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(new_n675), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n741), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n744), .A2(new_n731), .ZN(new_n751));
  INV_X1    g0551(.A(new_n662), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT95), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n730), .B(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n740), .A2(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n750), .A2(new_n755), .ZN(G399));
  INV_X1    g0556(.A(new_n214), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G41), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n547), .A2(G116), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n759), .A2(G1), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(new_n228), .B2(new_n759), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT28), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n716), .A2(KEYINPUT99), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT99), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n542), .A2(new_n765), .A3(new_n712), .A4(new_n714), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n687), .A2(KEYINPUT98), .A3(new_n705), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n704), .A2(KEYINPUT26), .A3(new_n539), .A4(new_n541), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(KEYINPUT98), .B1(new_n687), .B2(new_n705), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n697), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(KEYINPUT29), .B(new_n754), .C1(new_n767), .C2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n670), .A2(new_n697), .A3(new_n713), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(new_n744), .B2(new_n662), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n707), .A2(KEYINPUT92), .B1(new_n775), .B2(new_n542), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n731), .B1(new_n776), .B2(new_n710), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n773), .B1(KEYINPUT29), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n540), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n560), .A2(new_n564), .A3(new_n566), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n624), .A2(new_n625), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT97), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(KEYINPUT97), .B1(new_n702), .B2(new_n622), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n607), .B(new_n779), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT30), .ZN(new_n786));
  AOI21_X1  g0586(.A(G179), .B1(new_n622), .B2(new_n510), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n787), .A2(new_n694), .A3(new_n592), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n785), .A2(new_n786), .B1(new_n788), .B2(new_n529), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n503), .A2(KEYINPUT78), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n581), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n507), .B1(new_n506), .B2(new_n508), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n317), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n323), .A2(new_n588), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n794), .A2(G179), .A3(new_n584), .A4(new_n591), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n540), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n782), .B1(new_n780), .B2(new_n781), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n702), .A2(new_n622), .A3(KEYINPUT97), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n796), .A2(new_n799), .A3(KEYINPUT30), .ZN(new_n800));
  AOI211_X1 g0600(.A(KEYINPUT31), .B(new_n754), .C1(new_n789), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT31), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n785), .A2(new_n786), .ZN(new_n803));
  AND4_X1   g0603(.A1(new_n529), .A2(new_n787), .A3(new_n694), .A4(new_n592), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n803), .A2(new_n805), .A3(new_n800), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n802), .B1(new_n806), .B2(new_n731), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n744), .A2(new_n738), .A3(new_n675), .A4(new_n754), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n801), .A2(new_n807), .B1(new_n579), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G330), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n778), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n763), .B1(new_n812), .B2(G1), .ZN(G364));
  AND2_X1   g0613(.A1(new_n211), .A2(G13), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n210), .B1(new_n814), .B2(G45), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n758), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n747), .B2(G330), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(G330), .B2(new_n747), .ZN(new_n819));
  INV_X1    g0619(.A(new_n817), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n757), .A2(new_n290), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n821), .A2(G355), .B1(new_n593), .B2(new_n757), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n757), .A2(new_n279), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n228), .B2(G45), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n254), .A2(new_n505), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(G13), .A2(G33), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT100), .Z(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(G20), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n230), .B1(G20), .B2(new_n398), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(G179), .A2(G200), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G190), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G20), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n550), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n336), .A2(G179), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(G20), .A3(G190), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n220), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n837), .A2(new_n290), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n833), .A2(G20), .A3(new_n338), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n274), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT32), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n838), .A2(G20), .A3(new_n338), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT102), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n841), .B(new_n844), .C1(new_n380), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(G20), .A2(G179), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT101), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n338), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n336), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(G200), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G68), .A2(new_n852), .B1(new_n853), .B2(G77), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n850), .A2(G190), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n336), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n855), .A2(G200), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n854), .B1(new_n249), .B2(new_n857), .C1(new_n201), .C2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G322), .A2(new_n858), .B1(new_n856), .B2(G326), .ZN(new_n861));
  INV_X1    g0661(.A(G311), .ZN(new_n862));
  INV_X1    g0662(.A(new_n853), .ZN(new_n863));
  INV_X1    g0663(.A(new_n852), .ZN(new_n864));
  XOR2_X1   g0664(.A(KEYINPUT33), .B(G317), .Z(new_n865));
  OAI221_X1 g0665(.A(new_n861), .B1(new_n862), .B2(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(G303), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n290), .B1(new_n839), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n842), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(G329), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(G294), .ZN(new_n871));
  INV_X1    g0671(.A(G283), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n870), .B1(new_n871), .B2(new_n836), .C1(new_n847), .C2(new_n872), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n848), .A2(new_n860), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n820), .B(new_n832), .C1(new_n874), .C2(new_n830), .ZN(new_n875));
  INV_X1    g0675(.A(new_n829), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n875), .B1(new_n747), .B2(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n819), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(G396));
  NAND2_X1  g0679(.A1(new_n731), .A2(new_n402), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n397), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n403), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n681), .A2(new_n754), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n777), .B(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n817), .B1(new_n886), .B2(new_n810), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n810), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n830), .A2(new_n827), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n820), .B1(new_n369), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n830), .ZN(new_n891));
  AOI22_X1  g0691(.A1(G116), .A2(new_n853), .B1(new_n856), .B2(G303), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n892), .B1(new_n872), .B2(new_n864), .C1(new_n871), .C2(new_n859), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n847), .A2(new_n220), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n290), .B1(new_n842), .B2(new_n862), .C1(new_n839), .C2(new_n380), .ZN(new_n895));
  NOR4_X1   g0695(.A1(new_n893), .A2(new_n837), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(G132), .ZN(new_n897));
  OAI221_X1 g0697(.A(new_n279), .B1(new_n842), .B2(new_n897), .C1(new_n839), .C2(new_n249), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(G58), .B2(new_n835), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n202), .B2(new_n847), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT103), .Z(new_n901));
  INV_X1    g0701(.A(KEYINPUT34), .ZN(new_n902));
  AOI22_X1  g0702(.A1(G143), .A2(new_n858), .B1(new_n853), .B2(G159), .ZN(new_n903));
  INV_X1    g0703(.A(G137), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n903), .B1(new_n904), .B2(new_n857), .C1(new_n360), .C2(new_n864), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n901), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n905), .A2(new_n902), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n896), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n890), .B1(new_n891), .B2(new_n908), .C1(new_n885), .C2(new_n828), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n888), .A2(new_n909), .ZN(G384));
  INV_X1    g0710(.A(new_n474), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n911), .A2(KEYINPUT35), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(KEYINPUT35), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n912), .A2(new_n913), .A3(G116), .A4(new_n231), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT36), .Z(new_n915));
  OAI211_X1 g0715(.A(new_n229), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n210), .B(G13), .C1(new_n916), .C2(new_n250), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT104), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n301), .A2(new_n340), .ZN(new_n921));
  INV_X1    g0721(.A(new_n299), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n344), .B2(new_n345), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n263), .B(new_n293), .C1(new_n923), .C2(KEYINPUT16), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n924), .A2(new_n270), .B1(new_n327), .B2(new_n330), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n920), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n348), .A2(new_n349), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT16), .B1(new_n346), .B2(new_n299), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n270), .B1(new_n294), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n331), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(KEYINPUT104), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n727), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n926), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT105), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT37), .B1(new_n332), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n301), .A2(KEYINPUT105), .A3(new_n331), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n301), .A2(new_n727), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n927), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n933), .A2(KEYINPUT37), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n932), .B1(new_n351), .B2(new_n356), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n919), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n932), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n454), .B2(new_n455), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT37), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n348), .A2(new_n349), .B1(new_n929), .B2(new_n331), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n943), .B1(new_n946), .B2(KEYINPUT104), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n945), .B1(new_n947), .B2(new_n926), .ZN(new_n948));
  INV_X1    g0748(.A(new_n935), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n938), .ZN(new_n950));
  OAI211_X1 g0750(.A(KEYINPUT38), .B(new_n944), .C1(new_n948), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n942), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT39), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT106), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n453), .A2(new_n353), .A3(new_n341), .A4(new_n350), .ZN(new_n956));
  INV_X1    g0756(.A(new_n937), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n921), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n945), .B1(new_n959), .B2(new_n332), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n958), .B1(new_n960), .B2(new_n950), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT39), .B1(new_n961), .B2(new_n919), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n939), .A2(new_n935), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n965), .A2(KEYINPUT106), .A3(KEYINPUT38), .A4(new_n944), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n955), .A2(new_n962), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n953), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n450), .A2(new_n440), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(new_n731), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n717), .A2(new_n754), .A3(new_n885), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n883), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n731), .A2(new_n440), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n443), .A3(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n440), .B(new_n731), .C1(new_n450), .C2(new_n444), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(new_n952), .A3(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n680), .A2(new_n727), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n971), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n773), .B(new_n457), .C1(KEYINPUT29), .C2(new_n777), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n686), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n980), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(G330), .ZN(new_n984));
  AND3_X1   g0784(.A1(new_n809), .A2(new_n977), .A3(new_n885), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n952), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT40), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n961), .A2(new_n919), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n955), .A2(new_n989), .A3(new_n966), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n796), .A2(new_n799), .A3(KEYINPUT30), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT30), .B1(new_n796), .B2(new_n799), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n991), .A2(new_n992), .A3(new_n804), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT31), .B1(new_n993), .B2(new_n754), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n806), .A2(new_n802), .A3(new_n731), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n677), .A2(new_n578), .A3(new_n542), .A4(new_n754), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n884), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n998), .A2(KEYINPUT40), .A3(new_n977), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n990), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n988), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n457), .A2(new_n809), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n984), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n983), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n210), .B2(new_n814), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n983), .A2(new_n1004), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n918), .B1(new_n1006), .B2(new_n1007), .ZN(G367));
  OAI21_X1  g0808(.A(new_n831), .B1(new_n214), .B2(new_n393), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n823), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(new_n244), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n817), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G283), .A2(new_n853), .B1(new_n856), .B2(G311), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n871), .B2(new_n864), .C1(new_n867), .C2(new_n859), .ZN(new_n1014));
  INV_X1    g0814(.A(G317), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n290), .B1(new_n842), .B2(new_n1015), .C1(new_n845), .C2(new_n550), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n839), .ZN(new_n1017));
  AOI21_X1  g0817(.A(KEYINPUT46), .B1(new_n1017), .B2(G116), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1017), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n380), .B2(new_n836), .ZN(new_n1020));
  NOR4_X1   g0820(.A1(new_n1014), .A2(new_n1016), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT114), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G50), .A2(new_n853), .B1(new_n856), .B2(G143), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n858), .A2(G150), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n836), .A2(new_n202), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n845), .A2(new_n369), .B1(new_n839), .B2(new_n201), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n279), .B1(new_n842), .B2(new_n904), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n852), .A2(G159), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1023), .A2(new_n1024), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1022), .A2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT47), .Z(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(new_n891), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n731), .A2(new_n701), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n697), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n1034), .B2(new_n704), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT107), .Z(new_n1037));
  AOI211_X1 g0837(.A(new_n1012), .B(new_n1033), .C1(new_n829), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT111), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n737), .A2(new_n739), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n735), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n1042), .A3(new_n751), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n752), .A2(new_n754), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n542), .B1(new_n525), .B2(new_n754), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n715), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n731), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1040), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n755), .A2(KEYINPUT111), .A3(new_n1049), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1054), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1051), .A2(new_n1052), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT44), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n755), .B2(new_n1049), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1045), .A2(KEYINPUT44), .A3(new_n1050), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1055), .A2(new_n1057), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n749), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT112), .B1(new_n740), .B2(new_n751), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(new_n1043), .Z(new_n1065));
  XNOR2_X1  g0865(.A(new_n748), .B(KEYINPUT113), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n747), .A2(KEYINPUT113), .A3(G330), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1067), .B1(new_n1068), .B2(new_n1065), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1053), .A2(new_n1054), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n750), .A3(new_n1057), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1063), .A2(new_n812), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n812), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n758), .B(KEYINPUT41), .Z(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n816), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT43), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1037), .A2(new_n1077), .ZN(new_n1078));
  OR3_X1    g0878(.A1(new_n1043), .A2(KEYINPUT42), .A3(new_n1050), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n662), .B1(new_n521), .B2(new_n531), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n754), .B1(new_n1080), .B2(new_n1047), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT42), .B1(new_n1043), .B2(new_n1050), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT108), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1037), .A2(new_n1077), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1084), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1078), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT108), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1078), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n1092), .A3(new_n1086), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n750), .A2(new_n1050), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1089), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT109), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1094), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1089), .A2(new_n1093), .A3(KEYINPUT109), .A4(new_n1094), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1097), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1039), .B1(new_n1076), .B2(new_n1101), .ZN(G387));
  INV_X1    g0902(.A(new_n821), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1103), .A2(new_n760), .B1(G107), .B2(new_n214), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1010), .B1(new_n241), .B2(G45), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n760), .B(new_n505), .C1(new_n202), .C2(new_n369), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT115), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n256), .A2(G50), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT50), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1108), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1104), .B1(new_n1105), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n831), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n817), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n740), .A2(new_n876), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n836), .A2(new_n393), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n279), .B1(new_n842), .B2(new_n360), .C1(new_n839), .C2(new_n369), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(G97), .C2(new_n846), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G50), .A2(new_n858), .B1(new_n856), .B2(G159), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G68), .A2(new_n853), .B1(new_n852), .B2(new_n261), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n279), .B1(new_n869), .B2(G326), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n836), .A2(new_n872), .B1(new_n839), .B2(new_n871), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G303), .A2(new_n853), .B1(new_n858), .B2(G317), .ZN(new_n1125));
  INV_X1    g0925(.A(G322), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1125), .B1(new_n862), .B2(new_n864), .C1(new_n1126), .C2(new_n857), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT48), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1124), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1128), .B2(new_n1127), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT49), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1123), .B1(new_n593), .B2(new_n845), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1122), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1115), .B(new_n1116), .C1(new_n830), .C2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n1069), .B2(new_n816), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1069), .A2(new_n812), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n758), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1069), .A2(new_n812), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1136), .B1(new_n1138), .B2(new_n1139), .ZN(G393));
  INV_X1    g0940(.A(new_n1071), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n750), .B1(new_n1070), .B2(new_n1057), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1137), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(new_n758), .A3(new_n1072), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1050), .A2(new_n829), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT116), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G150), .A2(new_n856), .B1(new_n858), .B2(G159), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT51), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n290), .B1(new_n869), .B2(G143), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1149), .B1(new_n202), .B2(new_n839), .C1(new_n369), .C2(new_n836), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n249), .A2(new_n864), .B1(new_n863), .B2(new_n256), .ZN(new_n1151));
  OR4_X1    g0951(.A1(new_n894), .A2(new_n1148), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G311), .A2(new_n858), .B1(new_n856), .B2(G317), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT52), .Z(new_n1154));
  NOR2_X1   g0954(.A1(new_n836), .A2(new_n593), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n290), .B1(new_n842), .B2(new_n1126), .C1(new_n839), .C2(new_n872), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(G107), .C2(new_n846), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G294), .A2(new_n853), .B1(new_n852), .B2(G303), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1154), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n891), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n831), .B1(new_n550), .B2(new_n214), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1010), .A2(new_n248), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n817), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1146), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n816), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1144), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT117), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT117), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1144), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(G390));
  INV_X1    g0971(.A(new_n970), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n754), .B(new_n882), .C1(new_n767), .C2(new_n772), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1173), .A2(new_n883), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n977), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1172), .B(new_n990), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n972), .B2(new_n883), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n953), .B(new_n967), .C1(new_n1177), .C2(new_n970), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  AND4_X1   g0979(.A1(G330), .A2(new_n809), .A3(new_n885), .A4(new_n977), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n809), .A2(new_n977), .A3(new_n885), .A4(G330), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1176), .A2(new_n1178), .A3(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n816), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT119), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1181), .A2(KEYINPUT119), .A3(new_n816), .A4(new_n1183), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT118), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n977), .B1(new_n998), .B2(G330), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n973), .B1(new_n1190), .B2(new_n1180), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n809), .A2(G330), .A3(new_n885), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1175), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1193), .A2(new_n883), .A3(new_n1173), .A4(new_n1182), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n457), .A2(G330), .A3(new_n809), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n981), .A2(new_n686), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1189), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n981), .A2(new_n686), .A3(new_n1196), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT118), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1183), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1182), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1198), .B(new_n1201), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT118), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT118), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1181), .B(new_n1183), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1204), .A2(new_n1207), .A3(new_n758), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n889), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n817), .B1(new_n261), .B2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G97), .A2(new_n853), .B1(new_n856), .B2(G283), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n380), .B2(new_n864), .C1(new_n593), .C2(new_n859), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n279), .B(new_n840), .C1(G294), .C2(new_n869), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n369), .B2(new_n836), .C1(new_n202), .C2(new_n847), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT54), .B(G143), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT120), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G137), .A2(new_n852), .B1(new_n853), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n897), .B2(new_n859), .ZN(new_n1218));
  INV_X1    g1018(.A(G125), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n279), .B1(new_n842), .B2(new_n1219), .C1(new_n845), .C2(new_n249), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n856), .A2(G128), .B1(new_n1220), .B2(KEYINPUT121), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1017), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT53), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n839), .B2(new_n360), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1222), .A2(new_n1224), .B1(G159), .B2(new_n835), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1221), .B(new_n1225), .C1(KEYINPUT121), .C2(new_n1220), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1212), .A2(new_n1214), .B1(new_n1218), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1210), .B1(new_n1227), .B2(new_n830), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n968), .B2(new_n828), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1188), .A2(new_n1208), .A3(new_n1229), .ZN(G378));
  NAND2_X1  g1030(.A1(new_n365), .A2(new_n727), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n378), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1231), .B1(new_n685), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n685), .A2(new_n1232), .A3(new_n1231), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  AND4_X1   g1039(.A1(G330), .A2(new_n988), .A3(new_n1000), .A4(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1239), .B1(new_n1241), .B2(new_n1000), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n980), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n988), .A2(new_n1000), .A3(G330), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1239), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n978), .A2(new_n979), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1172), .B1(new_n953), .B2(new_n967), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1241), .A2(new_n1000), .A3(new_n1239), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1246), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1243), .A2(new_n1251), .A3(KEYINPUT122), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT122), .B1(new_n1243), .B2(new_n1251), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1207), .A2(new_n1199), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT57), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1243), .A2(new_n1251), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(KEYINPUT57), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n758), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1239), .A2(new_n828), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n817), .B1(G50), .B2(new_n1209), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n279), .A2(G41), .ZN(new_n1263));
  AOI211_X1 g1063(.A(G50), .B(new_n1263), .C1(new_n284), .C2(new_n497), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n380), .A2(new_n859), .B1(new_n857), .B2(new_n593), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G97), .B2(new_n852), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1263), .B1(new_n201), .B2(new_n845), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n839), .A2(new_n369), .B1(new_n842), .B2(new_n872), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1025), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1266), .B(new_n1269), .C1(new_n393), .C2(new_n863), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT58), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1264), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n284), .B(new_n497), .C1(new_n845), .C2(new_n274), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(G124), .B2(new_n869), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(G128), .A2(new_n858), .B1(new_n853), .B2(G137), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n897), .B2(new_n864), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1216), .A2(new_n1017), .B1(G150), .B2(new_n835), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n857), .B2(new_n1219), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT59), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1274), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1279), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1282), .A2(KEYINPUT59), .ZN(new_n1283));
  OAI221_X1 g1083(.A(new_n1272), .B1(new_n1271), .B2(new_n1270), .C1(new_n1281), .C2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1262), .B1(new_n1284), .B2(new_n830), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1261), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1254), .B2(new_n816), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1260), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(G375));
  NOR2_X1   g1091(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1292), .A2(new_n1075), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1175), .A2(new_n827), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n817), .B1(G68), .B2(new_n1209), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(G107), .A2(new_n853), .B1(new_n856), .B2(G294), .ZN(new_n1297));
  OAI221_X1 g1097(.A(new_n1297), .B1(new_n593), .B2(new_n864), .C1(new_n872), .C2(new_n859), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n290), .B1(new_n839), .B2(new_n550), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n1299), .B(new_n1117), .C1(G303), .C2(new_n869), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n369), .B2(new_n847), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n839), .A2(new_n274), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n279), .B1(new_n845), .B2(new_n201), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n1302), .B(new_n1303), .C1(G128), .C2(new_n869), .ZN(new_n1304));
  OAI221_X1 g1104(.A(new_n1304), .B1(new_n249), .B2(new_n836), .C1(new_n360), .C2(new_n863), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(G137), .A2(new_n858), .B1(new_n852), .B2(new_n1216), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n897), .B2(new_n857), .ZN(new_n1307));
  OAI22_X1  g1107(.A1(new_n1298), .A2(new_n1301), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  OR2_X1    g1108(.A1(new_n1308), .A2(KEYINPUT123), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n891), .B1(new_n1308), .B2(KEYINPUT123), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1296), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  AOI22_X1  g1111(.A1(new_n1200), .A2(new_n816), .B1(new_n1295), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1294), .A2(new_n1312), .ZN(G381));
  OR2_X1    g1113(.A1(G393), .A2(G396), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(G390), .A2(G384), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(G387), .ZN(new_n1316));
  INV_X1    g1116(.A(G381), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1315), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(KEYINPUT124), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT125), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G378), .A2(new_n1320), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1188), .A2(new_n1208), .A3(KEYINPUT125), .A4(new_n1229), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT124), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1315), .A2(new_n1325), .A3(new_n1316), .A4(new_n1317), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1319), .A2(new_n1290), .A3(new_n1324), .A4(new_n1326), .ZN(G407));
  NAND2_X1  g1127(.A1(new_n728), .A2(G213), .ZN(new_n1328));
  XOR2_X1   g1128(.A(new_n1328), .B(KEYINPUT126), .Z(new_n1329));
  NAND3_X1  g1129(.A1(new_n1290), .A2(new_n1324), .A3(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(G407), .A2(new_n1330), .A3(G213), .ZN(G409));
  NAND3_X1  g1131(.A1(new_n1198), .A2(new_n1201), .A3(new_n1293), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(KEYINPUT60), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT60), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1334), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n758), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(KEYINPUT127), .B1(new_n1333), .B2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT127), .ZN(new_n1339));
  AOI211_X1 g1139(.A(new_n1339), .B(new_n1336), .C1(new_n1332), .C2(KEYINPUT60), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1312), .B1(new_n1338), .B2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(G384), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  OAI211_X1 g1143(.A(G384), .B(new_n1312), .C1(new_n1338), .C2(new_n1340), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1329), .A2(G2897), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1343), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1345), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  OAI211_X1 g1148(.A(G378), .B(new_n1288), .C1(new_n1256), .C2(new_n1259), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT122), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1257), .A2(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1243), .A2(new_n1251), .A3(KEYINPUT122), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1351), .A2(new_n1255), .A3(new_n1075), .A4(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1287), .B1(new_n1257), .B2(new_n816), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1321), .A2(new_n1355), .A3(new_n1322), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1349), .A2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1329), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1159(.A(KEYINPUT61), .B1(new_n1348), .B2(new_n1359), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(G387), .A2(new_n1170), .A3(new_n1168), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1098), .B1(new_n1096), .B2(new_n1095), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1074), .B1(new_n1072), .B2(new_n812), .ZN(new_n1363));
  OAI211_X1 g1163(.A(new_n1362), .B(new_n1100), .C1(new_n1363), .C2(new_n816), .ZN(new_n1364));
  AND3_X1   g1164(.A1(new_n1144), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1169), .B1(new_n1144), .B2(new_n1166), .ZN(new_n1366));
  OAI211_X1 g1166(.A(new_n1364), .B(new_n1039), .C1(new_n1365), .C2(new_n1366), .ZN(new_n1367));
  XNOR2_X1  g1167(.A(G393), .B(new_n878), .ZN(new_n1368));
  AND3_X1   g1168(.A1(new_n1361), .A2(new_n1367), .A3(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1368), .B1(new_n1361), .B2(new_n1367), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT63), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1334), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1373));
  OAI21_X1  g1173(.A(new_n1339), .B1(new_n1373), .B2(new_n1336), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1333), .A2(KEYINPUT127), .A3(new_n1337), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1374), .A2(new_n1375), .ZN(new_n1376));
  AOI21_X1  g1176(.A(G384), .B1(new_n1376), .B2(new_n1312), .ZN(new_n1377));
  INV_X1    g1177(.A(new_n1344), .ZN(new_n1378));
  NOR2_X1   g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1379), .ZN(new_n1380));
  OAI21_X1  g1180(.A(new_n1372), .B1(new_n1359), .B2(new_n1380), .ZN(new_n1381));
  AOI21_X1  g1181(.A(new_n1329), .B1(new_n1349), .B2(new_n1356), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1382), .A2(KEYINPUT63), .A3(new_n1379), .ZN(new_n1383));
  NAND4_X1  g1183(.A1(new_n1360), .A2(new_n1371), .A3(new_n1381), .A4(new_n1383), .ZN(new_n1384));
  INV_X1    g1184(.A(KEYINPUT61), .ZN(new_n1385));
  INV_X1    g1185(.A(new_n1345), .ZN(new_n1386));
  OAI21_X1  g1186(.A(new_n1386), .B1(new_n1377), .B2(new_n1378), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n1343), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1387), .A2(new_n1388), .ZN(new_n1389));
  OAI21_X1  g1189(.A(new_n1385), .B1(new_n1389), .B2(new_n1382), .ZN(new_n1390));
  INV_X1    g1190(.A(KEYINPUT62), .ZN(new_n1391));
  AND4_X1   g1191(.A1(new_n1391), .A2(new_n1357), .A3(new_n1358), .A4(new_n1379), .ZN(new_n1392));
  AOI21_X1  g1192(.A(new_n1391), .B1(new_n1382), .B2(new_n1379), .ZN(new_n1393));
  NOR3_X1   g1193(.A1(new_n1390), .A2(new_n1392), .A3(new_n1393), .ZN(new_n1394));
  OAI21_X1  g1194(.A(new_n1384), .B1(new_n1394), .B2(new_n1371), .ZN(G405));
  OAI21_X1  g1195(.A(new_n1324), .B1(new_n1260), .B2(new_n1289), .ZN(new_n1396));
  AOI21_X1  g1196(.A(new_n1380), .B1(new_n1396), .B2(new_n1349), .ZN(new_n1397));
  INV_X1    g1197(.A(new_n1397), .ZN(new_n1398));
  NAND3_X1  g1198(.A1(new_n1380), .A2(new_n1396), .A3(new_n1349), .ZN(new_n1399));
  NAND3_X1  g1199(.A1(new_n1398), .A2(new_n1371), .A3(new_n1399), .ZN(new_n1400));
  INV_X1    g1200(.A(new_n1399), .ZN(new_n1401));
  OAI22_X1  g1201(.A1(new_n1401), .A2(new_n1397), .B1(new_n1369), .B2(new_n1370), .ZN(new_n1402));
  NAND2_X1  g1202(.A1(new_n1400), .A2(new_n1402), .ZN(G402));
endmodule


