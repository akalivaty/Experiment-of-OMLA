

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589;

  XNOR2_X1 U321 ( .A(n366), .B(n365), .ZN(n382) );
  INV_X1 U322 ( .A(G92GAT), .ZN(n348) );
  XNOR2_X1 U323 ( .A(n355), .B(n312), .ZN(n318) );
  NOR2_X1 U324 ( .A1(n290), .A2(n524), .ZN(n574) );
  XNOR2_X1 U325 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U326 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n326) );
  AND2_X1 U327 ( .A1(G231GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U328 ( .A(KEYINPUT54), .B(n397), .Z(n290) );
  NOR2_X1 U329 ( .A1(n367), .A2(n374), .ZN(n375) );
  XNOR2_X1 U330 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n365) );
  XOR2_X1 U331 ( .A(G1GAT), .B(G127GAT), .Z(n407) );
  XNOR2_X1 U332 ( .A(n311), .B(KEYINPUT76), .ZN(n312) );
  XNOR2_X1 U333 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U334 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U335 ( .A(n337), .B(n289), .ZN(n338) );
  XNOR2_X1 U336 ( .A(n339), .B(n338), .ZN(n343) );
  XNOR2_X1 U337 ( .A(n359), .B(n358), .ZN(n363) );
  XNOR2_X1 U338 ( .A(n367), .B(n326), .ZN(n558) );
  XNOR2_X1 U339 ( .A(n466), .B(G190GAT), .ZN(n467) );
  XNOR2_X1 U340 ( .A(n468), .B(n467), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n291) );
  XNOR2_X1 U342 ( .A(n291), .B(KEYINPUT7), .ZN(n351) );
  XOR2_X1 U343 ( .A(G22GAT), .B(G15GAT), .Z(n330) );
  XOR2_X1 U344 ( .A(n351), .B(n330), .Z(n293) );
  NAND2_X1 U345 ( .A1(G229GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U346 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U347 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n295) );
  XNOR2_X1 U348 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U350 ( .A(n297), .B(n296), .Z(n305) );
  XOR2_X1 U351 ( .A(G197GAT), .B(G50GAT), .Z(n299) );
  XNOR2_X1 U352 ( .A(G36GAT), .B(G29GAT), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U354 ( .A(G1GAT), .B(G113GAT), .Z(n301) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(G141GAT), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n575) );
  XNOR2_X1 U359 ( .A(G120GAT), .B(G148GAT), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n306), .B(G57GAT), .ZN(n398) );
  XOR2_X1 U361 ( .A(G64GAT), .B(G92GAT), .Z(n308) );
  XNOR2_X1 U362 ( .A(G176GAT), .B(G204GAT), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n387) );
  XNOR2_X1 U364 ( .A(n398), .B(n387), .ZN(n325) );
  XOR2_X1 U365 ( .A(KEYINPUT73), .B(G85GAT), .Z(n310) );
  XNOR2_X1 U366 ( .A(G99GAT), .B(G106GAT), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n355) );
  INV_X1 U368 ( .A(KEYINPUT31), .ZN(n311) );
  INV_X1 U369 ( .A(KEYINPUT32), .ZN(n314) );
  XNOR2_X1 U370 ( .A(G71GAT), .B(G78GAT), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n313), .B(KEYINPUT13), .ZN(n341) );
  XNOR2_X1 U372 ( .A(n314), .B(n341), .ZN(n316) );
  NAND2_X1 U373 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U374 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n323) );
  XOR2_X1 U376 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n320) );
  XNOR2_X1 U377 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U379 ( .A(KEYINPUT72), .B(n321), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n367) );
  NOR2_X1 U382 ( .A1(n575), .A2(n558), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n327), .B(KEYINPUT46), .ZN(n344) );
  XOR2_X1 U384 ( .A(KEYINPUT82), .B(KEYINPUT84), .Z(n329) );
  XNOR2_X1 U385 ( .A(KEYINPUT15), .B(KEYINPUT83), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n334) );
  XOR2_X1 U387 ( .A(n407), .B(G57GAT), .Z(n332) );
  XNOR2_X1 U388 ( .A(n330), .B(G155GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U390 ( .A(n334), .B(n333), .Z(n339) );
  XOR2_X1 U391 ( .A(KEYINPUT85), .B(KEYINPUT14), .Z(n336) );
  XNOR2_X1 U392 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U394 ( .A(G8GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n340), .B(G211GAT), .ZN(n386) );
  XNOR2_X1 U396 ( .A(n386), .B(n341), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n583) );
  XOR2_X1 U398 ( .A(KEYINPUT111), .B(n583), .Z(n547) );
  NOR2_X1 U399 ( .A1(n344), .A2(n547), .ZN(n345) );
  XNOR2_X1 U400 ( .A(KEYINPUT112), .B(n345), .ZN(n364) );
  XOR2_X1 U401 ( .A(KEYINPUT80), .B(KEYINPUT78), .Z(n347) );
  XNOR2_X1 U402 ( .A(KEYINPUT9), .B(KEYINPUT10), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n353) );
  NAND2_X1 U404 ( .A1(G232GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n359) );
  XNOR2_X1 U406 ( .A(G36GAT), .B(G190GAT), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n354), .B(G218GAT), .ZN(n390) );
  XNOR2_X1 U408 ( .A(n390), .B(n355), .ZN(n357) );
  XOR2_X1 U409 ( .A(G50GAT), .B(G162GAT), .Z(n423) );
  XOR2_X1 U410 ( .A(G29GAT), .B(G134GAT), .Z(n408) );
  XOR2_X1 U411 ( .A(n423), .B(n408), .Z(n356) );
  XOR2_X1 U412 ( .A(KEYINPUT11), .B(KEYINPUT65), .Z(n361) );
  XNOR2_X1 U413 ( .A(KEYINPUT67), .B(KEYINPUT79), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n363), .B(n362), .ZN(n568) );
  NAND2_X1 U416 ( .A1(n364), .A2(n568), .ZN(n366) );
  XNOR2_X1 U417 ( .A(n568), .B(KEYINPUT81), .ZN(n464) );
  NAND2_X1 U418 ( .A1(KEYINPUT36), .A2(n464), .ZN(n371) );
  INV_X1 U419 ( .A(KEYINPUT36), .ZN(n369) );
  INV_X1 U420 ( .A(n464), .ZN(n368) );
  NAND2_X1 U421 ( .A1(n369), .A2(n368), .ZN(n370) );
  NAND2_X1 U422 ( .A1(n371), .A2(n370), .ZN(n585) );
  NAND2_X1 U423 ( .A1(n583), .A2(n585), .ZN(n373) );
  XOR2_X1 U424 ( .A(KEYINPUT68), .B(KEYINPUT45), .Z(n372) );
  XOR2_X1 U425 ( .A(n373), .B(n372), .Z(n374) );
  NAND2_X1 U426 ( .A1(KEYINPUT114), .A2(n375), .ZN(n379) );
  INV_X1 U427 ( .A(KEYINPUT114), .ZN(n377) );
  INV_X1 U428 ( .A(n375), .ZN(n376) );
  NAND2_X1 U429 ( .A1(n377), .A2(n376), .ZN(n378) );
  NAND2_X1 U430 ( .A1(n379), .A2(n378), .ZN(n380) );
  NAND2_X1 U431 ( .A1(n380), .A2(n575), .ZN(n381) );
  NAND2_X1 U432 ( .A1(n382), .A2(n381), .ZN(n383) );
  XNOR2_X1 U433 ( .A(n383), .B(KEYINPUT48), .ZN(n537) );
  XOR2_X1 U434 ( .A(G197GAT), .B(KEYINPUT21), .Z(n422) );
  XOR2_X1 U435 ( .A(KEYINPUT96), .B(n422), .Z(n385) );
  NAND2_X1 U436 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n394) );
  XOR2_X1 U438 ( .A(n387), .B(n386), .Z(n392) );
  XOR2_X1 U439 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n389) );
  XNOR2_X1 U440 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n388) );
  XNOR2_X1 U441 ( .A(n389), .B(n388), .ZN(n447) );
  XNOR2_X1 U442 ( .A(n447), .B(n390), .ZN(n391) );
  XNOR2_X1 U443 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U444 ( .A(n394), .B(n393), .Z(n527) );
  XNOR2_X1 U445 ( .A(KEYINPUT122), .B(n527), .ZN(n395) );
  NAND2_X1 U446 ( .A1(n537), .A2(n395), .ZN(n396) );
  XNOR2_X1 U447 ( .A(n396), .B(KEYINPUT123), .ZN(n397) );
  XOR2_X1 U448 ( .A(n398), .B(KEYINPUT91), .Z(n400) );
  NAND2_X1 U449 ( .A1(G225GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U450 ( .A(n400), .B(n399), .ZN(n415) );
  XOR2_X1 U451 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n402) );
  XNOR2_X1 U452 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n401) );
  XNOR2_X1 U453 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U454 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n404) );
  XNOR2_X1 U455 ( .A(KEYINPUT5), .B(KEYINPUT90), .ZN(n403) );
  XNOR2_X1 U456 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U457 ( .A(n406), .B(n405), .Z(n413) );
  XOR2_X1 U458 ( .A(G113GAT), .B(KEYINPUT0), .Z(n443) );
  XOR2_X1 U459 ( .A(G85GAT), .B(n407), .Z(n410) );
  XNOR2_X1 U460 ( .A(G162GAT), .B(n408), .ZN(n409) );
  XNOR2_X1 U461 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U462 ( .A(n443), .B(n411), .ZN(n412) );
  XNOR2_X1 U463 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U464 ( .A(n415), .B(n414), .ZN(n421) );
  XNOR2_X1 U465 ( .A(KEYINPUT89), .B(KEYINPUT3), .ZN(n416) );
  XNOR2_X1 U466 ( .A(n416), .B(KEYINPUT88), .ZN(n417) );
  XOR2_X1 U467 ( .A(n417), .B(KEYINPUT2), .Z(n419) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(G155GAT), .ZN(n418) );
  XNOR2_X1 U469 ( .A(n419), .B(n418), .ZN(n436) );
  INV_X1 U470 ( .A(n436), .ZN(n420) );
  XNOR2_X1 U471 ( .A(n421), .B(n420), .ZN(n481) );
  XNOR2_X1 U472 ( .A(KEYINPUT95), .B(n481), .ZN(n524) );
  XOR2_X1 U473 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n425) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U475 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U476 ( .A(n426), .B(G106GAT), .Z(n431) );
  XOR2_X1 U477 ( .A(G78GAT), .B(G148GAT), .Z(n428) );
  XNOR2_X1 U478 ( .A(G22GAT), .B(G204GAT), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U480 ( .A(n429), .B(G218GAT), .ZN(n430) );
  XNOR2_X1 U481 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U482 ( .A(KEYINPUT23), .B(KEYINPUT72), .Z(n433) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U485 ( .A(n435), .B(n434), .Z(n438) );
  XNOR2_X1 U486 ( .A(n436), .B(G211GAT), .ZN(n437) );
  XNOR2_X1 U487 ( .A(n438), .B(n437), .ZN(n476) );
  NAND2_X1 U488 ( .A1(n574), .A2(n476), .ZN(n439) );
  XNOR2_X1 U489 ( .A(n439), .B(KEYINPUT55), .ZN(n458) );
  XOR2_X1 U490 ( .A(G134GAT), .B(G99GAT), .Z(n441) );
  XNOR2_X1 U491 ( .A(G43GAT), .B(G190GAT), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U493 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U495 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U496 ( .A(n446), .B(G71GAT), .Z(n449) );
  XNOR2_X1 U497 ( .A(G15GAT), .B(n447), .ZN(n448) );
  XNOR2_X1 U498 ( .A(n449), .B(n448), .ZN(n457) );
  XOR2_X1 U499 ( .A(G127GAT), .B(G176GAT), .Z(n451) );
  XNOR2_X1 U500 ( .A(G120GAT), .B(KEYINPUT87), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n451), .B(n450), .ZN(n455) );
  XOR2_X1 U502 ( .A(G183GAT), .B(KEYINPUT66), .Z(n453) );
  XNOR2_X1 U503 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n452) );
  XNOR2_X1 U504 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U505 ( .A(n455), .B(n454), .Z(n456) );
  XNOR2_X1 U506 ( .A(n457), .B(n456), .ZN(n539) );
  NAND2_X1 U507 ( .A1(n458), .A2(n539), .ZN(n571) );
  XNOR2_X1 U508 ( .A(n558), .B(KEYINPUT104), .ZN(n542) );
  NOR2_X1 U509 ( .A1(n571), .A2(n542), .ZN(n461) );
  XNOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n459), .B(G176GAT), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  INV_X1 U513 ( .A(n571), .ZN(n465) );
  NAND2_X1 U514 ( .A1(n465), .A2(n547), .ZN(n463) );
  XNOR2_X1 U515 ( .A(KEYINPUT124), .B(G183GAT), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n463), .B(n462), .ZN(G1350GAT) );
  NAND2_X1 U517 ( .A1(n465), .A2(n464), .ZN(n468) );
  XOR2_X1 U518 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n466) );
  XOR2_X1 U519 ( .A(KEYINPUT98), .B(KEYINPUT34), .Z(n487) );
  NOR2_X1 U520 ( .A1(n367), .A2(n575), .ZN(n469) );
  XNOR2_X1 U521 ( .A(n469), .B(KEYINPUT77), .ZN(n499) );
  INV_X1 U522 ( .A(n583), .ZN(n564) );
  NOR2_X1 U523 ( .A1(n464), .A2(n564), .ZN(n470) );
  XNOR2_X1 U524 ( .A(n470), .B(KEYINPUT16), .ZN(n485) );
  XNOR2_X1 U525 ( .A(n476), .B(KEYINPUT69), .ZN(n471) );
  XNOR2_X1 U526 ( .A(n471), .B(KEYINPUT28), .ZN(n538) );
  NOR2_X1 U527 ( .A1(n538), .A2(n539), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n527), .B(KEYINPUT27), .ZN(n478) );
  AND2_X1 U529 ( .A1(n478), .A2(n524), .ZN(n536) );
  NAND2_X1 U530 ( .A1(n472), .A2(n536), .ZN(n484) );
  NAND2_X1 U531 ( .A1(n539), .A2(n527), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n473), .A2(n476), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n474), .B(KEYINPUT97), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT25), .ZN(n480) );
  NOR2_X1 U535 ( .A1(n539), .A2(n476), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n477), .B(KEYINPUT26), .ZN(n573) );
  NAND2_X1 U537 ( .A1(n478), .A2(n573), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n480), .A2(n479), .ZN(n482) );
  NAND2_X1 U539 ( .A1(n482), .A2(n481), .ZN(n483) );
  NAND2_X1 U540 ( .A1(n484), .A2(n483), .ZN(n496) );
  NAND2_X1 U541 ( .A1(n485), .A2(n496), .ZN(n511) );
  NOR2_X1 U542 ( .A1(n499), .A2(n511), .ZN(n493) );
  NAND2_X1 U543 ( .A1(n493), .A2(n524), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U545 ( .A(G1GAT), .B(n488), .Z(G1324GAT) );
  XOR2_X1 U546 ( .A(G8GAT), .B(KEYINPUT99), .Z(n490) );
  NAND2_X1 U547 ( .A1(n493), .A2(n527), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U550 ( .A1(n493), .A2(n539), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  NAND2_X1 U552 ( .A1(n493), .A2(n538), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n494), .B(KEYINPUT100), .ZN(n495) );
  XNOR2_X1 U554 ( .A(G22GAT), .B(n495), .ZN(G1327GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT39), .B(KEYINPUT101), .Z(n502) );
  NAND2_X1 U556 ( .A1(n585), .A2(n496), .ZN(n497) );
  NOR2_X1 U557 ( .A1(n497), .A2(n583), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(KEYINPUT37), .ZN(n523) );
  NOR2_X1 U559 ( .A1(n523), .A2(n499), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT38), .B(n500), .ZN(n508) );
  NAND2_X1 U561 ( .A1(n524), .A2(n508), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U563 ( .A(G29GAT), .B(n503), .Z(G1328GAT) );
  NAND2_X1 U564 ( .A1(n508), .A2(n527), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n504), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT102), .B(KEYINPUT40), .Z(n506) );
  NAND2_X1 U567 ( .A1(n508), .A2(n539), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U569 ( .A(G43GAT), .B(n507), .Z(G1330GAT) );
  NAND2_X1 U570 ( .A1(n508), .A2(n538), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U572 ( .A(G57GAT), .B(KEYINPUT103), .Z(n513) );
  INV_X1 U573 ( .A(n542), .ZN(n510) );
  NAND2_X1 U574 ( .A1(n575), .A2(n510), .ZN(n522) );
  NOR2_X1 U575 ( .A1(n522), .A2(n511), .ZN(n519) );
  NAND2_X1 U576 ( .A1(n519), .A2(n524), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(n515) );
  XOR2_X1 U578 ( .A(KEYINPUT42), .B(KEYINPUT105), .Z(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U580 ( .A1(n519), .A2(n527), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(KEYINPUT106), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G64GAT), .B(n517), .ZN(G1333GAT) );
  NAND2_X1 U583 ( .A1(n539), .A2(n519), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U586 ( .A1(n519), .A2(n538), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  XOR2_X1 U588 ( .A(G85GAT), .B(KEYINPUT107), .Z(n526) );
  NOR2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n532) );
  NAND2_X1 U590 ( .A1(n532), .A2(n524), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n532), .A2(n527), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n530) );
  NAND2_X1 U595 ( .A1(n532), .A2(n539), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n534) );
  NAND2_X1 U599 ( .A1(n532), .A2(n538), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U601 ( .A(G106GAT), .B(n535), .Z(G1339GAT) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n554) );
  NOR2_X1 U603 ( .A1(n538), .A2(n554), .ZN(n540) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n546) );
  NOR2_X1 U605 ( .A1(n575), .A2(n546), .ZN(n541) );
  XOR2_X1 U606 ( .A(G113GAT), .B(n541), .Z(G1340GAT) );
  NOR2_X1 U607 ( .A1(n542), .A2(n546), .ZN(n544) );
  XNOR2_X1 U608 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U610 ( .A(G120GAT), .B(n545), .Z(G1341GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n549) );
  INV_X1 U612 ( .A(n546), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n551), .A2(n547), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n550), .Z(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U617 ( .A1(n551), .A2(n464), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  INV_X1 U619 ( .A(n554), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n555), .A2(n573), .ZN(n567) );
  NOR2_X1 U621 ( .A1(n575), .A2(n567), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1344GAT) );
  NOR2_X1 U624 ( .A1(n558), .A2(n567), .ZN(n563) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n560) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(KEYINPUT118), .B(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n567), .ZN(n565) );
  XOR2_X1 U631 ( .A(G155GAT), .B(n565), .Z(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT120), .B(n566), .ZN(G1346GAT) );
  NOR2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n570) );
  XNOR2_X1 U634 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1347GAT) );
  NOR2_X1 U636 ( .A1(n575), .A2(n571), .ZN(n572) );
  XOR2_X1 U637 ( .A(G169GAT), .B(n572), .Z(G1348GAT) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n579) );
  NOR2_X1 U639 ( .A1(n575), .A2(n579), .ZN(n577) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n581) );
  INV_X1 U644 ( .A(n579), .ZN(n586) );
  NAND2_X1 U645 ( .A1(n586), .A2(n367), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n586), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n588) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

