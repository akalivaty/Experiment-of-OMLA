//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT64), .ZN(G261));
  AOI21_X1  g031(.A(KEYINPUT65), .B1(new_n452), .B2(G2106), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n457), .B1(G567), .B2(new_n454), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n452), .A2(KEYINPUT65), .A3(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(G125), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n463), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  OAI211_X1 g050(.A(G137), .B(new_n467), .C1(new_n469), .C2(new_n470), .ZN(new_n476));
  INV_X1    g051(.A(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n469), .A2(new_n470), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n467), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n484), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n487), .A2(new_n493), .A3(G138), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n467), .C1(new_n469), .C2(new_n470), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n483), .A2(G126), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT67), .B(G114), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT68), .B1(new_n502), .B2(G2105), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT67), .A2(G114), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT67), .A2(G114), .ZN(new_n505));
  OAI211_X1 g080(.A(KEYINPUT68), .B(G2105), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n501), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT69), .ZN(new_n509));
  OAI21_X1  g084(.A(G2105), .B1(new_n504), .B2(new_n505), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n500), .B1(new_n512), .B2(new_n506), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n499), .B1(new_n509), .B2(new_n515), .ZN(G164));
  NAND2_X1  g091(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n524), .A2(new_n530), .ZN(G166));
  NAND3_X1  g106(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT72), .B(G89), .ZN(new_n534));
  OAI221_X1 g109(.A(new_n532), .B1(new_n528), .B2(new_n533), .C1(new_n526), .C2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT71), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT7), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n535), .A2(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n523), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n525), .A2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G52), .ZN(new_n545));
  INV_X1    g120(.A(new_n526), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G90), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n521), .A2(G56), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n523), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(KEYINPUT73), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n525), .A2(G43), .A3(G543), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n526), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n552), .A2(KEYINPUT73), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(new_n521), .A2(G65), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT75), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n523), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OR3_X1    g145(.A1(new_n528), .A2(KEYINPUT9), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT9), .B1(new_n528), .B2(new_n570), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n569), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n526), .A2(KEYINPUT74), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT74), .B1(new_n526), .B2(new_n574), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G299));
  OR2_X1    g153(.A1(new_n535), .A2(new_n539), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  AOI22_X1  g155(.A1(new_n546), .A2(G87), .B1(new_n544), .B2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  NAND3_X1  g158(.A1(new_n544), .A2(KEYINPUT77), .A3(G48), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n585));
  INV_X1    g160(.A(G48), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n528), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n584), .A2(new_n587), .B1(new_n546), .B2(G86), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n521), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n523), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n591), .A2(KEYINPUT76), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n591), .A2(KEYINPUT76), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n588), .B1(new_n592), .B2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n546), .A2(G85), .B1(new_n544), .B2(G47), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n523), .B2(new_n596), .ZN(G290));
  INV_X1    g172(.A(G868), .ZN(new_n598));
  NOR2_X1   g173(.A1(G301), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n546), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n526), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n600), .A2(new_n603), .B1(G54), .B2(new_n544), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT78), .B(G66), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n521), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G79), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n518), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n606), .B(KEYINPUT79), .C1(new_n607), .C2(new_n518), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n610), .A2(G651), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT80), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n604), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n613), .B1(new_n604), .B2(new_n612), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n599), .B1(new_n617), .B2(new_n598), .ZN(G321));
  XOR2_X1   g193(.A(G321), .B(KEYINPUT81), .Z(G284));
  NAND2_X1  g194(.A1(G299), .A2(new_n598), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n598), .B2(G168), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(new_n598), .B2(G168), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT82), .ZN(G148));
  NOR2_X1   g200(.A1(new_n560), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(new_n616), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n627), .A2(new_n623), .A3(new_n614), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n626), .B1(new_n628), .B2(G868), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n465), .A2(new_n478), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(G2100), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT84), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT85), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n483), .A2(G123), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n487), .A2(G135), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n467), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n637), .A2(new_n639), .A3(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT86), .ZN(new_n660));
  INV_X1    g235(.A(G14), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n657), .B2(new_n658), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(KEYINPUT17), .ZN(new_n671));
  INV_X1    g246(.A(new_n665), .ZN(new_n672));
  INV_X1    g247(.A(new_n666), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n668), .A3(new_n673), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(new_n667), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n670), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n685), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n687), .B(new_n690), .C1(new_n682), .C2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT88), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n694), .B(new_n698), .ZN(G229));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G32), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n483), .A2(G129), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n487), .A2(G141), .B1(G105), .B2(new_n478), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT26), .Z(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT95), .Z(new_n707));
  OAI21_X1  g282(.A(new_n701), .B1(new_n707), .B2(new_n700), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT96), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n708), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n700), .A2(G35), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G162), .B2(new_n700), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT29), .Z(new_n714));
  INV_X1    g289(.A(G2090), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n700), .B1(KEYINPUT24), .B2(G34), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(KEYINPUT24), .B2(G34), .ZN(new_n718));
  INV_X1    g293(.A(G160), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G29), .ZN(new_n720));
  INV_X1    g295(.A(G2084), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n700), .A2(G26), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n483), .A2(G128), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n487), .A2(G140), .ZN(new_n726));
  OR2_X1    g301(.A1(G104), .A2(G2105), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(new_n700), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2067), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT31), .B(G11), .Z(new_n733));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n700), .B1(new_n734), .B2(G28), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT97), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n735), .A2(new_n736), .B1(new_n734), .B2(G28), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n644), .B2(new_n700), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT98), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n732), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n700), .A2(G33), .ZN(new_n743));
  NAND2_X1  g318(.A1(G115), .A2(G2104), .ZN(new_n744));
  INV_X1    g319(.A(G127), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n482), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n467), .B1(new_n746), .B2(KEYINPUT94), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT94), .B2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT25), .ZN(new_n749));
  NAND2_X1  g324(.A1(G103), .A2(G2104), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G2105), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n487), .A2(G139), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n743), .B1(new_n754), .B2(new_n700), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G2072), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n716), .A2(new_n722), .A3(new_n742), .A4(new_n756), .ZN(new_n757));
  OAI22_X1  g332(.A1(new_n720), .A2(new_n721), .B1(new_n755), .B2(G2072), .ZN(new_n758));
  INV_X1    g333(.A(G16), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G21), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G168), .B2(new_n759), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(G1966), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n759), .A2(G5), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G301), .B2(G16), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  AOI22_X1  g342(.A1(G1966), .A2(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n700), .A2(G27), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G164), .B2(new_n700), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT99), .B(G2078), .Z(new_n771));
  OAI211_X1 g346(.A(new_n767), .B(new_n768), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  OR4_X1    g347(.A1(new_n711), .A2(new_n757), .A3(new_n758), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n714), .A2(new_n715), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n759), .A2(G20), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G299), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G1956), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT101), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n759), .A2(G4), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n617), .B2(new_n759), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT93), .B(G1348), .Z(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n783), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n759), .A2(G19), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n560), .B2(new_n759), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n792), .A2(G1341), .B1(new_n770), .B2(new_n771), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n793), .B1(G1341), .B2(new_n792), .C1(new_n781), .C2(new_n782), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n773), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT91), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n483), .A2(G119), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n487), .A2(G131), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n467), .A2(G107), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n800), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G25), .B(new_n804), .S(G29), .Z(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT35), .B(G1991), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n805), .B(new_n806), .Z(new_n807));
  AND2_X1   g382(.A1(new_n759), .A2(G24), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G290), .B2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT89), .B(G1986), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n807), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n759), .A2(G6), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G305), .B2(G16), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT32), .B(G1981), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT90), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n819), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT90), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n821), .A2(new_n822), .A3(new_n817), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n759), .A2(G23), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G288), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT33), .B(G1976), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(G1971), .ZN(new_n828));
  NOR2_X1   g403(.A1(G166), .A2(new_n759), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n759), .A2(G22), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OR3_X1    g406(.A1(new_n829), .A2(new_n828), .A3(new_n830), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n820), .A2(new_n823), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n813), .B1(new_n834), .B2(KEYINPUT34), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT34), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n823), .A2(new_n820), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT92), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n797), .A2(new_n798), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n839), .B1(new_n838), .B2(new_n840), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n799), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n838), .A2(new_n840), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT92), .ZN(new_n846));
  INV_X1    g421(.A(new_n799), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n847), .A3(new_n841), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n796), .B1(new_n844), .B2(new_n848), .ZN(G311));
  NAND2_X1  g424(.A1(new_n844), .A2(new_n848), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n795), .ZN(G150));
  NAND2_X1  g426(.A1(new_n544), .A2(G55), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(new_n526), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(new_n523), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT104), .B(G860), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n617), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT103), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n861), .B(new_n863), .ZN(new_n864));
  OAI221_X1 g439(.A(new_n852), .B1(new_n853), .B2(new_n526), .C1(new_n855), .C2(new_n523), .ZN(new_n865));
  OAI221_X1 g440(.A(new_n554), .B1(new_n555), .B2(new_n526), .C1(new_n552), .C2(KEYINPUT73), .ZN(new_n866));
  INV_X1    g441(.A(new_n558), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n557), .A2(new_n857), .A3(new_n558), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n864), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT39), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n858), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n860), .B1(new_n874), .B2(new_n875), .ZN(G145));
  XNOR2_X1  g451(.A(new_n707), .B(new_n730), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n878));
  INV_X1    g453(.A(G118), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(G2105), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n487), .A2(G142), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(KEYINPUT105), .Z(new_n882));
  AOI211_X1 g457(.A(new_n880), .B(new_n882), .C1(G130), .C2(new_n483), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n877), .B(new_n883), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n494), .A2(new_n496), .B1(new_n483), .B2(G126), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n513), .A2(new_n514), .ZN(new_n886));
  AOI211_X1 g461(.A(KEYINPUT69), .B(new_n500), .C1(new_n512), .C2(new_n506), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n754), .B(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n804), .B(new_n633), .Z(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n884), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G160), .B(new_n644), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(G162), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n892), .B2(new_n895), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(G395));
  XNOR2_X1  g476(.A(G305), .B(G290), .ZN(new_n902));
  XNOR2_X1  g477(.A(G303), .B(G288), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n902), .B(new_n903), .Z(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n870), .A2(KEYINPUT107), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n868), .A2(new_n869), .A3(new_n907), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n906), .A2(new_n623), .A3(new_n617), .A4(new_n908), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n868), .A2(new_n869), .A3(new_n907), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n907), .B1(new_n868), .B2(new_n869), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n628), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n604), .A2(new_n612), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(G299), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n604), .A2(new_n612), .A3(new_n577), .A4(new_n573), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT108), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n920));
  INV_X1    g495(.A(new_n918), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n913), .A2(new_n919), .A3(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n915), .A2(new_n917), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n909), .A2(new_n912), .A3(new_n927), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n924), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n926), .B1(new_n924), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n905), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n925), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n924), .A2(new_n926), .A3(new_n928), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n904), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(G868), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n857), .A2(G868), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(G295));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n941), .A3(new_n939), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n598), .B1(new_n931), .B2(new_n935), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT110), .B1(new_n943), .B2(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(G331));
  NAND3_X1  g520(.A1(G286), .A2(G301), .A3(KEYINPUT112), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n547), .A2(new_n545), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT112), .B1(new_n947), .B2(new_n542), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n543), .A2(new_n949), .A3(new_n545), .A4(new_n547), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n950), .A3(G168), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n946), .A2(new_n951), .A3(new_n868), .A4(new_n869), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT114), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n946), .A2(new_n951), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n870), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(new_n927), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n923), .A2(new_n919), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n952), .A2(KEYINPUT113), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n952), .A2(KEYINPUT113), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n958), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n904), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n905), .B(new_n958), .C1(new_n959), .C2(new_n962), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n897), .A4(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n967), .A2(KEYINPUT44), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n921), .A2(new_n922), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n970));
  OR3_X1    g545(.A1(new_n954), .A2(new_n870), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n952), .A2(new_n970), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n955), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n960), .A2(new_n961), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n969), .A2(new_n973), .B1(new_n974), .B2(new_n957), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n966), .B(new_n897), .C1(new_n905), .C2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n976), .A2(new_n977), .A3(KEYINPUT43), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n977), .B1(new_n976), .B2(KEYINPUT43), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n968), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n981));
  NOR2_X1   g556(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n974), .A2(new_n955), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n923), .A2(new_n919), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n983), .A2(new_n984), .B1(new_n953), .B2(new_n957), .ZN(new_n985));
  AOI21_X1  g560(.A(G37), .B1(new_n985), .B2(new_n905), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n965), .B1(new_n986), .B2(new_n964), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n981), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n980), .A2(new_n988), .ZN(G397));
  AOI21_X1  g564(.A(KEYINPUT120), .B1(new_n571), .B2(new_n572), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(KEYINPUT57), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(G299), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(G164), .B2(G1384), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT118), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n996), .B(new_n993), .C1(G164), .C2(G1384), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n993), .A2(G1384), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n476), .A2(G40), .A3(new_n479), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT66), .B1(new_n472), .B2(G2105), .ZN(new_n1001));
  AOI211_X1 g576(.A(new_n462), .B(new_n467), .C1(new_n471), .C2(new_n463), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT116), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n474), .A2(new_n1005), .A3(new_n1000), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n888), .A2(new_n998), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT56), .B(G2072), .Z(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(KEYINPUT121), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n995), .A2(new_n997), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  INV_X1    g588(.A(G1384), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n888), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n779), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n992), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1348), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1005), .B1(new_n474), .B2(new_n1000), .ZN(new_n1021));
  AOI211_X1 g596(.A(KEYINPUT116), .B(new_n999), .C1(new_n468), .C2(new_n473), .ZN(new_n1022));
  OAI22_X1  g597(.A1(G164), .A2(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1013), .B1(new_n888), .B2(new_n1014), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1019), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G164), .A2(G1384), .ZN(new_n1026));
  INV_X1    g601(.A(G2067), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(new_n1027), .A3(new_n1012), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n914), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1010), .A2(new_n1017), .A3(new_n992), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1018), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1996), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n995), .A2(new_n1032), .A3(new_n997), .A4(new_n1007), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1026), .A2(new_n1012), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT58), .B(G1341), .Z(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n560), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT123), .B1(new_n1039), .B2(KEYINPUT59), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n914), .A2(KEYINPUT60), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1025), .A2(new_n1028), .A3(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1025), .A2(new_n914), .A3(new_n1028), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT60), .B1(new_n1044), .B2(new_n1029), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1030), .A2(KEYINPUT61), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1040), .B1(KEYINPUT123), .B2(KEYINPUT59), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1037), .A2(new_n560), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT61), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1010), .A2(new_n1017), .A3(new_n1050), .A4(new_n992), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1047), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1031), .B1(new_n1046), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT119), .B(G2084), .Z(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1023), .A2(new_n1024), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1966), .B1(new_n1007), .B2(new_n994), .ZN(new_n1057));
  OAI21_X1  g632(.A(G8), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G286), .A2(G8), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(KEYINPUT51), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n1061));
  INV_X1    g636(.A(G1966), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n888), .A2(new_n998), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1012), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT45), .B1(new_n888), .B2(new_n1014), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1011), .A2(new_n1015), .A3(new_n1012), .A4(new_n1054), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1061), .B(G8), .C1(new_n1068), .C2(G286), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1059), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(KEYINPUT124), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n1072));
  AOI211_X1 g647(.A(new_n1072), .B(new_n1059), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1060), .B(new_n1069), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n995), .A2(new_n997), .A3(new_n1007), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(G2078), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1075), .A2(G2078), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1078), .A2(new_n1079), .B1(new_n1016), .B2(new_n765), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g656(.A(G301), .B(KEYINPUT54), .Z(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1079), .B1(new_n466), .B2(new_n467), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(new_n999), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1063), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1084), .B1(new_n1087), .B2(new_n1065), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n765), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n994), .A2(new_n1063), .A3(KEYINPUT125), .A4(new_n1086), .ZN(new_n1090));
  AND4_X1   g665(.A1(new_n1082), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1081), .A2(new_n1083), .B1(new_n1091), .B2(new_n1077), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1074), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G303), .A2(G8), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT55), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1076), .A2(new_n828), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1023), .A2(new_n1024), .A3(G2090), .ZN(new_n1098));
  OAI211_X1 g673(.A(G8), .B(new_n1096), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1076), .B2(new_n828), .ZN(new_n1100));
  INV_X1    g675(.A(G8), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1095), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G288), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G1976), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1034), .A2(G8), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT52), .ZN(new_n1106));
  INV_X1    g681(.A(G1981), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n588), .B(new_n1107), .C1(new_n592), .C2(new_n593), .ZN(new_n1108));
  INV_X1    g683(.A(new_n591), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n588), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n1110), .B2(new_n1107), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT49), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1108), .B(KEYINPUT49), .C1(new_n1110), .C2(new_n1107), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1113), .A2(G8), .A3(new_n1034), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(G1976), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT52), .B1(G288), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1034), .A2(G8), .A3(new_n1104), .A4(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1106), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1099), .A2(new_n1102), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1053), .A2(new_n1093), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(G8), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1119), .B1(new_n1123), .B2(new_n1095), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1058), .A2(G286), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(KEYINPUT63), .A3(new_n1099), .A4(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1099), .A2(new_n1102), .A3(new_n1120), .A4(new_n1125), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1074), .A2(KEYINPUT62), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1070), .B(KEYINPUT124), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1132), .A2(new_n1133), .A3(new_n1060), .A4(new_n1069), .ZN(new_n1134));
  AOI21_X1  g709(.A(G301), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1131), .A2(new_n1134), .A3(new_n1121), .A4(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1099), .A2(new_n1119), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1034), .A2(G8), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1115), .A2(new_n1116), .A3(new_n1103), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(new_n1108), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1122), .A2(new_n1130), .A3(new_n1136), .A4(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n729), .B(new_n1027), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT117), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n707), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1032), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1065), .A2(new_n1012), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(new_n1032), .A3(new_n707), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n804), .A2(new_n806), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n804), .A2(new_n806), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1147), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1148), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(G290), .B(G1986), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1147), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1142), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1147), .A2(new_n1032), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT46), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT47), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1151), .B(KEYINPUT126), .ZN(new_n1163));
  OAI22_X1  g738(.A1(new_n1162), .A2(new_n1163), .B1(G2067), .B2(new_n729), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1147), .ZN(new_n1165));
  NOR2_X1   g740(.A1(G290), .A2(G1986), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1147), .A2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT48), .Z(new_n1168));
  OAI211_X1 g743(.A(new_n1161), .B(new_n1165), .C1(new_n1153), .C2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1156), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g746(.A1(new_n982), .A2(new_n987), .ZN(new_n1173));
  NOR3_X1   g747(.A1(G229), .A2(new_n460), .A3(G227), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n663), .A2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g749(.A1(new_n1173), .A2(new_n899), .A3(new_n1175), .ZN(G308));
  NOR2_X1   g750(.A1(new_n899), .A2(new_n1175), .ZN(new_n1177));
  OAI21_X1  g751(.A(new_n1177), .B1(new_n987), .B2(new_n982), .ZN(G225));
endmodule


