//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(G148gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G141gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT78), .B(G148gat), .ZN(new_n205));
  INV_X1    g004(.A(G141gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n210), .B2(KEYINPUT2), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n206), .A2(G148gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n203), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n208), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n207), .A2(new_n211), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT79), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G141gat), .B(G148gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n216), .B1(new_n220), .B2(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n202), .A2(KEYINPUT78), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT78), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G148gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n203), .B1(new_n225), .B2(G141gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n215), .B1(new_n212), .B2(new_n209), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n221), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT79), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n229), .A3(KEYINPUT3), .ZN(new_n230));
  XOR2_X1   g029(.A(G113gat), .B(G120gat), .Z(new_n231));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n232));
  INV_X1    g031(.A(G134gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G127gat), .ZN(new_n234));
  INV_X1    g033(.A(G127gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G134gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n231), .A2(new_n232), .A3(new_n234), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n236), .ZN(new_n238));
  XNOR2_X1  g037(.A(G113gat), .B(G120gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(KEYINPUT1), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n221), .B(new_n218), .C1(new_n226), .C2(new_n227), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n219), .A2(new_n230), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n237), .A2(new_n240), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n217), .A3(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT4), .B1(new_n228), .B2(new_n241), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n243), .A2(new_n244), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT5), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n228), .B(new_n241), .ZN(new_n252));
  INV_X1    g051(.A(new_n244), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT80), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT80), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n250), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n250), .A2(KEYINPUT5), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n261));
  XNOR2_X1  g060(.A(G1gat), .B(G29gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G57gat), .B(G85gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT6), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n265), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n256), .A2(new_n259), .A3(new_n267), .A4(new_n258), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n260), .A2(KEYINPUT6), .A3(new_n265), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G8gat), .B(G36gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(G64gat), .B(G92gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G226gat), .ZN(new_n275));
  INV_X1    g074(.A(G233gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(KEYINPUT29), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n283));
  NAND3_X1  g082(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT24), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n283), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G183gat), .ZN(new_n289));
  INV_X1    g088(.A(G190gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G169gat), .ZN(new_n294));
  INV_X1    g093(.A(G176gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT23), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(G169gat), .B2(G176gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT25), .A4(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n281), .B1(new_n293), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n284), .A2(new_n283), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n291), .B(new_n288), .C1(new_n302), .C2(new_n282), .ZN(new_n303));
  INV_X1    g102(.A(new_n300), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT67), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT64), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n307), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n286), .A2(new_n287), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n308), .A2(new_n309), .A3(new_n291), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n284), .A2(KEYINPUT64), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n310), .A2(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT65), .A4(new_n299), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT25), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n280), .B1(new_n306), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n313), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n311), .A2(new_n308), .A3(new_n309), .A4(new_n291), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n322), .A2(KEYINPUT68), .A3(new_n301), .A4(new_n305), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(KEYINPUT27), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT27), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(KEYINPUT69), .ZN(new_n329));
  OAI211_X1 g128(.A(KEYINPUT70), .B(G183gat), .C1(new_n327), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n290), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n332), .B1(KEYINPUT27), .B2(new_n289), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n334));
  AOI21_X1  g133(.A(new_n333), .B1(new_n334), .B2(G183gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n325), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT28), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT70), .B1(new_n328), .B2(G183gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(new_n289), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n340), .A2(KEYINPUT71), .A3(new_n330), .A4(new_n290), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n336), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT27), .B(G183gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(KEYINPUT28), .A3(new_n290), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT72), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NOR3_X1   g146(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n286), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n279), .B1(new_n324), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n352), .B1(new_n342), .B2(new_n346), .ZN(new_n356));
  INV_X1    g155(.A(new_n277), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n306), .A2(new_n316), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n360));
  NOR2_X1   g159(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n361));
  INV_X1    g160(.A(G211gat), .ZN(new_n362));
  INV_X1    g161(.A(G218gat), .ZN(new_n363));
  OAI22_X1  g162(.A1(new_n360), .A2(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G197gat), .B(G204gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n367), .A3(new_n365), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n355), .A2(new_n359), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n371), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n324), .A2(new_n354), .A3(new_n277), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n293), .A2(new_n281), .A3(new_n300), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT67), .B1(new_n303), .B2(new_n304), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n322), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n340), .A2(new_n290), .A3(new_n330), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT28), .B1(new_n379), .B2(new_n325), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n345), .B1(new_n380), .B2(new_n341), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n378), .B1(new_n381), .B2(new_n352), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n278), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n373), .B1(new_n374), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n274), .B1(new_n372), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n374), .A2(new_n383), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n371), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n354), .A2(new_n277), .A3(new_n378), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n356), .B1(new_n317), .B2(new_n323), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n373), .B(new_n388), .C1(new_n389), .C2(new_n279), .ZN(new_n390));
  INV_X1    g189(.A(new_n274), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n385), .A2(new_n392), .A3(KEYINPUT30), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT30), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n387), .A2(new_n394), .A3(new_n390), .A4(new_n391), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n271), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT68), .B1(new_n377), .B2(new_n322), .ZN(new_n400));
  AND4_X1   g199(.A1(KEYINPUT68), .A2(new_n322), .A3(new_n301), .A4(new_n305), .ZN(new_n401));
  OAI22_X1  g200(.A1(new_n400), .A2(new_n401), .B1(new_n381), .B2(new_n352), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n241), .ZN(new_n403));
  INV_X1    g202(.A(G227gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n404), .A2(new_n276), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n324), .A2(new_n354), .A3(new_n245), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n408), .A2(KEYINPUT34), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(KEYINPUT34), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n324), .A2(new_n354), .A3(new_n245), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n245), .B1(new_n324), .B2(new_n354), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n405), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G15gat), .B(G43gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(G71gat), .B(G99gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  NAND4_X1  g216(.A1(new_n414), .A2(KEYINPUT32), .A3(KEYINPUT33), .A4(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT73), .ZN(new_n419));
  INV_X1    g218(.A(new_n417), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n420), .B1(new_n414), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n418), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n403), .A2(new_n407), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n424), .B1(new_n425), .B2(new_n405), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n422), .B2(KEYINPUT73), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n411), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n406), .B1(new_n403), .B2(new_n407), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n419), .B(new_n417), .C1(new_n429), .C2(KEYINPUT33), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n417), .A2(KEYINPUT33), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n429), .A2(new_n424), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(KEYINPUT73), .B(new_n417), .C1(new_n429), .C2(KEYINPUT33), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n414), .A2(KEYINPUT32), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n433), .A2(new_n436), .A3(new_n410), .A4(new_n409), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n428), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n364), .A2(new_n367), .A3(new_n365), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n367), .B1(new_n364), .B2(new_n365), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n217), .B1(new_n442), .B2(new_n218), .ZN(new_n443));
  OAI211_X1 g242(.A(G228gat), .B(G233gat), .C1(new_n443), .C2(KEYINPUT83), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n371), .B1(new_n439), .B2(new_n242), .ZN(new_n445));
  OAI21_X1  g244(.A(G22gat), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT29), .B1(new_n369), .B2(new_n370), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n228), .B1(new_n447), .B2(KEYINPUT3), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n242), .A2(new_n439), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n373), .ZN(new_n450));
  INV_X1    g249(.A(G22gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  XOR2_X1   g251(.A(G78gat), .B(G106gat), .Z(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n446), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n454), .B1(new_n446), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT31), .B(G50gat), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n458), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n446), .A2(new_n452), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n453), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n462), .B2(new_n455), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n444), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n458), .B1(new_n456), .B2(new_n457), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n460), .A3(new_n455), .ZN(new_n466));
  INV_X1    g265(.A(new_n444), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(KEYINPUT35), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n271), .A2(new_n396), .A3(KEYINPUT87), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n399), .A2(new_n438), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n260), .A2(new_n265), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT82), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .A4(new_n268), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n270), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n266), .B2(new_n268), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n396), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT74), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n433), .B2(new_n436), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n411), .B1(new_n482), .B2(KEYINPUT75), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT74), .B1(new_n411), .B2(KEYINPUT75), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n436), .A3(new_n433), .ZN(new_n485));
  AOI211_X1 g284(.A(new_n480), .B(new_n470), .C1(new_n483), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT35), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n473), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n464), .A2(KEYINPUT84), .A3(new_n468), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT84), .B1(new_n464), .B2(new_n468), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n269), .A2(KEYINPUT82), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n492), .A2(new_n270), .A3(new_n477), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n493), .B2(new_n396), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT85), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n244), .B1(new_n243), .B2(new_n249), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT39), .B1(new_n252), .B2(new_n253), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT39), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n265), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  AOI211_X1 g299(.A(new_n495), .B(KEYINPUT40), .C1(new_n498), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n243), .A2(new_n249), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(new_n499), .A3(new_n253), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n503), .B(new_n267), .C1(new_n496), .C2(new_n497), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT85), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n503), .A2(new_n267), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n496), .A2(new_n497), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n265), .A2(new_n260), .B1(new_n510), .B2(KEYINPUT40), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n393), .A2(new_n507), .A3(new_n395), .A4(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT86), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT37), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n387), .A2(new_n514), .A3(new_n390), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n386), .A2(new_n373), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n371), .B(new_n388), .C1(new_n389), .C2(new_n279), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT37), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT38), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n515), .A2(new_n518), .A3(new_n519), .A4(new_n274), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n520), .A2(new_n269), .A3(new_n270), .A4(new_n392), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n515), .A2(new_n274), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT37), .B1(new_n372), .B2(new_n384), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT38), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n470), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n494), .B1(new_n513), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n428), .A2(new_n529), .A3(new_n437), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT76), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n428), .A2(new_n437), .A3(KEYINPUT76), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n529), .B1(new_n483), .B2(new_n485), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n528), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n488), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G1gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT16), .ZN(new_n539));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540));
  MUX2_X1   g339(.A(new_n538), .B(new_n539), .S(new_n540), .Z(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT93), .B(G8gat), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n543), .A2(new_n544), .B1(G8gat), .B2(new_n541), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT21), .ZN(new_n548));
  XOR2_X1   g347(.A(G57gat), .B(G64gat), .Z(new_n549));
  INV_X1    g348(.A(KEYINPUT9), .ZN(new_n550));
  INV_X1    g349(.A(G71gat), .ZN(new_n551));
  INV_X1    g350(.A(G78gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G71gat), .B(G78gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n549), .A2(new_n553), .B1(new_n554), .B2(KEYINPUT96), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(KEYINPUT96), .B2(new_n554), .ZN(new_n556));
  AND3_X1   g355(.A1(KEYINPUT97), .A2(KEYINPUT98), .A3(G57gat), .ZN(new_n557));
  OAI21_X1  g356(.A(G64gat), .B1(KEYINPUT97), .B2(G57gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(KEYINPUT98), .A2(G57gat), .ZN(new_n559));
  OAI22_X1  g358(.A1(new_n557), .A2(new_n558), .B1(G64gat), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n553), .B(new_n554), .C1(new_n560), .C2(KEYINPUT99), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n560), .A2(KEYINPUT99), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n556), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n547), .B1(new_n548), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n548), .ZN(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n566), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G183gat), .B(G211gat), .Z(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n570), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT103), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT104), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(G29gat), .A2(G36gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT14), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT91), .ZN(new_n588));
  XNOR2_X1  g387(.A(G43gat), .B(G50gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT90), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT15), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n589), .A2(new_n590), .A3(KEYINPUT15), .ZN(new_n592));
  XOR2_X1   g391(.A(KEYINPUT89), .B(G29gat), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(G36gat), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n588), .A2(new_n591), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n587), .A2(KEYINPUT88), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n594), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n587), .A2(KEYINPUT88), .ZN(new_n598));
  OAI211_X1 g397(.A(KEYINPUT15), .B(new_n589), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  INV_X1    g400(.A(G85gat), .ZN(new_n602));
  INV_X1    g401(.A(G92gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(KEYINPUT8), .A2(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n602), .B2(new_n603), .ZN(new_n606));
  NAND3_X1  g405(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G99gat), .B(G106gat), .Z(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  AOI21_X1  g409(.A(new_n585), .B1(new_n600), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT102), .ZN(new_n612));
  INV_X1    g411(.A(new_n600), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT17), .ZN(new_n614));
  INV_X1    g413(.A(new_n610), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G190gat), .B(G218gat), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n580), .A2(new_n581), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n619), .A2(new_n620), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n584), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n626), .A2(new_n622), .A3(new_n621), .A4(new_n583), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n577), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n545), .A2(new_n546), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n600), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n630), .A2(new_n600), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n635));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT13), .Z(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n637), .B1(new_n632), .B2(new_n633), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT95), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n547), .A2(new_n614), .A3(new_n617), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n642), .A2(new_n631), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(KEYINPUT18), .A3(new_n636), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n636), .A3(new_n631), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G113gat), .B(G141gat), .ZN(new_n648));
  INV_X1    g447(.A(G197gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT11), .B(G169gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT12), .Z(new_n653));
  NAND4_X1  g452(.A1(new_n641), .A2(new_n644), .A3(new_n647), .A4(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n638), .A2(new_n644), .A3(new_n647), .A4(new_n640), .ZN(new_n655));
  INV_X1    g454(.A(new_n653), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT106), .Z(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n608), .A2(new_n609), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(KEYINPUT105), .ZN(new_n664));
  OR3_X1    g463(.A1(new_n563), .A2(new_n610), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n610), .B1(new_n563), .B2(new_n664), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT10), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n615), .A2(new_n668), .A3(new_n563), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n662), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n665), .A2(new_n661), .A3(new_n666), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G120gat), .B(G148gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(G176gat), .B(G204gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n629), .A2(new_n659), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n537), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT107), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n537), .A2(new_n682), .A3(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n478), .A2(new_n479), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G1gat), .ZN(G1324gat));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n688));
  INV_X1    g487(.A(new_n396), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G8gat), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT16), .B(G8gat), .Z(new_n692));
  NAND3_X1  g491(.A1(new_n684), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n688), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n684), .A2(new_n689), .A3(new_n692), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(KEYINPUT42), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT108), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(G8gat), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n684), .B2(new_n689), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT42), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n700), .B(new_n701), .C1(KEYINPUT42), .C2(new_n695), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n697), .A2(new_n702), .ZN(G1325gat));
  NAND2_X1  g502(.A1(new_n684), .A2(new_n438), .ZN(new_n704));
  INV_X1    g503(.A(G15gat), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT109), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n704), .A2(KEYINPUT109), .A3(new_n705), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n534), .A2(new_n535), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n705), .ZN(new_n710));
  AOI211_X1 g509(.A(new_n706), .B(new_n707), .C1(new_n684), .C2(new_n710), .ZN(G1326gat));
  INV_X1    g510(.A(new_n491), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n684), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(new_n451), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  INV_X1    g515(.A(new_n628), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n537), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n678), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n576), .A2(new_n658), .A3(new_n719), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n721), .A2(new_n493), .A3(new_n593), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT45), .Z(new_n723));
  NOR2_X1   g522(.A1(new_n628), .A2(KEYINPUT44), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n488), .A2(KEYINPUT111), .A3(new_n536), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT111), .B1(new_n488), .B2(new_n536), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n718), .A2(KEYINPUT44), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n720), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n685), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(KEYINPUT112), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(KEYINPUT112), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n593), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n723), .B1(new_n731), .B2(new_n733), .ZN(G1328gat));
  OR3_X1    g533(.A1(new_n721), .A2(G36gat), .A3(new_n396), .ZN(new_n735));
  OR3_X1    g534(.A1(new_n735), .A2(KEYINPUT113), .A3(KEYINPUT46), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n729), .A2(new_n689), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G36gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(KEYINPUT46), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT113), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n736), .A2(new_n738), .A3(new_n739), .A4(new_n740), .ZN(G1329gat));
  INV_X1    g540(.A(new_n438), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n721), .A2(G43gat), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n729), .A2(new_n708), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(G43gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g545(.A1(new_n721), .A2(G50gat), .A3(new_n491), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(KEYINPUT114), .ZN(new_n748));
  INV_X1    g547(.A(G50gat), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n729), .B2(new_n712), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(KEYINPUT48), .A2(G50gat), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n729), .B2(new_n470), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n747), .B1(KEYINPUT114), .B2(KEYINPUT48), .ZN(new_n754));
  OAI22_X1  g553(.A1(new_n751), .A2(KEYINPUT48), .B1(new_n753), .B2(new_n754), .ZN(G1331gat));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n712), .A2(new_n480), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT86), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n512), .B(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n469), .B1(new_n521), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n757), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n532), .A2(new_n533), .ZN(new_n763));
  INV_X1    g562(.A(new_n535), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AND4_X1   g564(.A1(new_n438), .A2(new_n399), .A3(new_n471), .A4(new_n472), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n483), .A2(new_n485), .ZN(new_n767));
  INV_X1    g566(.A(new_n480), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n767), .A2(new_n768), .A3(new_n469), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n766), .B1(new_n769), .B2(KEYINPUT35), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n756), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n488), .A2(new_n536), .A3(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n629), .A2(new_n658), .A3(new_n719), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n493), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT97), .B(G57gat), .Z(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1332gat));
  INV_X1    g577(.A(new_n775), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT49), .B(G64gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n689), .A3(new_n780), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n775), .A2(new_n396), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(KEYINPUT115), .Z(G1333gat));
  NAND3_X1  g583(.A1(new_n779), .A2(KEYINPUT117), .A3(new_n438), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n775), .B2(new_n742), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n551), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n773), .A2(G71gat), .A3(new_n708), .A4(new_n774), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT116), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT50), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n788), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1334gat));
  NOR2_X1   g594(.A1(new_n775), .A2(new_n491), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(new_n552), .ZN(G1335gat));
  NOR2_X1   g596(.A1(new_n577), .A2(new_n658), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n717), .B(new_n798), .C1(new_n765), .C2(new_n770), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n628), .B1(new_n488), .B2(new_n536), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(KEYINPUT51), .A3(new_n798), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n719), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(G85gat), .B1(new_n804), .B2(new_n685), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n798), .A2(new_n678), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n727), .B2(new_n728), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n493), .A2(new_n602), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(G1336gat));
  AOI21_X1  g608(.A(new_n603), .B1(new_n807), .B2(new_n689), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n801), .A2(new_n803), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n799), .A2(KEYINPUT118), .A3(new_n800), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n719), .A2(G92gat), .A3(new_n396), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT52), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n803), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n814), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n818), .A2(KEYINPUT52), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n816), .B1(new_n810), .B2(new_n819), .ZN(G1337gat));
  INV_X1    g619(.A(new_n806), .ZN(new_n821));
  INV_X1    g620(.A(new_n724), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n771), .B2(new_n772), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n802), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G99gat), .B1(new_n826), .B2(new_n709), .ZN(new_n827));
  INV_X1    g626(.A(G99gat), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n804), .A2(new_n828), .A3(new_n438), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(G1338gat));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n831));
  INV_X1    g630(.A(G106gat), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n807), .B2(new_n470), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n469), .A2(G106gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n678), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n712), .B(new_n821), .C1(new_n823), .C2(new_n825), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(G106gat), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n834), .A2(new_n678), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n812), .A2(new_n813), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n836), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n831), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n832), .B1(new_n807), .B2(new_n712), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n812), .A2(new_n813), .A3(new_n841), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT53), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G106gat), .B1(new_n826), .B2(new_n469), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n836), .A3(new_n835), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(KEYINPUT119), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n844), .A2(new_n850), .ZN(G1339gat));
  NOR2_X1   g650(.A1(new_n493), .A2(new_n689), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  OR3_X1    g652(.A1(new_n667), .A2(new_n662), .A3(new_n669), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(KEYINPUT54), .A3(new_n670), .ZN(new_n855));
  XNOR2_X1  g654(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n670), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n857), .A2(KEYINPUT121), .A3(new_n675), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT121), .B1(new_n857), .B2(new_n675), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n676), .ZN(new_n863));
  INV_X1    g662(.A(new_n652), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n634), .A2(new_n637), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n643), .A2(new_n636), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n654), .A2(new_n625), .A3(new_n627), .A4(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT55), .B(new_n855), .C1(new_n858), .C2(new_n859), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OR3_X1    g669(.A1(new_n863), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n658), .A2(new_n676), .A3(new_n869), .A4(new_n862), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n654), .A2(new_n678), .A3(new_n867), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n871), .B(new_n872), .C1(new_n875), .C2(new_n717), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n717), .B1(new_n873), .B2(new_n874), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n863), .A2(new_n868), .A3(new_n870), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT122), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n876), .A2(new_n576), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n577), .A2(new_n628), .A3(new_n659), .A4(new_n719), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n853), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n882), .A2(new_n767), .A3(new_n469), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n659), .A2(G113gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n742), .A2(new_n712), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G113gat), .B1(new_n890), .B2(new_n659), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(G1340gat));
  NOR2_X1   g691(.A1(new_n719), .A2(G120gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n885), .A2(new_n886), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G120gat), .B1(new_n890), .B2(new_n719), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1341gat));
  NOR3_X1   g695(.A1(new_n890), .A2(new_n235), .A3(new_n576), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n883), .A2(new_n577), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n235), .ZN(G1342gat));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n233), .A3(new_n717), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n901));
  OAI21_X1  g700(.A(G134gat), .B1(new_n890), .B2(new_n628), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(KEYINPUT56), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G1343gat));
  AOI211_X1 g703(.A(KEYINPUT57), .B(new_n469), .C1(new_n880), .C2(new_n881), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n708), .A2(new_n853), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n576), .B1(new_n877), .B2(new_n878), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n491), .B1(new_n907), .B2(new_n881), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n905), .A2(new_n659), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n206), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n469), .B1(new_n880), .B2(new_n881), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n906), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n658), .A2(new_n206), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT58), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  OAI221_X1 g717(.A(new_n918), .B1(new_n914), .B2(new_n915), .C1(new_n911), .C2(new_n206), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1344gat));
  INV_X1    g719(.A(new_n914), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n225), .A3(new_n678), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n910), .ZN(new_n923));
  AOI211_X1 g722(.A(KEYINPUT59), .B(new_n225), .C1(new_n923), .C2(new_n678), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n925));
  AOI211_X1 g724(.A(new_n909), .B(new_n469), .C1(new_n880), .C2(new_n881), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n908), .A2(KEYINPUT57), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n678), .B(new_n906), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n925), .B1(new_n928), .B2(G148gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n922), .B1(new_n924), .B2(new_n929), .ZN(G1345gat));
  AOI21_X1  g729(.A(G155gat), .B1(new_n921), .B2(new_n577), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n577), .A2(G155gat), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n923), .B2(new_n932), .ZN(G1346gat));
  AOI21_X1  g732(.A(G162gat), .B1(new_n921), .B2(new_n717), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n717), .A2(G162gat), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n923), .B2(new_n935), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n685), .A2(new_n396), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n889), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n938), .B1(new_n880), .B2(new_n881), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n294), .B1(new_n939), .B2(new_n658), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT125), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n880), .A2(new_n881), .ZN(new_n942));
  AOI211_X1 g741(.A(new_n396), .B(new_n470), .C1(new_n483), .C2(new_n485), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n685), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n294), .A3(new_n658), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n941), .A2(new_n949), .ZN(G1348gat));
  AOI21_X1  g749(.A(G176gat), .B1(new_n948), .B2(new_n678), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n719), .A2(new_n295), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n951), .B1(new_n939), .B2(new_n952), .ZN(G1349gat));
  INV_X1    g752(.A(new_n343), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n947), .A2(new_n954), .A3(new_n576), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n289), .B1(new_n939), .B2(new_n577), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT60), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n957), .B(new_n958), .ZN(G1350gat));
  AOI21_X1  g758(.A(new_n290), .B1(new_n939), .B2(new_n717), .ZN(new_n960));
  XOR2_X1   g759(.A(new_n960), .B(KEYINPUT61), .Z(new_n961));
  NAND3_X1  g760(.A1(new_n948), .A2(new_n290), .A3(new_n717), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1351gat));
  NAND2_X1  g762(.A1(new_n709), .A2(new_n937), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n913), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(new_n649), .A3(new_n658), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n926), .A2(new_n927), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n968), .A2(new_n659), .A3(new_n964), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n967), .B1(new_n969), .B2(new_n649), .ZN(G1352gat));
  OAI21_X1  g769(.A(new_n678), .B1(new_n926), .B2(new_n927), .ZN(new_n971));
  OAI21_X1  g770(.A(G204gat), .B1(new_n971), .B2(new_n964), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n719), .A2(G204gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n913), .A2(new_n965), .A3(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n975), .B1(new_n974), .B2(KEYINPUT62), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n974), .A2(new_n975), .A3(KEYINPUT62), .ZN(new_n977));
  OAI221_X1 g776(.A(new_n972), .B1(KEYINPUT62), .B2(new_n974), .C1(new_n976), .C2(new_n977), .ZN(G1353gat));
  NAND3_X1  g777(.A1(new_n966), .A2(new_n362), .A3(new_n577), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n577), .B(new_n965), .C1(new_n926), .C2(new_n927), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n980), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n980), .B2(G211gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  AOI21_X1  g782(.A(G218gat), .B1(new_n966), .B2(new_n717), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n964), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n628), .A2(new_n363), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n986), .B(KEYINPUT127), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n984), .B1(new_n985), .B2(new_n987), .ZN(G1355gat));
endmodule


