//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n208), .B1(new_n202), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n207), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n207), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G20), .ZN(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n222), .B(new_n225), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n249), .B1(G1), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G116), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n226), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G283), .ZN(new_n256));
  INV_X1    g0056(.A(G20), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n256), .B(new_n257), .C1(G33), .C2(new_n218), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT75), .B(G116), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n254), .B(new_n258), .C1(new_n259), .C2(new_n257), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n252), .A2(KEYINPUT75), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT75), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G116), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n267), .A2(KEYINPUT20), .A3(new_n254), .A4(new_n258), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n255), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n248), .A2(G13), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n266), .A2(G20), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT5), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT74), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(KEYINPUT74), .A3(KEYINPUT5), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n276), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(G1), .A3(G13), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(new_n286), .B2(G270), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G264), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G257), .A2(G1698), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n288), .B(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G303), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n289), .A2(G33), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT66), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n285), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n227), .A2(KEYINPUT66), .A3(new_n284), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT79), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n285), .A2(new_n300), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT66), .B1(new_n227), .B2(new_n284), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT79), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(new_n294), .A4(new_n298), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n287), .A2(new_n304), .A3(new_n309), .ZN(new_n310));
  AND4_X1   g0110(.A1(KEYINPUT21), .A2(new_n273), .A3(G169), .A4(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n269), .B2(new_n272), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT21), .B1(new_n313), .B2(new_n310), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n273), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n310), .A2(G200), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n269), .A2(new_n272), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n287), .A2(new_n304), .A3(new_n309), .A4(G190), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n315), .A2(KEYINPUT80), .A3(new_n318), .A4(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n273), .A2(new_n310), .A3(G169), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT21), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n313), .A2(KEYINPUT21), .A3(new_n310), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n326), .A2(new_n322), .A3(new_n318), .A4(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT80), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT3), .B(G33), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n291), .A2(G222), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G223), .A2(G1698), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n307), .B(new_n335), .C1(G77), .C2(new_n332), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n282), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n285), .A2(new_n337), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n336), .B(new_n339), .C1(new_n209), .C2(new_n341), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n342), .A2(G179), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n257), .A2(G33), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT68), .ZN(new_n345));
  XOR2_X1   g0145(.A(KEYINPUT8), .B(G58), .Z(new_n346));
  NOR2_X1   g0146(.A1(G20), .A2(G33), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n345), .A2(new_n346), .B1(G150), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n203), .A2(G20), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n254), .B(KEYINPUT67), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n249), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n202), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT67), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n254), .B(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n257), .A2(G1), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(G50), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n352), .A2(new_n354), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n342), .A2(new_n312), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n343), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT9), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n342), .A2(G200), .ZN(new_n365));
  INV_X1    g0165(.A(G190), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n342), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n352), .A2(KEYINPUT9), .A3(new_n354), .A4(new_n359), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n364), .A2(new_n365), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT10), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n365), .B2(KEYINPUT69), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n371), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n362), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n340), .A2(G238), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G97), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(G226), .A2(G1698), .ZN(new_n378));
  INV_X1    g0178(.A(G232), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(G1698), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n377), .B1(new_n380), .B2(new_n332), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n375), .B(new_n339), .C1(new_n381), .C2(new_n303), .ZN(new_n382));
  XOR2_X1   g0182(.A(new_n382), .B(KEYINPUT13), .Z(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT14), .B1(new_n383), .B2(new_n312), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n382), .A2(KEYINPUT13), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(KEYINPUT13), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT14), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n388), .A3(G169), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT70), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n387), .B2(new_n316), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n385), .A2(KEYINPUT70), .A3(G179), .A4(new_n386), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n384), .A2(new_n389), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n257), .A2(G68), .ZN(new_n394));
  INV_X1    g0194(.A(new_n347), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(new_n202), .ZN(new_n396));
  AOI211_X1 g0196(.A(new_n394), .B(new_n396), .C1(new_n345), .C2(G77), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT11), .ZN(new_n398));
  OR3_X1    g0198(.A1(new_n397), .A2(new_n398), .A3(new_n356), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n397), .B2(new_n356), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n271), .A2(new_n394), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n401), .B(KEYINPUT12), .ZN(new_n402));
  INV_X1    g0202(.A(new_n254), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(G68), .A3(new_n358), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n399), .A2(new_n400), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n393), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n387), .A2(new_n366), .ZN(new_n407));
  INV_X1    g0207(.A(G200), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n385), .B2(new_n386), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n407), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G238), .A2(G1698), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n332), .B(new_n412), .C1(new_n379), .C2(G1698), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n307), .B(new_n413), .C1(G107), .C2(new_n332), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(new_n339), .C1(new_n211), .C2(new_n341), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(G179), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n250), .A2(G20), .ZN(new_n417));
  XOR2_X1   g0217(.A(KEYINPUT15), .B(G87), .Z(new_n418));
  AOI22_X1  g0218(.A1(new_n417), .A2(new_n418), .B1(new_n346), .B2(new_n347), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n257), .B2(new_n210), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n254), .B1(new_n210), .B2(new_n353), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n403), .A2(G77), .A3(new_n358), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n415), .A2(new_n312), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n416), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n374), .A2(new_n406), .A3(new_n411), .A4(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  INV_X1    g0227(.A(G68), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT72), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n289), .B2(G33), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n250), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n290), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(KEYINPUT7), .A3(new_n257), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT7), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT71), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT71), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT7), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n332), .B2(G20), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n428), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g0240(.A(G58), .B(G68), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n441), .A2(G20), .B1(G159), .B2(new_n347), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n427), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT7), .B1(new_n332), .B2(G20), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n288), .A2(new_n290), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n438), .A3(new_n257), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n447), .A3(G68), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(KEYINPUT16), .A3(new_n442), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(new_n254), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n209), .A2(G1698), .ZN(new_n451));
  OR2_X1    g0251(.A1(G223), .A2(G1698), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n332), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G87), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n307), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n285), .A2(G232), .A3(new_n337), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n456), .A2(new_n366), .A3(new_n458), .A4(new_n339), .ZN(new_n459));
  AOI211_X1 g0259(.A(new_n457), .B(new_n338), .C1(new_n455), .C2(new_n307), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(G200), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n356), .A2(new_n346), .A3(new_n358), .ZN(new_n462));
  INV_X1    g0262(.A(new_n346), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n353), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n450), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT17), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n449), .A2(new_n254), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n465), .B1(new_n470), .B2(new_n444), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(KEYINPUT17), .A3(new_n461), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n433), .A2(new_n439), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G68), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT16), .B1(new_n474), .B2(new_n442), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n449), .A2(new_n254), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n338), .B1(new_n455), .B2(new_n307), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(G179), .A3(new_n458), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n460), .B2(new_n312), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n477), .A2(KEYINPUT18), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT18), .B1(new_n477), .B2(new_n480), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n469), .B(new_n472), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n415), .A2(new_n366), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n415), .A2(G200), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(new_n421), .A4(new_n422), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n426), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n288), .A2(new_n290), .A3(new_n257), .A4(G87), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT22), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT22), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n332), .A2(new_n492), .A3(new_n257), .A4(G87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n259), .A2(new_n417), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n257), .A2(G107), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT23), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT81), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT81), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n499), .B(KEYINPUT23), .C1(new_n257), .C2(G107), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n498), .A2(new_n500), .B1(new_n497), .B2(new_n496), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n494), .A2(new_n495), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT24), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT24), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n494), .A2(new_n504), .A3(new_n501), .A4(new_n495), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n254), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n271), .A2(new_n496), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT25), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n508), .A2(KEYINPUT25), .ZN(new_n510));
  INV_X1    g0310(.A(new_n251), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n356), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n510), .B1(new_n513), .B2(G107), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n219), .A2(G1698), .ZN(new_n515));
  OR2_X1    g0315(.A1(G250), .A2(G1698), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n332), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G294), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n307), .ZN(new_n520));
  INV_X1    g0320(.A(new_n283), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n281), .A2(G264), .A3(new_n285), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n408), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n520), .A2(new_n366), .A3(new_n521), .A4(new_n522), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n507), .A2(new_n509), .A3(new_n514), .A4(new_n526), .ZN(new_n527));
  XOR2_X1   g0327(.A(new_n418), .B(KEYINPUT78), .Z(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(new_n512), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n332), .A2(new_n257), .A3(G68), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT76), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT19), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n218), .B2(new_n344), .ZN(new_n537));
  XNOR2_X1  g0337(.A(KEYINPUT76), .B(KEYINPUT19), .ZN(new_n538));
  AOI21_X1  g0338(.A(G20), .B1(new_n538), .B2(new_n377), .ZN(new_n539));
  NOR3_X1   g0339(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n531), .B(new_n537), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n254), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n418), .A2(new_n249), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT77), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT77), .ZN(new_n546));
  AOI211_X1 g0346(.A(new_n546), .B(new_n543), .C1(new_n541), .C2(new_n254), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n530), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n248), .A2(G45), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n282), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n285), .A2(G250), .A3(new_n549), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  OR2_X1    g0352(.A1(G238), .A2(G1698), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n211), .A2(G1698), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n332), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n259), .A2(G33), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI211_X1 g0357(.A(new_n550), .B(new_n552), .C1(new_n557), .C2(new_n307), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n316), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n307), .ZN(new_n560));
  INV_X1    g0360(.A(new_n550), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(new_n551), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n312), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n548), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n560), .A2(new_n366), .A3(new_n561), .A4(new_n551), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n558), .B2(G200), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n513), .A2(G87), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n567), .B(new_n568), .C1(new_n545), .C2(new_n547), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n527), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n288), .A2(new_n290), .A3(G244), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT4), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(G1698), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n332), .A2(G244), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n575), .A3(new_n256), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n332), .A2(G250), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n291), .B1(new_n577), .B2(KEYINPUT4), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n307), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n283), .B1(new_n286), .B2(G257), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(G190), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n249), .A2(G97), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n512), .B2(new_n218), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n473), .A2(G107), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n395), .A2(new_n210), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT6), .ZN(new_n588));
  INV_X1    g0388(.A(G107), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n218), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G97), .A2(G107), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(KEYINPUT6), .A3(G97), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n257), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n585), .A2(new_n587), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n584), .B1(new_n596), .B2(new_n254), .ZN(new_n597));
  INV_X1    g0397(.A(new_n580), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT73), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n579), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(KEYINPUT73), .B(new_n307), .C1(new_n576), .C2(new_n578), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n581), .B(new_n597), .C1(new_n602), .C2(new_n408), .ZN(new_n603));
  INV_X1    g0403(.A(new_n601), .ZN(new_n604));
  INV_X1    g0404(.A(new_n256), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n571), .B2(new_n572), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n572), .B1(new_n332), .B2(G250), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n575), .C1(new_n291), .C2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT73), .B1(new_n608), .B2(new_n307), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n316), .B(new_n580), .C1(new_n604), .C2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n584), .ZN(new_n611));
  AOI211_X1 g0411(.A(new_n586), .B(new_n594), .C1(new_n473), .C2(G107), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(new_n403), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n579), .A2(new_n580), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n312), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n610), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n603), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n570), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n507), .A2(new_n509), .A3(new_n514), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n523), .A2(G169), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT82), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n520), .A2(new_n522), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT83), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(G179), .A4(new_n521), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT83), .B1(new_n523), .B2(new_n316), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT82), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n523), .A2(new_n626), .A3(G169), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n621), .A2(new_n624), .A3(new_n625), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n619), .A2(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n331), .A2(new_n489), .A3(new_n618), .A4(new_n629), .ZN(G372));
  INV_X1    g0430(.A(new_n565), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  AOI22_X1  g0432(.A1(G97), .A2(new_n417), .B1(new_n533), .B2(new_n535), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n257), .B1(new_n536), .B2(new_n376), .ZN(new_n634));
  INV_X1    g0434(.A(new_n540), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n403), .B1(new_n636), .B2(new_n531), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n546), .B1(new_n637), .B2(new_n543), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n542), .A2(KEYINPUT77), .A3(new_n544), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n529), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n559), .A2(new_n563), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n569), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n632), .B1(new_n642), .B2(new_n616), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n610), .A2(new_n613), .A3(new_n615), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(KEYINPUT26), .A3(new_n565), .A4(new_n569), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n631), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n326), .A2(new_n318), .A3(new_n327), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n629), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n618), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n489), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT18), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n478), .A2(G179), .A3(new_n458), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n312), .B1(new_n478), .B2(new_n458), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n652), .B1(new_n471), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n477), .A2(KEYINPUT18), .A3(new_n480), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n425), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n411), .A2(new_n659), .B1(new_n393), .B2(new_n405), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n469), .A2(new_n472), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n372), .A2(new_n373), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n362), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n651), .A2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(G330), .ZN(new_n666));
  INV_X1    g0466(.A(G13), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G20), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n271), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT84), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(KEYINPUT84), .A3(KEYINPUT27), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n672), .A2(new_n673), .A3(G213), .A4(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n320), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n331), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n647), .A2(new_n680), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n666), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n619), .B1(new_n628), .B2(new_n677), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(KEYINPUT85), .A3(new_n527), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT85), .B1(new_n684), .B2(new_n527), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n686), .A2(new_n687), .B1(new_n629), .B2(new_n678), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n629), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n678), .ZN(new_n691));
  INV_X1    g0491(.A(new_n687), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n647), .A2(new_n677), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n685), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n689), .A2(new_n691), .A3(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n223), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n635), .A2(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n230), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n650), .A2(new_n678), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n527), .A2(new_n565), .A3(new_n569), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n603), .A2(KEYINPUT87), .A3(new_n616), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT87), .B1(new_n603), .B2(new_n616), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n706), .B(new_n648), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n646), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n678), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n331), .A2(new_n618), .A3(new_n629), .A4(new_n678), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n304), .A2(new_n309), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(G179), .A3(new_n287), .A4(new_n558), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n622), .A2(new_n579), .A3(new_n580), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n580), .B1(new_n604), .B2(new_n609), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n310), .A2(new_n523), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n558), .A2(G179), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AND4_X1   g0522(.A1(new_n520), .A2(new_n579), .A3(new_n522), .A4(new_n580), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n317), .A3(KEYINPUT30), .A4(new_n558), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n718), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n677), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g0527(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n728));
  NOR2_X1   g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n666), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n705), .A2(new_n712), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n702), .B1(new_n733), .B2(G1), .ZN(G364));
  NAND2_X1  g0534(.A1(new_n668), .A2(G45), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n698), .A2(G1), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n681), .A2(new_n682), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT89), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n257), .A2(new_n366), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n316), .A2(G200), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G322), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n366), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n408), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G283), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n446), .B1(new_n746), .B2(new_n747), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n316), .A2(new_n408), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G317), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT33), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n757), .A2(KEYINPUT33), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n749), .A2(new_n745), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G311), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n749), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G329), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n760), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n744), .A2(new_n754), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n753), .B(new_n768), .C1(G326), .C2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G294), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n257), .B1(new_n764), .B2(G190), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n773), .A2(KEYINPUT91), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(KEYINPUT91), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n744), .A2(new_n750), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n771), .B1(new_n772), .B2(new_n776), .C1(new_n295), .C2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n746), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n756), .A2(G68), .B1(new_n779), .B2(G58), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n210), .B2(new_n761), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT32), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n765), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n766), .A2(KEYINPUT32), .A3(G159), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n776), .A2(new_n218), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT90), .ZN(new_n788));
  INV_X1    g0588(.A(G87), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n332), .B1(new_n777), .B2(new_n789), .C1(new_n751), .C2(new_n589), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n786), .B(new_n791), .C1(new_n788), .C2(new_n790), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n769), .A2(new_n202), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n778), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n226), .B1(G20), .B2(new_n312), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n742), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n696), .A2(new_n332), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n229), .A2(new_n279), .A3(G50), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n797), .B(new_n798), .C1(new_n243), .C2(new_n279), .ZN(new_n799));
  NAND3_X1  g0599(.A1(G355), .A2(new_n223), .A3(new_n332), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(G116), .C2(new_n223), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n794), .A2(new_n795), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n736), .B1(new_n743), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n738), .A2(new_n666), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT88), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n666), .B2(new_n738), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n803), .B1(new_n806), .B2(new_n736), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT92), .ZN(G396));
  NAND2_X1  g0608(.A1(new_n423), .A2(new_n677), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n487), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n425), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n425), .A2(new_n677), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n740), .ZN(new_n815));
  INV_X1    g0615(.A(new_n736), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n756), .A2(G150), .B1(new_n779), .B2(G143), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n817), .B1(new_n818), .B2(new_n769), .C1(new_n783), .C2(new_n761), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT34), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n332), .B1(new_n765), .B2(new_n821), .C1(new_n428), .C2(new_n751), .ZN(new_n822));
  INV_X1    g0622(.A(new_n776), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(new_n823), .B2(G58), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n820), .B(new_n824), .C1(new_n202), .C2(new_n777), .ZN(new_n825));
  XOR2_X1   g0625(.A(KEYINPUT94), .B(G283), .Z(new_n826));
  AOI22_X1  g0626(.A1(new_n756), .A2(new_n826), .B1(new_n762), .B2(new_n259), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n827), .B1(new_n589), .B2(new_n777), .C1(new_n772), .C2(new_n746), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n751), .A2(new_n789), .ZN(new_n829));
  INV_X1    g0629(.A(G311), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n446), .B1(new_n769), .B2(new_n295), .C1(new_n830), .C2(new_n765), .ZN(new_n831));
  OR4_X1    g0631(.A1(new_n787), .A2(new_n828), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n795), .A2(new_n739), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT93), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n833), .A2(new_n795), .B1(new_n210), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n815), .A2(new_n816), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n677), .B1(new_n646), .B2(new_n649), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(new_n814), .ZN(new_n840));
  INV_X1    g0640(.A(new_n731), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n816), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT95), .Z(new_n843));
  OR2_X1    g0643(.A1(new_n840), .A2(new_n841), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n838), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  NOR2_X1   g0646(.A1(new_n406), .A2(new_n677), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT38), .ZN(new_n848));
  INV_X1    g0648(.A(new_n675), .ZN(new_n849));
  INV_X1    g0649(.A(new_n449), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT16), .B1(new_n448), .B2(new_n442), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n850), .A2(new_n851), .A3(new_n356), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n849), .B1(new_n852), .B2(new_n465), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT17), .B1(new_n471), .B2(new_n461), .ZN(new_n854));
  AND4_X1   g0654(.A1(KEYINPUT17), .A2(new_n450), .A3(new_n461), .A4(new_n466), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n853), .B1(new_n856), .B2(new_n658), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n655), .A2(new_n675), .B1(new_n450), .B2(new_n466), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n450), .A2(new_n461), .A3(new_n466), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n852), .A2(new_n465), .B1(new_n480), .B2(new_n849), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n467), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n860), .A2(new_n861), .B1(new_n863), .B2(KEYINPUT37), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n848), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n853), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n483), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n863), .A2(KEYINPUT37), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n477), .B1(new_n480), .B2(new_n849), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(new_n467), .A3(new_n861), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n867), .A2(KEYINPUT38), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n865), .A2(new_n872), .A3(KEYINPUT39), .ZN(new_n873));
  INV_X1    g0673(.A(new_n872), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n471), .A2(new_n675), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT98), .B1(new_n483), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n870), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n861), .B1(new_n869), .B2(new_n467), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n483), .A2(KEYINPUT98), .A3(new_n875), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n877), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n874), .B1(new_n883), .B2(new_n848), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n847), .B(new_n873), .C1(new_n884), .C2(KEYINPUT39), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n656), .A2(new_n657), .A3(new_n675), .ZN(new_n886));
  INV_X1    g0686(.A(new_n814), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n650), .A2(new_n678), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n813), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n865), .A2(new_n872), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n405), .A2(new_n677), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n406), .A2(new_n411), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n405), .B(new_n677), .C1(new_n393), .C2(new_n410), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n889), .A2(new_n890), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n885), .A2(new_n886), .A3(new_n895), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n489), .B1(new_n897), .B2(new_n704), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n664), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n896), .B(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT99), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n728), .B1(new_n725), .B2(new_n677), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n901), .B1(new_n904), .B2(new_n902), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n713), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n814), .B1(new_n892), .B2(new_n893), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n906), .A2(KEYINPUT40), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT98), .ZN(new_n909));
  INV_X1    g0709(.A(new_n875), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n909), .B(new_n910), .C1(new_n856), .C2(new_n658), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n911), .A2(new_n876), .A3(new_n880), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n872), .B1(new_n912), .B2(KEYINPUT38), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n890), .A2(new_n906), .A3(new_n907), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n908), .A2(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n489), .A2(new_n906), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(G330), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n900), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n248), .B2(new_n668), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n592), .A2(new_n593), .ZN(new_n922));
  OAI211_X1 g0722(.A(G20), .B(new_n227), .C1(new_n922), .C2(KEYINPUT35), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n252), .B(new_n923), .C1(KEYINPUT35), .C2(new_n922), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT36), .Z(new_n925));
  AOI211_X1 g0725(.A(new_n210), .B(new_n230), .C1(G58), .C2(G68), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT96), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(G50), .B2(new_n428), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(G1), .A3(new_n667), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n921), .A2(new_n925), .A3(new_n929), .ZN(G367));
  NAND2_X1  g0730(.A1(new_n613), .A2(new_n677), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n707), .B2(new_n708), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n644), .A2(new_n677), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT101), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n690), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n677), .B1(new_n937), .B2(new_n616), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n694), .A2(new_n932), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n939), .B(KEYINPUT42), .Z(new_n940));
  INV_X1    g0740(.A(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n638), .A2(new_n639), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n678), .B1(new_n942), .B2(new_n568), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n631), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n642), .B2(new_n943), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n938), .A2(new_n940), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n935), .A2(new_n689), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n941), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT100), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n948), .B(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n947), .B(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n697), .B(KEYINPUT41), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n694), .A2(new_n691), .A3(new_n934), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT45), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n694), .A2(new_n691), .ZN(new_n958));
  INV_X1    g0758(.A(new_n934), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT44), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT44), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n958), .A2(new_n962), .A3(new_n959), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n957), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n689), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT102), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n683), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n694), .B1(new_n688), .B2(new_n693), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(new_n732), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n957), .A2(new_n689), .A3(new_n961), .A4(new_n963), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT103), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n966), .A2(new_n971), .A3(KEYINPUT103), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n954), .B1(new_n977), .B2(new_n733), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n735), .A2(G1), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n952), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(G150), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n332), .B1(new_n746), .B2(new_n981), .C1(new_n755), .C2(new_n783), .ZN(new_n982));
  INV_X1    g0782(.A(new_n751), .ZN(new_n983));
  INV_X1    g0783(.A(new_n777), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n983), .A2(G77), .B1(new_n984), .B2(G58), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n818), .B2(new_n765), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n982), .B(new_n986), .C1(G143), .C2(new_n770), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n202), .B2(new_n761), .C1(new_n428), .C2(new_n776), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n756), .A2(G294), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n762), .A2(new_n826), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n984), .A2(KEYINPUT46), .A3(G116), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n446), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n751), .A2(new_n218), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G311), .B2(new_n770), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n295), .B2(new_n746), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT46), .B1(new_n984), .B2(new_n259), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n992), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n589), .B2(new_n776), .C1(new_n757), .C2(new_n765), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n988), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT104), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT47), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n736), .B1(new_n1001), .B2(new_n795), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n418), .A2(new_n696), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n797), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n796), .B(new_n1003), .C1(new_n239), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n742), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1002), .B(new_n1005), .C1(new_n1006), .C2(new_n945), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n980), .A2(new_n1007), .ZN(G387));
  INV_X1    g0808(.A(new_n971), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n698), .B1(new_n970), .B2(new_n732), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n762), .A2(G303), .B1(new_n756), .B2(G311), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n757), .B2(new_n746), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(KEYINPUT105), .B(G322), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1013), .B1(new_n770), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT106), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1016), .A2(KEYINPUT48), .B1(new_n823), .B2(new_n826), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(KEYINPUT48), .B2(new_n1016), .C1(new_n772), .C2(new_n777), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT49), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n766), .A2(G326), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n332), .B1(new_n983), .B2(new_n259), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n463), .A2(new_n755), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n528), .A2(new_n776), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n777), .A2(new_n210), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n769), .A2(new_n783), .B1(new_n746), .B2(new_n202), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(G150), .C2(new_n766), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n446), .B(new_n993), .C1(G68), .C2(new_n762), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1024), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n797), .B1(new_n236), .B2(new_n279), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n699), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1034), .A2(new_n223), .A3(new_n332), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n428), .A2(new_n210), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n346), .A2(new_n202), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1034), .B1(new_n1038), .B2(KEYINPUT50), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n279), .C1(KEYINPUT50), .C2(new_n1038), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1036), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(G107), .B2(new_n223), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1032), .A2(new_n795), .B1(new_n796), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n816), .C1(new_n688), .C2(new_n1006), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n979), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1011), .B(new_n1044), .C1(new_n1045), .C2(new_n970), .ZN(G393));
  OAI221_X1 g0846(.A(new_n796), .B1(new_n218), .B2(new_n223), .C1(new_n246), .C2(new_n1004), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n446), .B1(new_n751), .B2(new_n589), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n755), .A2(new_n295), .B1(new_n761), .B2(new_n772), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n984), .C2(new_n826), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n766), .A2(new_n1014), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n823), .A2(new_n259), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n769), .A2(new_n757), .B1(new_n746), .B2(new_n830), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT52), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G50), .A2(new_n756), .B1(new_n766), .B2(G143), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n428), .B2(new_n777), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1057), .A2(new_n446), .A3(new_n829), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n769), .A2(new_n981), .B1(new_n746), .B2(new_n783), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT51), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(new_n210), .C2(new_n776), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n463), .A2(new_n761), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n736), .B1(new_n1063), .B2(new_n795), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1047), .B(new_n1064), .C1(new_n936), .C2(new_n1006), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT107), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n966), .A2(new_n1066), .A3(new_n972), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n972), .A2(new_n1066), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1065), .B1(new_n1069), .B2(new_n1045), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n1069), .A2(new_n1009), .B1(new_n975), .B2(new_n976), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1070), .B1(new_n1071), .B2(new_n697), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(G390));
  NAND2_X1  g0873(.A1(new_n984), .A2(G150), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT53), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n446), .B1(new_n1074), .B2(KEYINPUT53), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n766), .A2(G125), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n983), .A2(G50), .B1(new_n779), .B2(G132), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n776), .A2(new_n783), .B1(new_n818), .B2(new_n755), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT54), .B(G143), .Z(new_n1081));
  AOI21_X1  g0881(.A(new_n1080), .B1(new_n762), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT110), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1079), .B(new_n1083), .C1(G128), .C2(new_n770), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G294), .A2(new_n766), .B1(new_n770), .B2(G283), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n218), .B2(new_n761), .C1(new_n252), .C2(new_n746), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n776), .A2(new_n210), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n755), .A2(new_n589), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n446), .B1(new_n777), .B2(new_n789), .C1(new_n751), .C2(new_n428), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n795), .B1(new_n1084), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n835), .A2(new_n463), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n816), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT111), .ZN(new_n1094));
  OR2_X1    g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n873), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT39), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n913), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1095), .B1(new_n1098), .B2(new_n741), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT112), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n847), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n894), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n677), .B1(new_n646), .B2(new_n709), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n812), .B1(new_n1104), .B2(new_n811), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n913), .B(new_n1102), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n847), .B1(new_n889), .B2(new_n894), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1098), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n814), .A2(new_n666), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n906), .A2(new_n894), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT108), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n906), .A2(new_n1109), .A3(KEYINPUT108), .A4(new_n894), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1108), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n727), .A2(new_n730), .A3(new_n887), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1116), .A2(new_n1103), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1106), .B(new_n1117), .C1(new_n1098), .C2(new_n1107), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1115), .A2(new_n979), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1101), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n906), .A2(new_n1109), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1117), .B(new_n1105), .C1(new_n894), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1116), .A2(new_n1103), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1112), .A2(new_n1123), .A3(new_n1113), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n889), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n489), .A2(G330), .A3(new_n906), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n898), .A2(new_n664), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n873), .B1(new_n884), .B2(KEYINPUT39), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n812), .B1(new_n839), .B2(new_n887), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1102), .B1(new_n1132), .B2(new_n1103), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n883), .A2(new_n848), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n847), .B1(new_n1134), .B2(new_n872), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n710), .A2(new_n678), .A3(new_n811), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n894), .B1(new_n1136), .B2(new_n812), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1131), .A2(new_n1133), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1114), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1118), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1130), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1128), .B1(new_n1125), .B2(new_n1122), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n1118), .A3(new_n1115), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1141), .A2(new_n1143), .A3(new_n697), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(KEYINPUT109), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT109), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1141), .A2(new_n1143), .A3(new_n1146), .A4(new_n697), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1120), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(G378));
  INV_X1    g0949(.A(KEYINPUT55), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n374), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(KEYINPUT55), .B(new_n362), .C1(new_n372), .C2(new_n373), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n360), .A2(new_n849), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT56), .Z(new_n1156));
  NAND3_X1  g0956(.A1(new_n1152), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1156), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1159), .A3(new_n740), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n834), .A2(new_n202), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n983), .A2(G58), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n210), .B2(new_n777), .C1(new_n752), .C2(new_n765), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n755), .A2(new_n218), .B1(new_n746), .B2(new_n589), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n332), .B(new_n1164), .C1(G116), .C2(new_n770), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1165), .B(new_n277), .C1(new_n528), .C2(new_n761), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1163), .B(new_n1166), .C1(G68), .C2(new_n823), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT58), .Z(new_n1168));
  NOR2_X1   g0968(.A1(new_n776), .A2(new_n981), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n756), .A2(G132), .B1(new_n779), .B2(G128), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G125), .A2(new_n770), .B1(new_n984), .B2(new_n1081), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1169), .B(new_n1172), .C1(G137), .C2(new_n762), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT59), .ZN(new_n1174));
  AOI21_X1  g0974(.A(G41), .B1(new_n766), .B2(G124), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G33), .B1(new_n983), .B2(G159), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1168), .B(new_n1177), .C1(G50), .C2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n736), .B1(new_n1179), .B2(new_n795), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1160), .A2(new_n1161), .A3(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT113), .ZN(new_n1182));
  MUX2_X1   g0982(.A(new_n1116), .B(new_n1121), .S(new_n1103), .Z(new_n1183));
  AOI22_X1  g0983(.A1(new_n1183), .A2(new_n1105), .B1(new_n1124), .B2(new_n889), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1129), .B1(new_n1140), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n885), .A2(new_n886), .A3(new_n895), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n908), .A2(new_n913), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT114), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1157), .A2(new_n1159), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n914), .A2(new_n915), .ZN(new_n1190));
  AND4_X1   g0990(.A1(G330), .A2(new_n1187), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1189), .B1(new_n916), .B2(G330), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1186), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1189), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n890), .A2(new_n906), .A3(new_n907), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT40), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n1195), .A2(KEYINPUT40), .B1(new_n884), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1197), .B2(new_n666), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n916), .A2(G330), .A3(new_n1189), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n896), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1193), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n698), .B1(new_n1185), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1182), .B1(new_n1202), .B2(KEYINPUT57), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1200), .B(KEYINPUT117), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT115), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1198), .A2(new_n1205), .A3(new_n1199), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1186), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT116), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(KEYINPUT115), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1198), .A2(new_n1205), .A3(new_n1199), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(KEYINPUT116), .A3(new_n1186), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1204), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n698), .A2(KEYINPUT57), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n979), .B1(new_n1185), .B2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1203), .B1(new_n1215), .B2(new_n1217), .ZN(G375));
  NAND3_X1  g1018(.A1(new_n1122), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1130), .A2(new_n953), .A3(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1162), .A2(new_n332), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT119), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n761), .A2(new_n981), .B1(new_n769), .B2(new_n821), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n756), .A2(new_n1081), .B1(new_n766), .B2(G128), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n818), .B2(new_n746), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n202), .B2(new_n776), .C1(new_n783), .C2(new_n777), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n755), .A2(new_n266), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n446), .B1(new_n751), .B2(new_n210), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n769), .A2(new_n772), .B1(new_n746), .B2(new_n752), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(G107), .C2(new_n762), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n765), .A2(new_n295), .B1(new_n777), .B2(new_n218), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT118), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1026), .A2(new_n1231), .A3(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1227), .B1(new_n1228), .B2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT120), .Z(new_n1236));
  AOI21_X1  g1036(.A(new_n736), .B1(new_n1236), .B2(new_n795), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n835), .A2(new_n428), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1103), .A2(new_n739), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1184), .B2(new_n1045), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1220), .A2(new_n1242), .ZN(G381));
  AND2_X1   g1043(.A1(new_n1101), .A2(new_n1119), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1144), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(G375), .A2(G384), .A3(G381), .A4(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n980), .A2(new_n1072), .A3(new_n1007), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  OR2_X1    g1048(.A1(G396), .A2(G393), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1246), .A2(new_n1248), .A3(new_n1250), .ZN(G407));
  NAND2_X1  g1051(.A1(G407), .A2(G213), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1185), .A2(new_n1201), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(KEYINPUT57), .A3(new_n697), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1182), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT117), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1200), .B(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(KEYINPUT116), .B1(new_n1213), .B2(new_n1186), .ZN(new_n1259));
  AOI211_X1 g1059(.A(new_n1209), .B(new_n896), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1217), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1256), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1244), .A2(new_n1144), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n676), .A2(G213), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1264), .A3(new_n1266), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(KEYINPUT121), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1252), .A2(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(KEYINPUT122), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1219), .A2(new_n1271), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1125), .A2(new_n1122), .A3(new_n1128), .A4(KEYINPUT60), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1130), .A3(new_n697), .A4(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT123), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1122), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1142), .B1(new_n1277), .B2(KEYINPUT60), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n698), .B1(new_n1219), .B2(new_n1271), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(KEYINPUT123), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1281), .B2(new_n1242), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n845), .B(new_n1241), .C1(new_n1276), .C2(new_n1280), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(G375), .A2(new_n1148), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1185), .A2(new_n953), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1261), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1182), .B1(new_n1201), .B2(new_n979), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1245), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1265), .B(new_n1284), .C1(new_n1285), .C2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT62), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1266), .A2(G2897), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT123), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1242), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n845), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1281), .A2(G384), .A3(new_n1242), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1293), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1294), .A2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1289), .B1(new_n1215), .B2(new_n1286), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n1263), .A2(G378), .B1(new_n1303), .B2(new_n1264), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1302), .B1(new_n1304), .B2(new_n1266), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT61), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1289), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1261), .B2(new_n1287), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(G375), .A2(new_n1148), .B1(new_n1308), .B2(new_n1245), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n1265), .A4(new_n1284), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1292), .A2(new_n1305), .A3(new_n1306), .A4(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT125), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1072), .B1(new_n980), .B2(new_n1007), .ZN(new_n1314));
  XOR2_X1   g1114(.A(G396), .B(G393), .Z(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1248), .A2(new_n1314), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G387), .A2(G390), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1315), .B1(new_n1318), .B2(new_n1247), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1313), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1316), .B1(new_n1248), .B2(new_n1314), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1318), .A2(new_n1247), .A3(new_n1315), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(new_n1322), .A3(KEYINPUT125), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1320), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1312), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT124), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1326), .B1(new_n1304), .B2(new_n1266), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1309), .A2(KEYINPUT124), .A3(new_n1265), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1327), .A2(new_n1302), .A3(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT61), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1291), .A2(new_n1331), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1309), .A2(KEYINPUT63), .A3(new_n1265), .A4(new_n1284), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1329), .A2(new_n1330), .A3(new_n1332), .A4(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1325), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(KEYINPUT126), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT126), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1325), .A2(new_n1334), .A3(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1336), .A2(new_n1338), .ZN(G405));
  NAND2_X1  g1139(.A1(G375), .A2(new_n1264), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1340), .B1(new_n1148), .B2(G375), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(new_n1341), .B(new_n1284), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1343));
  OR3_X1    g1143(.A1(new_n1342), .A2(KEYINPUT127), .A3(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT127), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1346));
  AND3_X1   g1146(.A1(new_n1344), .A2(new_n1345), .A3(new_n1346), .ZN(G402));
endmodule


