//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  AND2_X1   g003(.A1(new_n189), .A2(G221), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT81), .Z(new_n191));
  INV_X1    g005(.A(KEYINPUT86), .ZN(new_n192));
  INV_X1    g006(.A(G469), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G110), .B(G140), .ZN(new_n195));
  INV_X1    g009(.A(G953), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n196), .A2(G227), .ZN(new_n197));
  XOR2_X1   g011(.A(new_n195), .B(new_n197), .Z(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT64), .B1(new_n199), .B2(G134), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G137), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n199), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT11), .B1(new_n199), .B2(G134), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT65), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n202), .B2(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n199), .A2(KEYINPUT11), .A3(G134), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n210), .A2(new_n200), .A3(new_n203), .A4(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n208), .A2(G131), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n212), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT66), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n208), .A2(new_n214), .A3(KEYINPUT66), .A4(G131), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT84), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(KEYINPUT84), .A3(new_n220), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G104), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G107), .ZN(new_n227));
  INV_X1    g041(.A(G107), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G104), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G101), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT3), .B1(new_n226), .B2(G107), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n228), .A3(G104), .ZN(new_n234));
  INV_X1    g048(.A(G101), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n232), .A2(new_n234), .A3(new_n235), .A4(new_n227), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n236), .A2(KEYINPUT82), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(KEYINPUT82), .ZN(new_n238));
  OAI211_X1 g052(.A(KEYINPUT10), .B(new_n231), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n240));
  INV_X1    g054(.A(G143), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G146), .ZN(new_n242));
  OR2_X1    g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  XNOR2_X1  g058(.A(G143), .B(G146), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(new_n240), .ZN(new_n246));
  INV_X1    g060(.A(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n242), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(G128), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n243), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  OR3_X1    g066(.A1(new_n239), .A2(new_n252), .A3(KEYINPUT83), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT83), .B1(new_n239), .B2(new_n252), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n232), .A2(new_n234), .A3(new_n227), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G101), .ZN(new_n256));
  OAI211_X1 g070(.A(KEYINPUT4), .B(new_n256), .C1(new_n237), .C2(new_n238), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n249), .A2(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n245), .A2(new_n244), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT0), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n245), .A2(KEYINPUT0), .A3(new_n244), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OR2_X1    g076(.A1(new_n256), .A2(KEYINPUT4), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n257), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT10), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n231), .B1(new_n237), .B2(new_n238), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n267));
  OAI22_X1  g081(.A1(new_n246), .A2(new_n250), .B1(new_n267), .B2(new_n242), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n265), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n253), .A2(new_n254), .A3(new_n264), .A4(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n198), .B1(new_n225), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n252), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(new_n266), .B2(new_n269), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n219), .A2(new_n220), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT85), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT12), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n274), .A2(new_n275), .A3(new_n276), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n223), .A2(new_n224), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n270), .A2(new_n264), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n254), .A4(new_n253), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n271), .A2(new_n275), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n198), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n188), .B(new_n194), .C1(new_n282), .C2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n192), .A2(new_n193), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n198), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n225), .A2(new_n271), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n281), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n285), .A2(new_n286), .A3(new_n198), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n193), .B1(new_n295), .B2(new_n188), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n191), .B1(new_n290), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G214), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(G119), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G116), .ZN(new_n300));
  INV_X1    g114(.A(G116), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G119), .ZN(new_n302));
  INV_X1    g116(.A(G113), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n303), .A2(KEYINPUT2), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(KEYINPUT2), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n300), .B(new_n302), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n300), .A2(new_n302), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT2), .B(G113), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n306), .A2(new_n309), .A3(KEYINPUT68), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT68), .B1(new_n306), .B2(new_n309), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n257), .A2(new_n312), .A3(new_n263), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n236), .A2(KEYINPUT82), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n236), .A2(KEYINPUT82), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n314), .A2(new_n315), .B1(G101), .B2(new_n230), .ZN(new_n316));
  INV_X1    g130(.A(new_n306), .ZN(new_n317));
  MUX2_X1   g131(.A(new_n300), .B(new_n307), .S(KEYINPUT5), .Z(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(G113), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g135(.A(G110), .B(G122), .Z(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n322), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n313), .A2(new_n324), .A3(new_n320), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(KEYINPUT6), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G125), .B1(new_n260), .B2(new_n261), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n243), .B(new_n328), .C1(new_n246), .C2(new_n250), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT87), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n329), .A2(new_n330), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n327), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT88), .B(G224), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n196), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n329), .A2(new_n330), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n331), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n327), .A3(new_n336), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n321), .A2(new_n343), .A3(new_n322), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n326), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT89), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n326), .A2(new_n342), .A3(KEYINPUT89), .A4(new_n344), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G210), .B1(G237), .B2(G902), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT90), .B1(new_n332), .B2(new_n333), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n339), .A2(new_n352), .A3(new_n331), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n353), .A3(new_n327), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n336), .A2(KEYINPUT7), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n316), .B(new_n319), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n322), .B(KEYINPUT8), .Z(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OR2_X1    g173(.A1(new_n337), .A2(KEYINPUT91), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT7), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n337), .B2(KEYINPUT91), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n340), .A2(new_n327), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n356), .A2(new_n325), .A3(new_n359), .A4(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n364), .A2(new_n188), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n349), .A2(new_n350), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n350), .B1(new_n349), .B2(new_n365), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n298), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G237), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n196), .A3(G214), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n370), .A2(new_n241), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n241), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n217), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT17), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n372), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G131), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n370), .B(G143), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n217), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT17), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT74), .ZN(new_n381));
  INV_X1    g195(.A(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G125), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n328), .A2(G140), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT73), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .A4(KEYINPUT16), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT16), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT73), .B1(new_n383), .B2(KEYINPUT16), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n381), .B1(new_n389), .B2(G146), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT16), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n391), .B(KEYINPUT73), .C1(KEYINPUT16), .C2(new_n383), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n247), .B1(new_n392), .B2(new_n386), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n389), .A2(KEYINPUT74), .A3(G146), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n374), .B(new_n380), .C1(new_n394), .C2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G113), .B(G122), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n226), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n373), .A2(KEYINPUT18), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT18), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n377), .B1(new_n401), .B2(new_n217), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n383), .A2(new_n384), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(G146), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n400), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n397), .A2(new_n399), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n399), .B1(new_n397), .B2(new_n405), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n188), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G475), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT20), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n375), .A2(G131), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT92), .B1(new_n411), .B2(new_n373), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n389), .A2(G146), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n403), .B(KEYINPUT19), .Z(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n247), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT92), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n376), .A2(new_n378), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n412), .A2(new_n413), .A3(new_n415), .A4(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n399), .B1(new_n418), .B2(new_n405), .ZN(new_n419));
  INV_X1    g233(.A(new_n405), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n392), .A2(new_n247), .A3(new_n386), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n413), .A2(new_n421), .A3(new_n381), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n411), .A2(new_n373), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n395), .A2(new_n422), .B1(new_n423), .B2(new_n379), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n420), .B1(new_n424), .B2(new_n374), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n419), .B1(new_n425), .B2(new_n399), .ZN(new_n426));
  NOR2_X1   g240(.A1(G475), .A2(G902), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT93), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n410), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n397), .A2(new_n399), .A3(new_n405), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n418), .A2(new_n405), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n430), .B1(new_n431), .B2(new_n399), .ZN(new_n432));
  INV_X1    g246(.A(new_n428), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(KEYINPUT20), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n409), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G128), .B(G143), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT13), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n241), .A2(G128), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n439), .A2(KEYINPUT13), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n438), .A2(G134), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(new_n202), .ZN(new_n442));
  INV_X1    g256(.A(G122), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G116), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n301), .A2(G122), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(new_n228), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n228), .B1(new_n444), .B2(new_n445), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n442), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT14), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n444), .A2(new_n445), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G107), .B1(new_n445), .B2(new_n450), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n244), .A2(G143), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n439), .A2(new_n454), .A3(new_n202), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n202), .B1(new_n439), .B2(new_n454), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI22_X1  g271(.A1(new_n441), .A2(new_n449), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT72), .B(G217), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n187), .A2(new_n196), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT94), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT94), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n187), .A2(new_n462), .A3(new_n196), .A4(new_n459), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT95), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n438), .A2(G134), .A3(new_n440), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n467), .B(new_n442), .C1(new_n448), .C2(new_n447), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n461), .A2(new_n463), .ZN(new_n469));
  OAI221_X1 g283(.A(new_n446), .B1(new_n455), .B2(new_n456), .C1(new_n451), .C2(new_n452), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n465), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n468), .A2(new_n469), .A3(new_n470), .A4(KEYINPUT95), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n188), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G478), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(KEYINPUT15), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n476), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n472), .A2(new_n188), .A3(new_n473), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT96), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n477), .A2(KEYINPUT96), .A3(new_n479), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(G234), .A2(G237), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(G952), .A3(new_n196), .ZN(new_n486));
  XOR2_X1   g300(.A(KEYINPUT21), .B(G898), .Z(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(G902), .A3(G953), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n436), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n297), .A2(new_n368), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n219), .A2(new_n262), .A3(new_n220), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n202), .A2(G137), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n199), .A2(G134), .ZN(new_n495));
  OAI21_X1  g309(.A(G131), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n251), .B(new_n496), .C1(G131), .C2(new_n212), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n493), .B1(new_n492), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n312), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n312), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n492), .A2(new_n501), .A3(new_n497), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n503));
  NAND3_X1  g317(.A1(new_n369), .A2(new_n196), .A3(G210), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT26), .B(G101), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n500), .A2(new_n502), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT31), .ZN(new_n509));
  INV_X1    g323(.A(new_n502), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT28), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n492), .A2(new_n497), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n312), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT28), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n502), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n511), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n507), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT31), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n500), .A2(new_n519), .A3(new_n502), .A4(new_n507), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n509), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n509), .A2(KEYINPUT70), .A3(new_n518), .A4(new_n520), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(G472), .A2(G902), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT32), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(KEYINPUT32), .A3(new_n526), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n513), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n510), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n511), .A2(new_n515), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n533), .B1(new_n534), .B2(new_n532), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT29), .A3(new_n507), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n500), .A2(new_n502), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n537), .A2(new_n507), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n516), .A2(new_n517), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n188), .B(new_n536), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n529), .A2(new_n530), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n299), .A2(G128), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n244), .A2(G119), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT24), .B(G110), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT23), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n299), .B2(G128), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n244), .A2(KEYINPUT23), .A3(G119), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n545), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G110), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n422), .A2(new_n395), .A3(new_n549), .A4(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G110), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n551), .A2(new_n552), .A3(new_n556), .A4(new_n545), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT75), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n547), .A2(new_n548), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n558), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n403), .A2(G146), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n389), .B2(G146), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n562), .A2(new_n564), .A3(KEYINPUT76), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT76), .B1(new_n562), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n555), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT77), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n196), .A2(G221), .A3(G234), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT22), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(G137), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n555), .B(KEYINPUT77), .C1(new_n565), .C2(new_n566), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n567), .A2(new_n572), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n459), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(G234), .B2(new_n188), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G902), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n581), .B(KEYINPUT79), .Z(new_n582));
  NAND2_X1  g396(.A1(new_n577), .A2(new_n188), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT78), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT25), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n577), .A2(new_n584), .A3(new_n585), .A4(new_n188), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n579), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n544), .A2(KEYINPUT80), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT80), .B1(new_n544), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n491), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  AOI21_X1  g409(.A(G902), .B1(new_n523), .B2(new_n524), .ZN(new_n596));
  INV_X1    g410(.A(G472), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(KEYINPUT97), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n596), .B(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n297), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n591), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n602));
  INV_X1    g416(.A(new_n474), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n602), .B1(new_n603), .B2(G478), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n474), .A2(KEYINPUT99), .A3(new_n475), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n472), .A2(new_n607), .A3(new_n473), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n465), .A2(KEYINPUT33), .A3(new_n471), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(G478), .A3(new_n188), .A4(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n610), .A2(KEYINPUT98), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(KEYINPUT98), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n435), .ZN(new_n614));
  INV_X1    g428(.A(new_n298), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n349), .A2(new_n365), .ZN(new_n616));
  INV_X1    g430(.A(new_n350), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n349), .A2(new_n350), .A3(new_n365), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n615), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n489), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n601), .A2(new_n614), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT34), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(new_n484), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n436), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n601), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT35), .B(G107), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  AND2_X1   g443(.A1(new_n569), .A2(new_n574), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n580), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n589), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n599), .A2(new_n637), .A3(new_n491), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT37), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n556), .ZN(G12));
  NOR2_X1   g454(.A1(new_n297), .A2(new_n368), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n488), .A2(G900), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n486), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n625), .A2(new_n436), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT101), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n544), .A2(new_n641), .A3(new_n637), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  NAND2_X1  g461(.A1(new_n618), .A2(new_n619), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT38), .Z(new_n649));
  XOR2_X1   g463(.A(new_n643), .B(KEYINPUT39), .Z(new_n650));
  NOR2_X1   g464(.A1(new_n297), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n537), .A2(new_n517), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n532), .B(new_n502), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n655), .B(new_n188), .C1(new_n507), .C2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G472), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n529), .A2(new_n530), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n615), .B1(new_n482), .B2(new_n483), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n435), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n635), .B1(new_n651), .B2(new_n652), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n654), .A2(new_n659), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G143), .ZN(G45));
  NAND3_X1  g478(.A1(new_n613), .A2(new_n435), .A3(new_n643), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT103), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n613), .A2(new_n435), .A3(new_n667), .A4(new_n643), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n544), .A2(new_n641), .A3(new_n637), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G146), .ZN(G48));
  NOR2_X1   g486(.A1(new_n621), .A2(new_n614), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n282), .A2(new_n287), .ZN(new_n674));
  OAI21_X1  g488(.A(G469), .B1(new_n674), .B2(G902), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n285), .A2(new_n278), .A3(new_n280), .A4(new_n198), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n285), .A2(new_n286), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n676), .B1(new_n677), .B2(new_n198), .ZN(new_n678));
  INV_X1    g492(.A(new_n289), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n188), .A3(new_n679), .A4(new_n194), .ZN(new_n680));
  INV_X1    g494(.A(new_n190), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n675), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n544), .A2(new_n673), .A3(new_n591), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT104), .ZN(new_n684));
  INV_X1    g498(.A(new_n591), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT32), .B1(new_n525), .B2(new_n526), .ZN(new_n686));
  INV_X1    g500(.A(new_n526), .ZN(new_n687));
  AOI211_X1 g501(.A(new_n528), .B(new_n687), .C1(new_n523), .C2(new_n524), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n685), .B1(new_n689), .B2(new_n543), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n690), .A2(new_n691), .A3(new_n673), .A4(new_n682), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n684), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT41), .B(G113), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT105), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n693), .B(new_n695), .ZN(G15));
  NOR2_X1   g510(.A1(new_n621), .A2(new_n626), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n544), .A2(new_n697), .A3(new_n591), .A4(new_n682), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  INV_X1    g513(.A(new_n490), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n675), .A2(new_n680), .A3(new_n681), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n368), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n544), .A2(new_n700), .A3(new_n637), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  INV_X1    g518(.A(new_n596), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n509), .B(new_n520), .C1(new_n535), .C2(new_n507), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n705), .A2(G472), .B1(new_n526), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n661), .B1(new_n366), .B2(new_n367), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT106), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n648), .A2(new_n710), .A3(new_n661), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n682), .A2(new_n489), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n707), .A2(new_n712), .A3(new_n591), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NAND2_X1  g529(.A1(new_n706), .A2(new_n526), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n635), .B(new_n716), .C1(new_n596), .C2(new_n597), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n669), .A2(new_n368), .A3(new_n701), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n719), .A3(KEYINPUT107), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n620), .A2(new_n682), .A3(new_n668), .A4(new_n666), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n721), .B1(new_n722), .B2(new_n717), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(KEYINPUT108), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(KEYINPUT108), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n681), .B1(new_n290), .B2(new_n296), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n618), .A2(new_n298), .A3(new_n619), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n669), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n690), .A2(new_n728), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n544), .A2(new_n591), .A3(new_n732), .A4(new_n729), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n727), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n217), .ZN(G33));
  NOR2_X1   g551(.A1(new_n730), .A2(new_n731), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n690), .A2(new_n645), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G134), .ZN(G36));
  XNOR2_X1  g554(.A(new_n295), .B(KEYINPUT45), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(G469), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n193), .A2(new_n188), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(new_n742), .B2(new_n744), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(new_n748), .A3(new_n680), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n681), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  OR3_X1    g565(.A1(new_n750), .A2(new_n751), .A3(new_n650), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n599), .B1(new_n589), .B2(new_n634), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n436), .A2(new_n613), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT43), .Z(new_n755));
  AOI21_X1  g569(.A(KEYINPUT44), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n731), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n755), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n751), .B1(new_n750), .B2(new_n650), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n752), .A2(new_n757), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  NOR3_X1   g575(.A1(new_n544), .A2(new_n591), .A3(new_n731), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n749), .A2(KEYINPUT47), .A3(new_n681), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT47), .B1(new_n749), .B2(new_n681), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n670), .B(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n730), .B1(new_n709), .B2(new_n711), .ZN(new_n768));
  INV_X1    g582(.A(new_n643), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n635), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(new_n659), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n768), .A2(new_n659), .A3(KEYINPUT110), .A4(new_n770), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n724), .A2(new_n646), .A3(new_n671), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n767), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n773), .A2(new_n774), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT107), .B1(new_n718), .B2(new_n719), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n722), .A2(new_n717), .A3(new_n721), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n646), .B(new_n671), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n778), .A2(new_n781), .A3(KEYINPUT52), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n698), .A2(new_n703), .A3(new_n714), .ZN(new_n784));
  INV_X1    g598(.A(new_n614), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(new_n436), .B2(new_n480), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n621), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n599), .A3(new_n600), .A4(new_n591), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(new_n638), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n693), .A2(new_n784), .A3(new_n594), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n297), .A2(new_n435), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n731), .A2(new_n480), .A3(new_n769), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n544), .A2(new_n637), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n718), .A2(new_n732), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n735), .A3(new_n733), .A4(new_n739), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n790), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT53), .B1(new_n783), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n733), .A2(new_n735), .A3(new_n739), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n795), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n594), .A2(new_n789), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n693), .A4(new_n784), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n775), .A2(new_n776), .A3(new_n767), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT52), .B1(new_n778), .B2(new_n781), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n803), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n799), .B1(new_n808), .B2(KEYINPUT111), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n803), .B2(new_n806), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n783), .A2(KEYINPUT53), .A3(new_n798), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n809), .A2(KEYINPUT54), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n486), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n755), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n731), .A2(new_n701), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n690), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT48), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(KEYINPUT113), .A3(new_n821), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n659), .A2(new_n818), .A3(new_n486), .A4(new_n685), .ZN(new_n823));
  INV_X1    g637(.A(new_n613), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n436), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n819), .A2(new_n718), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n707), .A2(new_n591), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n827), .A2(new_n816), .A3(new_n701), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n649), .A2(new_n615), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n828), .A2(KEYINPUT50), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT50), .B1(new_n828), .B2(new_n830), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n825), .B(new_n826), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n827), .A2(new_n816), .ZN(new_n835));
  INV_X1    g649(.A(new_n731), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n675), .A2(new_n680), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n191), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n763), .A2(new_n764), .A3(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n834), .B(KEYINPUT51), .C1(new_n837), .C2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n763), .A2(new_n764), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n839), .B(KEYINPUT112), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n837), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n842), .B1(new_n845), .B2(new_n833), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n196), .A2(G952), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n820), .B(KEYINPUT113), .Z(new_n848));
  AOI21_X1  g662(.A(new_n847), .B1(new_n848), .B2(KEYINPUT48), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n822), .A2(new_n841), .A3(new_n846), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n823), .A2(new_n435), .A3(new_n613), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n810), .A2(new_n811), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n814), .A2(new_n850), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n828), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n368), .ZN(new_n856));
  OAI22_X1  g670(.A1(new_n854), .A2(new_n856), .B1(G952), .B2(G953), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n591), .B(new_n191), .C1(KEYINPUT49), .C2(new_n838), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n754), .B(new_n858), .C1(KEYINPUT49), .C2(new_n838), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n298), .A3(new_n649), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n857), .B1(new_n659), .B2(new_n860), .ZN(G75));
  NOR2_X1   g675(.A1(new_n196), .A2(G952), .ZN(new_n862));
  OAI211_X1 g676(.A(G210), .B(G902), .C1(new_n808), .C2(new_n799), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n326), .A2(new_n344), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(new_n342), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT55), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n188), .B1(new_n810), .B2(new_n811), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT56), .B1(new_n871), .B2(G210), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n872), .B2(KEYINPUT114), .ZN(new_n873));
  AND4_X1   g687(.A1(KEYINPUT114), .A2(new_n863), .A3(new_n864), .A4(new_n870), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n867), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(KEYINPUT115), .B(new_n867), .C1(new_n873), .C2(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(G51));
  NAND2_X1  g693(.A1(new_n810), .A2(new_n811), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT54), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n853), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n744), .B(KEYINPUT57), .Z(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT116), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n882), .A2(new_n887), .A3(new_n884), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n678), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n871), .A2(new_n742), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT117), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n862), .B1(new_n889), .B2(new_n891), .ZN(G54));
  AND3_X1   g706(.A1(new_n871), .A2(KEYINPUT58), .A3(G475), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n893), .A2(new_n894), .A3(new_n432), .ZN(new_n895));
  INV_X1    g709(.A(new_n862), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n893), .B2(new_n432), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n893), .B2(new_n432), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n895), .A2(new_n897), .A3(new_n898), .ZN(G60));
  NAND2_X1  g713(.A1(new_n608), .A2(new_n609), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT59), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n882), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n904), .A2(KEYINPUT119), .A3(new_n896), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT119), .B1(new_n904), .B2(new_n896), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n814), .A2(new_n853), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n901), .B1(new_n907), .B2(new_n903), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(G63));
  XNOR2_X1  g723(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n910));
  XOR2_X1   g724(.A(KEYINPUT121), .B(KEYINPUT60), .Z(new_n911));
  NAND2_X1  g725(.A1(G217), .A2(G902), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n880), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n576), .A3(new_n575), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n896), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n632), .A2(new_n633), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n910), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT122), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n916), .A2(new_n918), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT61), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n923), .B(new_n910), .C1(new_n916), .C2(new_n918), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n920), .A2(new_n922), .A3(new_n924), .ZN(G66));
  NAND2_X1  g739(.A1(new_n790), .A2(new_n196), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT123), .Z(new_n927));
  AOI21_X1  g741(.A(new_n196), .B1(new_n487), .B2(new_n335), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT124), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT125), .Z(new_n931));
  INV_X1    g745(.A(G898), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n868), .B1(new_n932), .B2(G953), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G69));
  NOR2_X1   g748(.A1(new_n498), .A2(new_n499), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n414), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n760), .A2(new_n765), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n776), .A2(new_n663), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n786), .A2(new_n731), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n651), .B(new_n942), .C1(new_n592), .C2(new_n593), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n938), .A2(new_n940), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n937), .B1(new_n944), .B2(new_n196), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n752), .A2(new_n690), .A3(new_n712), .A4(new_n759), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n946), .A2(new_n735), .A3(new_n733), .A4(new_n739), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n760), .A2(new_n765), .A3(new_n776), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n196), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n196), .A2(G900), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT126), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n936), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n196), .B1(G227), .B2(G900), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n953), .B(new_n954), .Z(G72));
  XNOR2_X1  g769(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n597), .A2(new_n188), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(new_n957), .Z(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n944), .B2(new_n790), .ZN(new_n960));
  INV_X1    g774(.A(new_n655), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n862), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n947), .A2(new_n948), .A3(new_n790), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n517), .B(new_n537), .C1(new_n963), .C2(new_n958), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n958), .B1(new_n538), .B2(new_n508), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n809), .A2(new_n813), .A3(new_n965), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n962), .A2(new_n964), .A3(new_n966), .ZN(G57));
endmodule


