//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403, new_n1404, new_n1405, new_n1406;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  OAI22_X1  g0021(.A1(new_n218), .A2(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT66), .B(G238), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n223), .B(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT65), .Z(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n212), .B1(new_n215), .B2(new_n217), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n225), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT10), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G226), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  OAI211_X1 g0059(.A(G1), .B(G13), .C1(new_n259), .C2(new_n254), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G274), .A3(new_n256), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT67), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT3), .B(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G223), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n265), .A2(new_n266), .B1(new_n218), .B2(new_n264), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n264), .A2(G222), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n253), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT67), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n258), .A2(new_n271), .A3(new_n261), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n263), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G200), .ZN(new_n274));
  INV_X1    g0074(.A(G190), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(new_n273), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n213), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT68), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G58), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n207), .A2(G33), .ZN(new_n287));
  OR2_X1    g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n207), .A2(new_n259), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(G150), .A2(new_n290), .B1(new_n203), .B2(G20), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n280), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n202), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n278), .B(new_n213), .C1(G1), .C2(new_n207), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n294), .B1(new_n296), .B2(new_n202), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT69), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT9), .B1(new_n292), .B2(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n252), .B1(new_n277), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n277), .A2(new_n303), .A3(new_n252), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n289), .A2(KEYINPUT71), .ZN(new_n308));
  INV_X1    g0108(.A(new_n281), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n289), .A2(KEYINPUT71), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n311), .B1(new_n207), .B2(new_n218), .C1(new_n287), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n279), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n296), .A2(G77), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n314), .B(new_n315), .C1(G77), .C2(new_n293), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n260), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n261), .B1(new_n318), .B2(new_n219), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n264), .A2(G232), .A3(new_n268), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n320), .B1(new_n220), .B2(new_n264), .C1(new_n265), .C2(new_n226), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n319), .B1(new_n321), .B2(new_n253), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n316), .B1(new_n322), .B2(G190), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n322), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n299), .B1(new_n326), .B2(new_n273), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT70), .A2(G179), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT70), .A2(G179), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n327), .B1(new_n331), .B2(new_n273), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n316), .B1(new_n322), .B2(G169), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n322), .A2(new_n330), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n307), .A2(new_n325), .A3(new_n332), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n264), .A2(G226), .A3(new_n268), .ZN(new_n338));
  AND3_X1   g0138(.A1(KEYINPUT72), .A2(G33), .A3(G97), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT72), .B1(G33), .B2(G97), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n338), .B(new_n341), .C1(new_n265), .C2(new_n234), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n253), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n260), .A2(G274), .A3(new_n256), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT73), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n345), .A2(new_n346), .B1(new_n257), .B2(G238), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n261), .A2(KEYINPUT73), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n344), .A2(new_n349), .A3(KEYINPUT13), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT13), .ZN(new_n351));
  INV_X1    g0151(.A(G238), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n261), .A2(KEYINPUT73), .B1(new_n318), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(KEYINPUT73), .B2(new_n261), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n354), .B2(new_n343), .ZN(new_n355));
  OAI21_X1  g0155(.A(G200), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n293), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n357), .A2(KEYINPUT12), .A3(new_n225), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT12), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n293), .B2(G68), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n358), .B(new_n360), .C1(new_n225), .C2(new_n295), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT74), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n362), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n289), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n287), .A2(new_n218), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n279), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT11), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n367), .A2(new_n368), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n363), .A2(new_n364), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT13), .B1(new_n344), .B2(new_n349), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n354), .A2(new_n351), .A3(new_n343), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(G190), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n356), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(G169), .B1(new_n350), .B2(new_n355), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT14), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n373), .A2(G179), .A3(new_n374), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT14), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(G169), .C1(new_n350), .C2(new_n355), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n377), .B1(new_n383), .B2(new_n371), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n284), .A2(new_n225), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n386), .A2(new_n201), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(G20), .B1(G159), .B2(new_n290), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT75), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT3), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(G33), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n259), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT76), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n390), .ZN(new_n395));
  NAND2_X1  g0195(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(G33), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(KEYINPUT77), .A2(KEYINPUT7), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n207), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G68), .ZN(new_n401));
  AOI21_X1  g0201(.A(G20), .B1(new_n393), .B2(new_n397), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT16), .B(new_n388), .C1(new_n401), .C2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(G20), .ZN(new_n408));
  AOI21_X1  g0208(.A(G33), .B1(new_n395), .B2(new_n396), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n390), .A2(G33), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n408), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n407), .B1(new_n264), .B2(G20), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n225), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n388), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n406), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n405), .A2(new_n279), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n357), .B1(new_n283), .B2(new_n285), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT78), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n419), .B(new_n420), .C1(new_n286), .C2(new_n296), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n286), .A2(new_n296), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT78), .B1(new_n422), .B2(new_n418), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n417), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT79), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  MUX2_X1   g0227(.A(G223), .B(G226), .S(G1698), .Z(new_n428));
  NAND3_X1  g0228(.A1(new_n393), .A2(new_n428), .A3(new_n397), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G87), .ZN(new_n430));
  XOR2_X1   g0230(.A(new_n430), .B(KEYINPUT80), .Z(new_n431));
  AOI21_X1  g0231(.A(new_n260), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n261), .B1(new_n318), .B2(new_n234), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT81), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n261), .B(KEYINPUT81), .C1(new_n318), .C2(new_n234), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n433), .A2(new_n436), .A3(new_n437), .A4(new_n330), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT82), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n326), .B1(new_n432), .B2(new_n434), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n438), .B2(new_n440), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n417), .A2(KEYINPUT79), .A3(new_n424), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n427), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT18), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n417), .A2(KEYINPUT79), .A3(new_n424), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT79), .B1(new_n417), .B2(new_n424), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT18), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(new_n443), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n324), .B1(new_n432), .B2(new_n434), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n433), .A2(new_n275), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n436), .A2(new_n437), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n417), .A2(new_n455), .A3(new_n424), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT17), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n417), .A2(new_n455), .A3(new_n424), .A4(KEYINPUT17), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n446), .A2(new_n451), .A3(new_n461), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n337), .A2(new_n385), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n255), .A2(G1), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT5), .B(G41), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n253), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G270), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n466), .A2(new_n260), .A3(G274), .A4(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT90), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n221), .A2(new_n268), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n393), .A2(new_n397), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT88), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT88), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n393), .A2(new_n397), .A3(new_n476), .A4(new_n473), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n393), .A2(new_n397), .A3(G257), .A4(new_n268), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n410), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G303), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT89), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT89), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n478), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n472), .B1(new_n488), .B2(new_n253), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n478), .A2(new_n483), .A3(new_n486), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n486), .B1(new_n478), .B2(new_n483), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n472), .B(new_n253), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n471), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G283), .ZN(new_n495));
  INV_X1    g0295(.A(G97), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n207), .C1(G33), .C2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(new_n279), .C1(new_n207), .C2(G116), .ZN(new_n498));
  XOR2_X1   g0298(.A(new_n498), .B(KEYINPUT20), .Z(new_n499));
  NOR2_X1   g0299(.A1(new_n293), .A2(G116), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n280), .B(new_n293), .C1(G1), .C2(new_n259), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n502), .B2(G116), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n326), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n494), .A2(KEYINPUT21), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n253), .B1(new_n490), .B2(new_n491), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT90), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n492), .ZN(new_n510));
  INV_X1    g0310(.A(G179), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n505), .A2(new_n511), .A3(new_n470), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n470), .B1(new_n509), .B2(new_n492), .ZN(new_n516));
  INV_X1    g0316(.A(new_n506), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT91), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(KEYINPUT91), .B(new_n515), .C1(new_n516), .C2(new_n517), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n514), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(G190), .B(new_n471), .C1(new_n489), .C2(new_n493), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n505), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n516), .A2(new_n324), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT92), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n494), .A2(G200), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT92), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(new_n505), .A4(new_n523), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  OR3_X1    g0331(.A1(new_n255), .A2(KEYINPUT84), .A3(G1), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n206), .A2(G45), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT84), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n532), .A2(new_n260), .A3(new_n534), .A4(G250), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n260), .A2(G274), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(new_n536), .B2(new_n533), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(G238), .A2(G1698), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n219), .B2(G1698), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n393), .A2(new_n540), .A3(new_n397), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n253), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT85), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n260), .B1(new_n541), .B2(new_n542), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT85), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n546), .A2(new_n537), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n326), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n546), .A2(new_n537), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT85), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n547), .B1(new_n546), .B2(new_n537), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n330), .A3(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n393), .A2(new_n397), .A3(new_n207), .A4(G68), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT19), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n287), .B2(new_n496), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT19), .B1(new_n339), .B2(new_n340), .ZN(new_n558));
  INV_X1    g0358(.A(G87), .ZN(new_n559));
  NOR2_X1   g0359(.A1(G97), .A2(G107), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n558), .A2(new_n207), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n279), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n312), .A2(new_n357), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n501), .A2(new_n312), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT86), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT86), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n562), .A2(new_n567), .A3(new_n563), .A4(new_n564), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n549), .A2(new_n553), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n408), .ZN(new_n570));
  AND2_X1   g0370(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n571));
  NOR2_X1   g0371(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n259), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n570), .B1(new_n573), .B2(new_n410), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT7), .B1(new_n481), .B2(new_n207), .ZN(new_n575));
  OAI21_X1  g0375(.A(G107), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT6), .ZN(new_n577));
  AND2_X1   g0377(.A1(G97), .A2(G107), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(new_n560), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n220), .A2(KEYINPUT6), .A3(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n280), .B1(new_n576), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n357), .A2(new_n496), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n501), .B2(new_n496), .ZN(new_n585));
  OAI21_X1  g0385(.A(KEYINPUT83), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n220), .B1(new_n412), .B2(new_n413), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n581), .A2(G20), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n290), .A2(G77), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n279), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT83), .ZN(new_n592));
  INV_X1    g0392(.A(new_n585), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT4), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n595), .A2(new_n219), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n264), .A2(new_n268), .A3(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n480), .A2(new_n410), .A3(G250), .A4(G1698), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n597), .A2(new_n495), .A3(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n393), .A2(new_n397), .A3(G244), .A4(new_n268), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n595), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n253), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n466), .A2(new_n465), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n260), .ZN(new_n605));
  INV_X1    g0405(.A(G257), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n469), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(G200), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n260), .B1(new_n599), .B2(new_n601), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n610), .A2(G190), .A3(new_n607), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n586), .B(new_n594), .C1(new_n609), .C2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n545), .B2(new_n548), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n551), .A2(G190), .A3(new_n552), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n502), .A2(G87), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n562), .A2(new_n563), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(G169), .B1(new_n610), .B2(new_n607), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n597), .A2(new_n495), .A3(new_n598), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n595), .B2(new_n600), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n331), .B(new_n608), .C1(new_n620), .C2(new_n260), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n576), .A2(new_n582), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n585), .B1(new_n623), .B2(new_n279), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n569), .A2(new_n612), .A3(new_n617), .A4(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT87), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n624), .B1(new_n618), .B2(new_n621), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n594), .A2(new_n586), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n603), .A2(new_n275), .A3(new_n608), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n610), .A2(new_n607), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n632), .B1(G200), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n630), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n635), .A2(KEYINPUT87), .A3(new_n617), .A4(new_n569), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n469), .B1(new_n605), .B2(new_n221), .ZN(new_n637));
  NOR2_X1   g0437(.A1(G250), .A2(G1698), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n606), .B2(G1698), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n393), .A2(new_n639), .A3(new_n397), .ZN(new_n640));
  XNOR2_X1  g0440(.A(KEYINPUT94), .B(G294), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G33), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n260), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n275), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(G200), .B2(new_n644), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n357), .A2(KEYINPUT25), .A3(new_n220), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(KEYINPUT25), .B1(new_n357), .B2(new_n220), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n501), .A2(new_n220), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT22), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(new_n559), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n393), .A2(new_n397), .A3(new_n207), .A4(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n559), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n264), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n652), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n542), .A2(G20), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT23), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n207), .B2(G107), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n220), .A2(KEYINPUT23), .A3(G20), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n654), .A2(new_n657), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT24), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT22), .B1(new_n264), .B2(new_n655), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n660), .A2(new_n661), .ZN(new_n666));
  INV_X1    g0466(.A(new_n658), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT24), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(new_n654), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT93), .B1(new_n672), .B2(new_n279), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT93), .ZN(new_n674));
  AOI211_X1 g0474(.A(new_n674), .B(new_n280), .C1(new_n664), .C2(new_n671), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n646), .B(new_n651), .C1(new_n673), .C2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n663), .A2(KEYINPUT24), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n670), .B1(new_n669), .B2(new_n654), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n279), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n674), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n672), .A2(KEYINPUT93), .A3(new_n279), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n650), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NOR4_X1   g0482(.A1(new_n637), .A2(new_n643), .A3(KEYINPUT95), .A4(new_n511), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT95), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n644), .B2(new_n326), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n644), .A2(G179), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n676), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n629), .A2(new_n636), .A3(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n464), .A2(new_n531), .A3(new_n690), .ZN(G372));
  NAND2_X1  g0491(.A1(new_n438), .A2(new_n440), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT82), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n421), .A2(new_n423), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n402), .A2(new_n403), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n225), .B1(new_n402), .B2(new_n399), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n415), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n280), .B1(new_n699), .B2(KEYINPUT16), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n696), .B1(new_n700), .B2(new_n416), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT96), .B1(new_n695), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT96), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n443), .A2(new_n703), .A3(new_n425), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(new_n704), .A3(KEYINPUT18), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n695), .A2(new_n701), .A3(KEYINPUT96), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n703), .B1(new_n443), .B2(new_n425), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n450), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n383), .A2(new_n371), .B1(new_n376), .B2(new_n335), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n705), .B(new_n708), .C1(new_n709), .C2(new_n460), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT97), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT97), .ZN(new_n712));
  INV_X1    g0512(.A(new_n306), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n304), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(new_n711), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n332), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT98), .Z(new_n717));
  OAI211_X1 g0517(.A(new_n614), .B(new_n616), .C1(new_n324), .C2(new_n550), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n553), .B(new_n565), .C1(G169), .C2(new_n550), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT26), .ZN(new_n722));
  INV_X1    g0522(.A(new_n631), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n721), .A2(new_n722), .A3(new_n622), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n569), .A2(new_n630), .A3(new_n617), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT26), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n724), .A2(new_n719), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n516), .A2(new_n517), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n728), .A2(KEYINPUT21), .B1(new_n510), .B2(new_n512), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n682), .A2(new_n687), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n494), .A2(new_n506), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT91), .B1(new_n731), .B2(new_n515), .ZN(new_n732));
  INV_X1    g0532(.A(new_n521), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n729), .B(new_n730), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n721), .A2(new_n635), .A3(new_n676), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n727), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n717), .B1(new_n464), .B2(new_n737), .ZN(G369));
  INV_X1    g0538(.A(G330), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT27), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT27), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(G213), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G343), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n505), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n522), .A2(new_n530), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n747), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n739), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n682), .A2(new_n746), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n730), .A2(new_n746), .B1(new_n688), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n730), .A2(new_n745), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n520), .A2(new_n521), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n745), .B1(new_n757), .B2(new_n729), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n756), .B1(new_n758), .B2(new_n689), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n755), .A2(new_n759), .ZN(G399));
  INV_X1    g0560(.A(new_n210), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G41), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n206), .ZN(new_n763));
  INV_X1    g0563(.A(G116), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n560), .A2(new_n559), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n217), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n763), .A2(new_n766), .B1(new_n767), .B2(new_n762), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT28), .Z(new_n769));
  INV_X1    g0569(.A(new_n468), .ZN(new_n770));
  NOR4_X1   g0570(.A1(new_n770), .A2(new_n637), .A3(new_n643), .A4(new_n511), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n771), .A2(new_n633), .A3(new_n552), .A4(new_n551), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n509), .B2(new_n492), .ZN(new_n773));
  NOR4_X1   g0573(.A1(new_n633), .A2(new_n331), .A3(new_n550), .A4(new_n644), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI22_X1  g0575(.A1(KEYINPUT30), .A2(new_n773), .B1(new_n516), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n772), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n489), .B2(new_n493), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT30), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(KEYINPUT31), .B(new_n745), .C1(new_n776), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n778), .A2(new_n779), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n494), .A2(new_n774), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n773), .A2(KEYINPUT30), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(KEYINPUT31), .B1(new_n786), .B2(new_n745), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  AND4_X1   g0588(.A1(new_n629), .A2(new_n636), .A3(new_n689), .A4(new_n746), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n530), .A2(new_n757), .A3(new_n729), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n739), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n734), .A2(new_n736), .ZN(new_n793));
  INV_X1    g0593(.A(new_n727), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(KEYINPUT29), .B1(new_n795), .B2(new_n746), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n723), .A2(new_n622), .ZN(new_n797));
  OAI21_X1  g0597(.A(KEYINPUT26), .B1(new_n797), .B2(new_n720), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n798), .B(new_n719), .C1(KEYINPUT26), .C2(new_n725), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(new_n734), .B2(new_n736), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT29), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n800), .A2(new_n801), .A3(new_n745), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n792), .B1(new_n796), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(KEYINPUT99), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n801), .B1(new_n737), .B2(new_n745), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n735), .B1(new_n522), .B2(new_n730), .ZN(new_n806));
  OAI211_X1 g0606(.A(KEYINPUT29), .B(new_n746), .C1(new_n806), .C2(new_n799), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT99), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n808), .A2(new_n809), .A3(new_n792), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n804), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n769), .B1(new_n811), .B2(G1), .ZN(G364));
  NAND2_X1  g0612(.A1(new_n207), .A2(G13), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT100), .Z(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G45), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n763), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n752), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n749), .A2(new_n751), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(G330), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n213), .B1(G20), .B2(new_n326), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT106), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n207), .A2(new_n324), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n331), .A2(G190), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT103), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n826), .A2(KEYINPUT103), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G326), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n207), .A2(G190), .ZN(new_n833));
  NOR2_X1   g0633(.A1(G179), .A2(G200), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n264), .B1(new_n836), .B2(G329), .ZN(new_n837));
  INV_X1    g0637(.A(new_n641), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n275), .A2(G179), .A3(G200), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n207), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n837), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n331), .A2(new_n324), .A3(new_n833), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n841), .B1(G311), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n207), .A2(new_n275), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(new_n511), .A3(G200), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT104), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n331), .A2(new_n275), .A3(new_n824), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(KEYINPUT33), .B(G317), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n851), .A2(G303), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n833), .A2(new_n511), .A3(G200), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT105), .Z(new_n857));
  NAND3_X1  g0657(.A1(new_n331), .A2(new_n324), .A3(new_n845), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n857), .A2(G283), .B1(G322), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n832), .A2(new_n844), .A3(new_n855), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n840), .A2(new_n496), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n481), .B(new_n862), .C1(new_n843), .C2(G77), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n857), .A2(G107), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n863), .B(new_n864), .C1(new_n284), .C2(new_n858), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n836), .A2(G159), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT32), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n852), .A2(new_n225), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n850), .A2(new_n559), .ZN(new_n869));
  NOR4_X1   g0669(.A1(new_n865), .A2(new_n867), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n831), .A2(G50), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n823), .A2(new_n861), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n861), .A2(new_n823), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n822), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(G13), .A2(G33), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(G20), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(new_n821), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n210), .A2(new_n264), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT101), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n880), .A2(G355), .B1(new_n764), .B2(new_n761), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n881), .A2(KEYINPUT102), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(KEYINPUT102), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n398), .A2(new_n210), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n255), .B2(new_n767), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n255), .B2(new_n250), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n882), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n816), .B(new_n874), .C1(new_n878), .C2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n877), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n888), .B1(new_n819), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n820), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(G396));
  NAND2_X1  g0692(.A1(new_n316), .A2(new_n745), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n325), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n336), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n335), .A2(new_n746), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n737), .B2(new_n745), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n746), .B(new_n899), .C1(new_n806), .C2(new_n727), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n817), .B1(new_n903), .B2(new_n792), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n792), .B2(new_n903), .ZN(new_n905));
  AOI22_X1  g0705(.A1(G150), .A2(new_n853), .B1(new_n843), .B2(G159), .ZN(new_n906));
  XNOR2_X1  g0706(.A(KEYINPUT109), .B(G143), .ZN(new_n907));
  INV_X1    g0707(.A(G137), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n906), .B1(new_n858), .B2(new_n907), .C1(new_n830), .C2(new_n908), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT34), .Z(new_n910));
  AOI21_X1  g0710(.A(new_n398), .B1(G132), .B2(new_n836), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n284), .B2(new_n840), .ZN(new_n912));
  INV_X1    g0712(.A(new_n857), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n225), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n850), .A2(new_n202), .ZN(new_n915));
  NOR4_X1   g0715(.A1(new_n910), .A2(new_n912), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n857), .A2(G87), .ZN(new_n917));
  INV_X1    g0717(.A(G311), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n917), .B1(new_n918), .B2(new_n835), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT108), .Z(new_n920));
  OAI21_X1  g0720(.A(new_n481), .B1(new_n850), .B2(new_n220), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT107), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n831), .A2(G303), .ZN(new_n923));
  INV_X1    g0723(.A(G283), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n764), .A2(new_n842), .B1(new_n852), .B2(new_n924), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n862), .B(new_n925), .C1(G294), .C2(new_n859), .ZN(new_n926));
  AND4_X1   g0726(.A1(new_n920), .A2(new_n922), .A3(new_n923), .A4(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n821), .B1(new_n916), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n821), .A2(new_n875), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n816), .B1(new_n218), .B2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n928), .B(new_n930), .C1(new_n899), .C2(new_n876), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n905), .A2(new_n931), .ZN(G384));
  NOR2_X1   g0732(.A1(new_n699), .A2(KEYINPUT16), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n405), .A2(new_n279), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n424), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n743), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n462), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT37), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n456), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n449), .B2(new_n443), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n447), .A2(new_n448), .A3(new_n743), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n935), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n937), .B(new_n456), .C1(new_n946), .C2(new_n695), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT37), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n939), .A2(new_n949), .A3(KEYINPUT38), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n708), .A2(new_n461), .A3(new_n705), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n702), .A2(new_n704), .A3(new_n456), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT37), .B1(new_n952), .B2(new_n943), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n951), .A2(new_n943), .B1(new_n953), .B2(new_n945), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n950), .B1(new_n954), .B2(KEYINPUT38), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT39), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n383), .A2(new_n371), .A3(new_n746), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT38), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n460), .B1(KEYINPUT18), .B2(new_n445), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n937), .B1(new_n961), .B2(new_n451), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n942), .A2(new_n944), .B1(new_n947), .B2(KEYINPUT37), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(new_n950), .A3(KEYINPUT39), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n957), .A2(new_n959), .A3(new_n965), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n708), .A2(new_n705), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(new_n936), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n964), .A2(new_n950), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n371), .B(new_n745), .C1(new_n383), .C2(new_n377), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n371), .A2(new_n745), .ZN(new_n972));
  AOI21_X1  g0772(.A(KEYINPUT110), .B1(new_n384), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n382), .A2(new_n380), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n373), .A2(new_n374), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n381), .B1(new_n975), .B2(G169), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n371), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  AND4_X1   g0777(.A1(KEYINPUT110), .A2(new_n977), .A3(new_n376), .A4(new_n972), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n971), .B1(new_n973), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n970), .B(new_n980), .C1(new_n902), .C2(new_n897), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n969), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n805), .A2(new_n807), .A3(new_n463), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n717), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n982), .B(new_n984), .Z(new_n985));
  NAND2_X1  g0785(.A1(new_n979), .A2(new_n899), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n788), .A2(new_n790), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(new_n955), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n986), .B1(new_n790), .B2(new_n788), .ZN(new_n990));
  AOI21_X1  g0790(.A(KEYINPUT40), .B1(new_n964), .B2(new_n950), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n989), .A2(KEYINPUT40), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n464), .B1(new_n788), .B2(new_n790), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n739), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n994), .B2(new_n993), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n985), .A2(new_n996), .B1(new_n206), .B2(new_n814), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT111), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n998), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n985), .A2(new_n996), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n1004));
  NOR4_X1   g0804(.A1(new_n1003), .A2(new_n215), .A3(new_n1004), .A4(new_n764), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT36), .ZN(new_n1006));
  OR3_X1    g0806(.A1(new_n217), .A2(new_n218), .A3(new_n386), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n206), .B(G13), .C1(new_n1007), .C2(new_n246), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1002), .A2(new_n1009), .ZN(G367));
  OAI221_X1 g0810(.A(new_n878), .B1(new_n210), .B2(new_n312), .C1(new_n241), .C2(new_n884), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n817), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT113), .Z(new_n1013));
  AOI22_X1  g0813(.A1(G303), .A2(new_n859), .B1(new_n853), .B2(new_n641), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n924), .B2(new_n842), .C1(new_n830), .C2(new_n918), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n851), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT46), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n850), .B2(new_n764), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n840), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(G107), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n398), .ZN(new_n1021));
  INV_X1    g0821(.A(G317), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n856), .A2(new_n496), .B1(new_n835), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1016), .A2(new_n1018), .A3(new_n1020), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n830), .A2(new_n907), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n851), .A2(G58), .B1(G159), .B2(new_n853), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1019), .A2(G68), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n264), .B1(new_n856), .B2(new_n218), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G137), .B2(new_n836), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G150), .A2(new_n859), .B1(new_n843), .B2(G50), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1015), .A2(new_n1025), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT47), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n822), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1013), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n616), .A2(new_n746), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n721), .A2(new_n1038), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n719), .A2(new_n1038), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n877), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n635), .B1(new_n631), .B2(new_n746), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n723), .A2(new_n622), .A3(new_n745), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n758), .A2(new_n689), .A3(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1046), .A2(KEYINPUT42), .B1(new_n630), .B2(new_n746), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n750), .A2(new_n689), .A3(new_n746), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n756), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1045), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(KEYINPUT42), .B2(new_n1049), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n1047), .A2(new_n1053), .B1(KEYINPUT43), .B2(new_n1054), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(KEYINPUT43), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n755), .A2(new_n1051), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1059));
  AND3_X1   g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1058), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n815), .A2(G1), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT44), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n759), .B2(new_n1045), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1050), .A2(KEYINPUT44), .A3(new_n1051), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1048), .A2(new_n1049), .A3(new_n1045), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT45), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n759), .A2(KEYINPUT45), .A3(new_n1045), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT112), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n752), .A2(new_n1074), .A3(new_n754), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n1068), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1075), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1048), .B1(new_n754), .B2(new_n758), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n752), .B(new_n1079), .Z(new_n1080));
  OAI21_X1  g0880(.A(new_n811), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n762), .B(KEYINPUT41), .Z(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1064), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1042), .B1(new_n1063), .B2(new_n1084), .ZN(G387));
  XNOR2_X1  g0885(.A(new_n752), .B(new_n1079), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n809), .B1(new_n808), .B2(new_n792), .ZN(new_n1087));
  AOI211_X1 g0887(.A(KEYINPUT99), .B(new_n791), .C1(new_n805), .C2(new_n807), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n804), .A2(new_n810), .A3(new_n1080), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n1090), .A3(new_n762), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n754), .A2(new_n889), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n880), .A2(new_n765), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n237), .A2(new_n255), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n884), .ZN(new_n1095));
  OR3_X1    g0895(.A1(new_n281), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1096));
  OAI21_X1  g0896(.A(KEYINPUT50), .B1(new_n281), .B2(G50), .ZN(new_n1097));
  AOI21_X1  g0897(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1096), .A2(new_n766), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1095), .A2(new_n1099), .B1(new_n220), .B2(new_n761), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n878), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n817), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n851), .A2(G77), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n202), .B2(new_n858), .C1(new_n225), .C2(new_n842), .ZN(new_n1104));
  INV_X1    g0904(.A(G159), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n830), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(G150), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1021), .B1(new_n1107), .B2(new_n835), .C1(new_n312), .C2(new_n840), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n913), .A2(new_n496), .B1(new_n286), .B2(new_n852), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1104), .A2(new_n1106), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT114), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n856), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1112), .A2(G116), .B1(new_n836), .B2(G326), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n850), .A2(new_n838), .B1(new_n924), .B2(new_n840), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n918), .A2(new_n852), .B1(new_n858), .B2(new_n1022), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(G303), .B2(new_n843), .ZN(new_n1116));
  INV_X1    g0916(.A(G322), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n830), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT48), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1114), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n1119), .B2(new_n1118), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT49), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n398), .B(new_n1113), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1111), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1102), .B1(new_n1125), .B2(new_n821), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1086), .A2(new_n1064), .B1(new_n1092), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1091), .A2(new_n1127), .ZN(G393));
  AND3_X1   g0928(.A1(new_n1068), .A2(new_n1073), .A3(new_n755), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n755), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1051), .A2(new_n877), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n878), .B1(new_n496), .B2(new_n210), .C1(new_n245), .C2(new_n884), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n817), .A2(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n830), .A2(new_n1022), .B1(new_n918), .B2(new_n858), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT52), .Z(new_n1136));
  AOI21_X1  g0936(.A(new_n264), .B1(new_n836), .B2(G322), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n864), .B(new_n1137), .C1(new_n764), .C2(new_n840), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G303), .A2(new_n853), .B1(new_n843), .B2(G294), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n924), .B2(new_n850), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n1136), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n830), .A2(new_n1107), .B1(new_n1105), .B2(new_n858), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT51), .Z(new_n1143));
  OAI221_X1 g0943(.A(new_n1021), .B1(new_n218), .B2(new_n840), .C1(new_n835), .C2(new_n907), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n851), .A2(G68), .B1(new_n309), .B2(new_n843), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1145), .B(new_n917), .C1(new_n202), .C2(new_n852), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1134), .B1(new_n1148), .B2(new_n821), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1131), .A2(new_n1064), .B1(new_n1132), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n762), .B1(new_n1078), .B2(new_n1089), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1130), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1068), .A2(new_n1073), .A3(new_n755), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n811), .A2(new_n1086), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1150), .B1(new_n1151), .B2(new_n1154), .ZN(G390));
  NAND4_X1  g0955(.A1(new_n988), .A2(G330), .A3(new_n899), .A4(new_n979), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n964), .A2(new_n950), .A3(KEYINPUT39), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n956), .B2(new_n955), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n737), .A2(new_n745), .A3(new_n900), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n979), .B1(new_n1160), .B2(new_n898), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1159), .B1(new_n1161), .B2(new_n958), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n955), .A2(new_n958), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n746), .B1(new_n806), .B2(new_n799), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n897), .B1(new_n1164), .B2(new_n896), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1163), .B1(new_n1165), .B2(new_n979), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1157), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1156), .A2(KEYINPUT115), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT115), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n791), .A2(new_n1169), .A3(new_n899), .A4(new_n979), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n957), .A2(new_n965), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n980), .B1(new_n902), .B2(new_n897), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n959), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n800), .A2(new_n745), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n898), .B1(new_n1176), .B2(new_n895), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n958), .B(new_n955), .C1(new_n1177), .C2(new_n980), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1172), .A2(new_n1175), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1167), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n979), .B1(new_n791), .B2(new_n899), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1182), .A2(new_n1168), .A3(new_n1177), .A4(new_n1170), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n902), .A2(new_n897), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1156), .A2(KEYINPUT116), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1184), .B1(new_n1185), .B2(new_n1181), .ZN(new_n1186));
  AOI211_X1 g0986(.A(KEYINPUT116), .B(new_n979), .C1(new_n791), .C2(new_n899), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1183), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n717), .B(new_n983), .C1(new_n464), .C2(new_n792), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1180), .A2(new_n1191), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1167), .A2(new_n1188), .A3(new_n1179), .A4(new_n1190), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n762), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1173), .A2(new_n875), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n286), .A2(new_n929), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n831), .A2(G128), .ZN(new_n1197));
  INV_X1    g0997(.A(G125), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n264), .B1(new_n835), .B2(new_n1198), .C1(new_n202), .C2(new_n856), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G159), .B2(new_n1019), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT54), .B(G143), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n908), .A2(new_n852), .B1(new_n842), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G132), .B2(new_n859), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n850), .A2(new_n1107), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT53), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1197), .A2(new_n1200), .A3(new_n1203), .A4(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n842), .A2(new_n496), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1207), .B(new_n914), .C1(G107), .C2(new_n853), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n264), .B(new_n869), .C1(G294), .C2(new_n836), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1208), .B(new_n1209), .C1(new_n924), .C2(new_n830), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n858), .A2(new_n764), .B1(new_n840), .B2(new_n218), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT117), .Z(new_n1212));
  OAI21_X1  g1012(.A(new_n1206), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n816), .B(new_n1196), .C1(new_n1213), .C2(new_n821), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1195), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1064), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1215), .B1(new_n1180), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1194), .A2(new_n1218), .ZN(G378));
  XOR2_X1   g1019(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n711), .A2(new_n714), .A3(new_n332), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n299), .A2(new_n743), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT119), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1223), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n711), .A2(new_n714), .A3(new_n332), .A4(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1225), .B1(new_n1224), .B2(new_n1227), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1221), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT119), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1224), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1220), .A3(new_n1233), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1230), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n992), .B2(new_n739), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1230), .A2(new_n1234), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT40), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(new_n990), .B2(new_n955), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n987), .A2(new_n991), .A3(new_n988), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1237), .B(G330), .C1(new_n1239), .C2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1236), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n982), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1236), .A2(new_n982), .A3(new_n1241), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1235), .A2(new_n875), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n929), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n817), .B1(G50), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n398), .A2(new_n254), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1250), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n853), .B2(G97), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1252), .B1(new_n220), .B2(new_n858), .C1(new_n312), .C2(new_n842), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1112), .A2(G58), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n836), .A2(G283), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1103), .A2(new_n1028), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1253), .B(new_n1256), .C1(G116), .C2(new_n831), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1251), .B1(new_n1257), .B2(KEYINPUT58), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(KEYINPUT58), .B2(new_n1257), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n853), .A2(G132), .B1(G150), .B2(new_n1019), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n908), .B2(new_n842), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1201), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n851), .A2(new_n1262), .B1(G128), .B2(new_n859), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT118), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n1261), .B(new_n1264), .C1(G125), .C2(new_n831), .ZN(new_n1265));
  XOR2_X1   g1065(.A(new_n1265), .B(KEYINPUT59), .Z(new_n1266));
  AOI211_X1 g1066(.A(G33), .B(G41), .C1(new_n1112), .C2(G159), .ZN(new_n1267));
  INV_X1    g1067(.A(G124), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1267), .B1(new_n1268), .B2(new_n835), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1259), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1249), .B1(new_n1270), .B2(new_n821), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1246), .A2(new_n1064), .B1(new_n1247), .B2(new_n1271), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1162), .A2(new_n1166), .A3(new_n1171), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1156), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1189), .B1(new_n1275), .B2(new_n1188), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1236), .A2(new_n982), .A3(new_n1241), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n982), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT57), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n762), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1188), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1190), .B1(new_n1180), .B2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT57), .B1(new_n1282), .B2(new_n1246), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1272), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT120), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(G375));
  OAI211_X1 g1089(.A(new_n1189), .B(new_n1183), .C1(new_n1187), .C2(new_n1186), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1191), .A2(new_n1083), .A3(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n979), .A2(new_n876), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(KEYINPUT121), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n264), .B1(new_n836), .B2(G303), .ZN(new_n1294));
  OAI221_X1 g1094(.A(new_n1294), .B1(new_n312), .B2(new_n840), .C1(new_n852), .C2(new_n764), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n857), .A2(G77), .B1(G107), .B2(new_n843), .ZN(new_n1296));
  OAI221_X1 g1096(.A(new_n1296), .B1(new_n496), .B2(new_n850), .C1(new_n924), .C2(new_n858), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1295), .B(new_n1297), .C1(G294), .C2(new_n831), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1112), .A2(G58), .B1(new_n836), .B2(G128), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1299), .B(new_n1021), .C1(new_n202), .C2(new_n840), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(G137), .A2(new_n859), .B1(new_n853), .B2(new_n1262), .ZN(new_n1301));
  OAI221_X1 g1101(.A(new_n1301), .B1(new_n1107), .B2(new_n842), .C1(new_n1105), .C2(new_n850), .ZN(new_n1302));
  AOI211_X1 g1102(.A(new_n1300), .B(new_n1302), .C1(G132), .C2(new_n831), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n821), .B1(new_n1298), .B2(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1304), .B(new_n817), .C1(G68), .C2(new_n1248), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1293), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1188), .B2(new_n1064), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1291), .A2(new_n1307), .ZN(G381));
  AND3_X1   g1108(.A1(new_n1091), .A2(new_n891), .A3(new_n1127), .ZN(new_n1309));
  INV_X1    g1109(.A(G384), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(KEYINPUT122), .ZN(new_n1312));
  NOR4_X1   g1112(.A1(G387), .A2(G378), .A3(G390), .A4(G381), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1312), .B(new_n1313), .C1(new_n1287), .C2(new_n1288), .ZN(G407));
  INV_X1    g1114(.A(new_n762), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1180), .B2(new_n1191), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1217), .B1(new_n1316), .B2(new_n1193), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1318));
  OAI211_X1 g1118(.A(G407), .B(G213), .C1(new_n1318), .C2(G343), .ZN(G409));
  OAI211_X1 g1119(.A(G378), .B(new_n1272), .C1(new_n1280), .C2(new_n1283), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1282), .A2(new_n1083), .A3(new_n1246), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1246), .A2(new_n1064), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1247), .A2(new_n1271), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1317), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1320), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n744), .A2(G213), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n744), .A2(G213), .A3(G2897), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  XOR2_X1   g1130(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n1331));
  NAND2_X1  g1131(.A1(new_n1290), .A2(new_n1331), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1156), .A2(KEYINPUT116), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1182), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1187), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(new_n1184), .A3(new_n1335), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1336), .A2(KEYINPUT60), .A3(new_n1189), .A4(new_n1183), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1332), .A2(new_n762), .A3(new_n1337), .A4(new_n1191), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1338), .A2(G384), .A3(new_n1307), .ZN(new_n1339));
  AOI21_X1  g1139(.A(G384), .B1(new_n1338), .B2(new_n1307), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1330), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1338), .A2(new_n1307), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1310), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1338), .A2(G384), .A3(new_n1307), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1344), .A3(new_n1329), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1341), .A2(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(KEYINPUT61), .B1(new_n1328), .B2(new_n1346), .ZN(new_n1347));
  AOI22_X1  g1147(.A1(new_n1320), .A2(new_n1325), .B1(G213), .B2(new_n744), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1348), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1326), .A2(new_n1327), .A3(new_n1349), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT62), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1353), .A2(KEYINPUT126), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1352), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1347), .A2(new_n1351), .A3(new_n1355), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1152), .A2(new_n1064), .A3(new_n1153), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1149), .A2(new_n1132), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1080), .B1(new_n804), .B2(new_n810), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1075), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1068), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1315), .B1(new_n1360), .B2(new_n1365), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1089), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1359), .B1(new_n1366), .B2(new_n1367), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n891), .B1(new_n1091), .B2(new_n1127), .ZN(new_n1369));
  NOR3_X1   g1169(.A1(new_n1368), .A2(new_n1309), .A3(new_n1369), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1091), .A2(new_n891), .A3(new_n1127), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(G393), .A2(G396), .ZN(new_n1372));
  AOI21_X1  g1172(.A(G390), .B1(new_n1371), .B2(new_n1372), .ZN(new_n1373));
  OAI21_X1  g1173(.A(G387), .B1(new_n1370), .B2(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1042), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1376), .A2(new_n1216), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1375), .B1(new_n1377), .B2(new_n1062), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1372), .A2(G390), .A3(new_n1371), .ZN(new_n1379));
  OAI21_X1  g1179(.A(new_n1368), .B1(new_n1309), .B2(new_n1369), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1378), .A2(new_n1379), .A3(new_n1380), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1374), .A2(new_n1381), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1356), .A2(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(KEYINPUT61), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1374), .A2(new_n1384), .A3(new_n1381), .ZN(new_n1385));
  INV_X1    g1185(.A(KEYINPUT124), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1385), .A2(new_n1386), .ZN(new_n1387));
  NAND4_X1  g1187(.A1(new_n1374), .A2(new_n1381), .A3(KEYINPUT124), .A4(new_n1384), .ZN(new_n1388));
  AOI22_X1  g1188(.A1(new_n1387), .A2(new_n1388), .B1(new_n1328), .B2(new_n1346), .ZN(new_n1389));
  INV_X1    g1189(.A(KEYINPUT125), .ZN(new_n1390));
  NAND4_X1  g1190(.A1(new_n1348), .A2(new_n1390), .A3(KEYINPUT63), .A4(new_n1349), .ZN(new_n1391));
  INV_X1    g1191(.A(KEYINPUT63), .ZN(new_n1392));
  OAI21_X1  g1192(.A(KEYINPUT125), .B1(new_n1352), .B2(new_n1392), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1352), .A2(new_n1392), .ZN(new_n1394));
  NAND4_X1  g1194(.A1(new_n1389), .A2(new_n1391), .A3(new_n1393), .A4(new_n1394), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1383), .A2(new_n1395), .ZN(G405));
  INV_X1    g1196(.A(new_n1349), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1382), .A2(new_n1397), .ZN(new_n1398));
  NAND3_X1  g1198(.A1(new_n1374), .A2(new_n1381), .A3(new_n1349), .ZN(new_n1399));
  INV_X1    g1199(.A(new_n1288), .ZN(new_n1400));
  AOI21_X1  g1200(.A(G378), .B1(new_n1400), .B2(new_n1286), .ZN(new_n1401));
  INV_X1    g1201(.A(new_n1284), .ZN(new_n1402));
  NOR2_X1   g1202(.A1(new_n1402), .A2(new_n1317), .ZN(new_n1403));
  OAI211_X1 g1203(.A(new_n1398), .B(new_n1399), .C1(new_n1401), .C2(new_n1403), .ZN(new_n1404));
  NAND2_X1  g1204(.A1(new_n1398), .A2(new_n1399), .ZN(new_n1405));
  OAI211_X1 g1205(.A(new_n1405), .B(new_n1318), .C1(new_n1317), .C2(new_n1402), .ZN(new_n1406));
  AND2_X1   g1206(.A1(new_n1404), .A2(new_n1406), .ZN(G402));
endmodule


