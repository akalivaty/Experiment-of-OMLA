

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U320 ( .A(n496), .B(KEYINPUT111), .ZN(n497) );
  XNOR2_X1 U321 ( .A(n498), .B(n497), .ZN(n499) );
  NOR2_X1 U322 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U323 ( .A(n305), .B(n384), .ZN(n306) );
  NOR2_X1 U324 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U325 ( .A(n307), .B(n306), .ZN(n309) );
  NOR2_X1 U326 ( .A1(n552), .A2(n551), .ZN(n564) );
  XOR2_X1 U327 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n450) );
  XOR2_X1 U328 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n289) );
  XNOR2_X1 U329 ( .A(G176GAT), .B(G204GAT), .ZN(n288) );
  XNOR2_X1 U330 ( .A(n289), .B(n288), .ZN(n291) );
  INV_X1 U331 ( .A(n291), .ZN(n290) );
  XOR2_X1 U332 ( .A(G92GAT), .B(G64GAT), .Z(n424) );
  NAND2_X1 U333 ( .A1(n290), .A2(n424), .ZN(n294) );
  INV_X1 U334 ( .A(n424), .ZN(n292) );
  NAND2_X1 U335 ( .A1(n292), .A2(n291), .ZN(n293) );
  NAND2_X1 U336 ( .A1(n294), .A2(n293), .ZN(n296) );
  NAND2_X1 U337 ( .A1(G230GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U339 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n298) );
  XNOR2_X1 U340 ( .A(KEYINPUT80), .B(KEYINPUT76), .ZN(n297) );
  XOR2_X1 U341 ( .A(n298), .B(n297), .Z(n299) );
  XNOR2_X1 U342 ( .A(n300), .B(n299), .ZN(n307) );
  XNOR2_X1 U343 ( .A(G99GAT), .B(G71GAT), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n301), .B(G120GAT), .ZN(n377) );
  XNOR2_X1 U345 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n302), .B(KEYINPUT74), .ZN(n359) );
  XNOR2_X1 U347 ( .A(n377), .B(n359), .ZN(n305) );
  XOR2_X1 U348 ( .A(G78GAT), .B(G148GAT), .Z(n304) );
  XNOR2_X1 U349 ( .A(G106GAT), .B(KEYINPUT77), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n384) );
  XNOR2_X1 U351 ( .A(G85GAT), .B(KEYINPUT78), .ZN(n308) );
  XNOR2_X1 U352 ( .A(n308), .B(KEYINPUT79), .ZN(n333) );
  XNOR2_X1 U353 ( .A(n309), .B(n333), .ZN(n474) );
  XNOR2_X1 U354 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n310), .B(G8GAT), .ZN(n360) );
  XOR2_X1 U356 ( .A(n360), .B(G197GAT), .Z(n312) );
  XOR2_X1 U357 ( .A(G141GAT), .B(G22GAT), .Z(n388) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(n388), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n317) );
  XNOR2_X1 U360 ( .A(G43GAT), .B(G15GAT), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n313), .B(G113GAT), .ZN(n367) );
  XOR2_X1 U362 ( .A(n367), .B(KEYINPUT67), .Z(n315) );
  NAND2_X1 U363 ( .A1(G229GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U365 ( .A(n317), .B(n316), .Z(n327) );
  XOR2_X1 U366 ( .A(G50GAT), .B(G29GAT), .Z(n319) );
  XNOR2_X1 U367 ( .A(KEYINPUT7), .B(KEYINPUT70), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U369 ( .A(n320), .B(KEYINPUT8), .Z(n322) );
  XNOR2_X1 U370 ( .A(G36GAT), .B(KEYINPUT69), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n341) );
  XOR2_X1 U372 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n324) );
  XNOR2_X1 U373 ( .A(KEYINPUT72), .B(KEYINPUT68), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n341), .B(n325), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n327), .B(n326), .ZN(n569) );
  XNOR2_X1 U377 ( .A(n569), .B(KEYINPUT73), .ZN(n553) );
  NAND2_X1 U378 ( .A1(n474), .A2(n553), .ZN(n462) );
  XOR2_X1 U379 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n329) );
  XNOR2_X1 U380 ( .A(KEYINPUT10), .B(KEYINPUT9), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U382 ( .A(n330), .B(G92GAT), .Z(n332) );
  XOR2_X1 U383 ( .A(G218GAT), .B(G162GAT), .Z(n387) );
  XNOR2_X1 U384 ( .A(G43GAT), .B(n387), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n337) );
  XOR2_X1 U386 ( .A(KEYINPUT65), .B(n333), .Z(n335) );
  NAND2_X1 U387 ( .A1(G232GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U389 ( .A(n337), .B(n336), .Z(n343) );
  XOR2_X1 U390 ( .A(G106GAT), .B(G134GAT), .Z(n339) );
  XNOR2_X1 U391 ( .A(G190GAT), .B(G99GAT), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U394 ( .A(n343), .B(n342), .ZN(n538) );
  INV_X1 U395 ( .A(n538), .ZN(n563) );
  XOR2_X1 U396 ( .A(G155GAT), .B(G78GAT), .Z(n345) );
  XNOR2_X1 U397 ( .A(G22GAT), .B(G211GAT), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U399 ( .A(G127GAT), .B(G71GAT), .Z(n347) );
  XNOR2_X1 U400 ( .A(G15GAT), .B(G183GAT), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U402 ( .A(n349), .B(n348), .Z(n354) );
  XOR2_X1 U403 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n351) );
  NAND2_X1 U404 ( .A1(G231GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U406 ( .A(KEYINPUT81), .B(n352), .ZN(n353) );
  XNOR2_X1 U407 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U408 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n356) );
  XNOR2_X1 U409 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U411 ( .A(n358), .B(n357), .Z(n362) );
  XNOR2_X1 U412 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U413 ( .A(n362), .B(n361), .ZN(n561) );
  INV_X1 U414 ( .A(n561), .ZN(n578) );
  NOR2_X1 U415 ( .A1(n563), .A2(n578), .ZN(n363) );
  XNOR2_X1 U416 ( .A(n363), .B(KEYINPUT16), .ZN(n448) );
  XOR2_X1 U417 ( .A(KEYINPUT86), .B(KEYINPUT84), .Z(n369) );
  XOR2_X1 U418 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n365) );
  NAND2_X1 U419 ( .A1(G227GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n369), .B(n368), .ZN(n371) );
  XNOR2_X1 U423 ( .A(G134GAT), .B(G127GAT), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n370), .B(KEYINPUT0), .ZN(n415) );
  XOR2_X1 U425 ( .A(n371), .B(n415), .Z(n379) );
  XOR2_X1 U426 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n373) );
  XNOR2_X1 U427 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U429 ( .A(n374), .B(G183GAT), .Z(n376) );
  XNOR2_X1 U430 ( .A(G169GAT), .B(G176GAT), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n432) );
  XNOR2_X1 U432 ( .A(n432), .B(n377), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n552) );
  INV_X1 U434 ( .A(n552), .ZN(n511) );
  XNOR2_X1 U435 ( .A(n511), .B(KEYINPUT87), .ZN(n436) );
  XOR2_X1 U436 ( .A(KEYINPUT90), .B(G211GAT), .Z(n381) );
  XNOR2_X1 U437 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U439 ( .A(G197GAT), .B(n382), .Z(n425) );
  XNOR2_X1 U440 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n383), .B(KEYINPUT2), .ZN(n414) );
  XNOR2_X1 U442 ( .A(n384), .B(n414), .ZN(n396) );
  XOR2_X1 U443 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n386) );
  XNOR2_X1 U444 ( .A(KEYINPUT24), .B(KEYINPUT89), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n392) );
  XOR2_X1 U446 ( .A(KEYINPUT88), .B(n387), .Z(n390) );
  XNOR2_X1 U447 ( .A(G50GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U449 ( .A(n392), .B(n391), .Z(n394) );
  NAND2_X1 U450 ( .A1(G228GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n425), .B(n397), .ZN(n547) );
  XNOR2_X1 U454 ( .A(KEYINPUT28), .B(n547), .ZN(n514) );
  XOR2_X1 U455 ( .A(G162GAT), .B(G148GAT), .Z(n399) );
  XNOR2_X1 U456 ( .A(G113GAT), .B(G141GAT), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U458 ( .A(G29GAT), .B(G85GAT), .Z(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n421) );
  XOR2_X1 U460 ( .A(KEYINPUT99), .B(KEYINPUT97), .Z(n403) );
  XNOR2_X1 U461 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U463 ( .A(KEYINPUT96), .B(KEYINPUT94), .Z(n405) );
  XNOR2_X1 U464 ( .A(G120GAT), .B(KEYINPUT95), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(n406), .ZN(n419) );
  XOR2_X1 U467 ( .A(KEYINPUT4), .B(G57GAT), .Z(n409) );
  XNOR2_X1 U468 ( .A(KEYINPUT98), .B(KEYINPUT93), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U470 ( .A(KEYINPUT1), .B(KEYINPUT92), .Z(n411) );
  XNOR2_X1 U471 ( .A(KEYINPUT6), .B(KEYINPUT91), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U473 ( .A(n413), .B(n412), .Z(n417) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n423) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n545) );
  XOR2_X1 U480 ( .A(n424), .B(G218GAT), .Z(n427) );
  XNOR2_X1 U481 ( .A(G36GAT), .B(n425), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U483 ( .A(KEYINPUT100), .B(KEYINPUT81), .Z(n429) );
  NAND2_X1 U484 ( .A1(G226GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U486 ( .A(n431), .B(n430), .Z(n434) );
  XNOR2_X1 U487 ( .A(G8GAT), .B(n432), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n541) );
  XOR2_X1 U489 ( .A(n541), .B(KEYINPUT27), .Z(n441) );
  NAND2_X1 U490 ( .A1(n545), .A2(n441), .ZN(n510) );
  NOR2_X1 U491 ( .A1(n514), .A2(n510), .ZN(n435) );
  NAND2_X1 U492 ( .A1(n436), .A2(n435), .ZN(n447) );
  INV_X1 U493 ( .A(n545), .ZN(n445) );
  XOR2_X1 U494 ( .A(KEYINPUT101), .B(KEYINPUT25), .Z(n439) );
  NOR2_X1 U495 ( .A1(n552), .A2(n541), .ZN(n437) );
  NOR2_X1 U496 ( .A1(n547), .A2(n437), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n443) );
  NAND2_X1 U498 ( .A1(n547), .A2(n552), .ZN(n440) );
  XOR2_X1 U499 ( .A(n440), .B(KEYINPUT26), .Z(n567) );
  NAND2_X1 U500 ( .A1(n441), .A2(n567), .ZN(n442) );
  NAND2_X1 U501 ( .A1(n443), .A2(n442), .ZN(n444) );
  NAND2_X1 U502 ( .A1(n445), .A2(n444), .ZN(n446) );
  NAND2_X1 U503 ( .A1(n447), .A2(n446), .ZN(n459) );
  NAND2_X1 U504 ( .A1(n448), .A2(n459), .ZN(n475) );
  NOR2_X1 U505 ( .A1(n462), .A2(n475), .ZN(n456) );
  NAND2_X1 U506 ( .A1(n456), .A2(n545), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U508 ( .A(G1GAT), .B(n451), .Z(G1324GAT) );
  XOR2_X1 U509 ( .A(G8GAT), .B(KEYINPUT103), .Z(n453) );
  INV_X1 U510 ( .A(n541), .ZN(n489) );
  NAND2_X1 U511 ( .A1(n456), .A2(n489), .ZN(n452) );
  XNOR2_X1 U512 ( .A(n453), .B(n452), .ZN(G1325GAT) );
  XOR2_X1 U513 ( .A(G15GAT), .B(KEYINPUT35), .Z(n455) );
  NAND2_X1 U514 ( .A1(n456), .A2(n511), .ZN(n454) );
  XNOR2_X1 U515 ( .A(n455), .B(n454), .ZN(G1326GAT) );
  NAND2_X1 U516 ( .A1(n456), .A2(n514), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n457), .B(KEYINPUT104), .ZN(n458) );
  XNOR2_X1 U518 ( .A(G22GAT), .B(n458), .ZN(G1327GAT) );
  XOR2_X1 U519 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n465) );
  XOR2_X1 U520 ( .A(KEYINPUT36), .B(n538), .Z(n581) );
  NAND2_X1 U521 ( .A1(n581), .A2(n459), .ZN(n460) );
  NOR2_X1 U522 ( .A1(n561), .A2(n460), .ZN(n461) );
  XNOR2_X1 U523 ( .A(KEYINPUT37), .B(n461), .ZN(n487) );
  NOR2_X1 U524 ( .A1(n487), .A2(n462), .ZN(n463) );
  XNOR2_X1 U525 ( .A(KEYINPUT38), .B(n463), .ZN(n471) );
  NAND2_X1 U526 ( .A1(n545), .A2(n471), .ZN(n464) );
  XNOR2_X1 U527 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U528 ( .A(G29GAT), .B(n466), .Z(G1328GAT) );
  NAND2_X1 U529 ( .A1(n471), .A2(n489), .ZN(n467) );
  XNOR2_X1 U530 ( .A(n467), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U531 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n469) );
  NAND2_X1 U532 ( .A1(n471), .A2(n511), .ZN(n468) );
  XNOR2_X1 U533 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U534 ( .A(G43GAT), .B(n470), .Z(G1330GAT) );
  NAND2_X1 U535 ( .A1(n471), .A2(n514), .ZN(n472) );
  XNOR2_X1 U536 ( .A(n472), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n477) );
  INV_X1 U538 ( .A(KEYINPUT41), .ZN(n473) );
  XNOR2_X1 U539 ( .A(n474), .B(n473), .ZN(n530) );
  INV_X1 U540 ( .A(n530), .ZN(n558) );
  NAND2_X1 U541 ( .A1(n569), .A2(n558), .ZN(n486) );
  NOR2_X1 U542 ( .A1(n486), .A2(n475), .ZN(n482) );
  NAND2_X1 U543 ( .A1(n482), .A2(n545), .ZN(n476) );
  XNOR2_X1 U544 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U545 ( .A(G57GAT), .B(n478), .ZN(G1332GAT) );
  NAND2_X1 U546 ( .A1(n489), .A2(n482), .ZN(n479) );
  XNOR2_X1 U547 ( .A(n479), .B(KEYINPUT108), .ZN(n480) );
  XNOR2_X1 U548 ( .A(G64GAT), .B(n480), .ZN(G1333GAT) );
  NAND2_X1 U549 ( .A1(n511), .A2(n482), .ZN(n481) );
  XNOR2_X1 U550 ( .A(n481), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n484) );
  NAND2_X1 U552 ( .A1(n482), .A2(n514), .ZN(n483) );
  XNOR2_X1 U553 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U554 ( .A(G78GAT), .B(n485), .Z(G1335GAT) );
  NOR2_X1 U555 ( .A1(n487), .A2(n486), .ZN(n492) );
  NAND2_X1 U556 ( .A1(n545), .A2(n492), .ZN(n488) );
  XNOR2_X1 U557 ( .A(G85GAT), .B(n488), .ZN(G1336GAT) );
  NAND2_X1 U558 ( .A1(n489), .A2(n492), .ZN(n490) );
  XNOR2_X1 U559 ( .A(n490), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U560 ( .A1(n511), .A2(n492), .ZN(n491) );
  XNOR2_X1 U561 ( .A(n491), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n494) );
  NAND2_X1 U563 ( .A1(n492), .A2(n514), .ZN(n493) );
  XNOR2_X1 U564 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U565 ( .A(G106GAT), .B(n495), .Z(G1339GAT) );
  XOR2_X1 U566 ( .A(G113GAT), .B(KEYINPUT115), .Z(n516) );
  NOR2_X1 U567 ( .A1(n530), .A2(n569), .ZN(n498) );
  INV_X1 U568 ( .A(KEYINPUT46), .ZN(n496) );
  NOR2_X1 U569 ( .A1(n499), .A2(n561), .ZN(n500) );
  XNOR2_X1 U570 ( .A(n500), .B(KEYINPUT112), .ZN(n501) );
  NAND2_X1 U571 ( .A1(n501), .A2(n538), .ZN(n502) );
  XNOR2_X1 U572 ( .A(n502), .B(KEYINPUT47), .ZN(n508) );
  NAND2_X1 U573 ( .A1(n561), .A2(n581), .ZN(n504) );
  XNOR2_X1 U574 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n503) );
  XNOR2_X1 U575 ( .A(n504), .B(n503), .ZN(n505) );
  NAND2_X1 U576 ( .A1(n505), .A2(n474), .ZN(n506) );
  NOR2_X1 U577 ( .A1(n553), .A2(n506), .ZN(n507) );
  XNOR2_X1 U578 ( .A(n509), .B(KEYINPUT48), .ZN(n540) );
  NOR2_X1 U579 ( .A1(n540), .A2(n510), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n527), .A2(n511), .ZN(n512) );
  XNOR2_X1 U581 ( .A(KEYINPUT114), .B(n512), .ZN(n513) );
  NOR2_X1 U582 ( .A1(n514), .A2(n513), .ZN(n523) );
  NAND2_X1 U583 ( .A1(n523), .A2(n553), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(G1340GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n518) );
  NAND2_X1 U586 ( .A1(n523), .A2(n558), .ZN(n517) );
  XNOR2_X1 U587 ( .A(n518), .B(n517), .ZN(n520) );
  XOR2_X1 U588 ( .A(G120GAT), .B(KEYINPUT116), .Z(n519) );
  XNOR2_X1 U589 ( .A(n520), .B(n519), .ZN(G1341GAT) );
  NAND2_X1 U590 ( .A1(n523), .A2(n561), .ZN(n521) );
  XNOR2_X1 U591 ( .A(n521), .B(KEYINPUT50), .ZN(n522) );
  XNOR2_X1 U592 ( .A(G127GAT), .B(n522), .ZN(G1342GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n525) );
  NAND2_X1 U594 ( .A1(n523), .A2(n563), .ZN(n524) );
  XNOR2_X1 U595 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U596 ( .A(G134GAT), .B(n526), .ZN(G1343GAT) );
  NAND2_X1 U597 ( .A1(n527), .A2(n567), .ZN(n537) );
  NOR2_X1 U598 ( .A1(n569), .A2(n537), .ZN(n529) );
  XNOR2_X1 U599 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n528) );
  XNOR2_X1 U600 ( .A(n529), .B(n528), .ZN(G1344GAT) );
  NOR2_X1 U601 ( .A1(n530), .A2(n537), .ZN(n535) );
  XOR2_X1 U602 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n532) );
  XNOR2_X1 U603 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n531) );
  XNOR2_X1 U604 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U605 ( .A(KEYINPUT120), .B(n533), .ZN(n534) );
  XNOR2_X1 U606 ( .A(n535), .B(n534), .ZN(G1345GAT) );
  NOR2_X1 U607 ( .A1(n578), .A2(n537), .ZN(n536) );
  XOR2_X1 U608 ( .A(G155GAT), .B(n536), .Z(G1346GAT) );
  NOR2_X1 U609 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U610 ( .A(G162GAT), .B(n539), .Z(G1347GAT) );
  INV_X1 U611 ( .A(KEYINPUT54), .ZN(n543) );
  NOR2_X1 U612 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U613 ( .A(n543), .B(n542), .ZN(n544) );
  NOR2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(KEYINPUT64), .B(n546), .ZN(n568) );
  INV_X1 U616 ( .A(n568), .ZN(n548) );
  XNOR2_X1 U617 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n564), .A2(n553), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n556) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT123), .B(n557), .Z(n560) );
  NAND2_X1 U625 ( .A1(n564), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n564), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1351GAT) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n580) );
  NOR2_X1 U633 ( .A1(n569), .A2(n580), .ZN(n574) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n571) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT59), .B(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n474), .A2(n580), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n580), .ZN(n579) );
  XOR2_X1 U644 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  INV_X1 U645 ( .A(n580), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

