//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G87), .A2(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n217), .B1(new_n202), .B2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n216), .B(new_n219), .C1(G107), .C2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G116), .A2(G270), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n210), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n208), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT65), .Z(new_n235));
  NAND2_X1  g0035(.A1(new_n228), .A2(new_n214), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G50), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n213), .B(new_n232), .C1(new_n235), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G222), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n259), .B(new_n261), .C1(new_n262), .C2(new_n260), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G41), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G1), .A3(G13), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n263), .B(new_n266), .C1(G77), .C2(new_n259), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT66), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT66), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n270), .B(new_n207), .C1(G41), .C2(G45), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n269), .A2(G274), .A3(new_n265), .A4(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT67), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n265), .A2(new_n273), .A3(new_n268), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n265), .B2(new_n268), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n267), .B(new_n272), .C1(new_n224), .C2(new_n276), .ZN(new_n277));
  OR2_X1    g0077(.A1(new_n277), .A2(G179), .ZN(new_n278));
  OAI21_X1  g0078(.A(G20), .B1(new_n236), .B2(G50), .ZN(new_n279));
  INV_X1    g0079(.A(G150), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n208), .A2(G33), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  OAI221_X1 g0084(.A(new_n279), .B1(new_n280), .B2(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n286), .A2(KEYINPUT68), .A3(new_n233), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT68), .B1(new_n286), .B2(new_n233), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n285), .A2(new_n289), .B1(new_n223), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n289), .A2(new_n291), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT69), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(new_n208), .B2(G1), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n207), .A2(KEYINPUT69), .A3(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n293), .A2(G50), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n277), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n278), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n300), .B(KEYINPUT9), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT71), .ZN(new_n306));
  INV_X1    g0106(.A(G190), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n277), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n277), .A2(G200), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OR3_X1    g0111(.A1(new_n309), .A2(KEYINPUT10), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT10), .B1(new_n309), .B2(new_n311), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n304), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n229), .A2(G1698), .ZN(new_n315));
  AND2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n315), .B1(G226), .B2(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n266), .ZN(new_n321));
  OAI21_X1  g0121(.A(G238), .B1(new_n274), .B2(new_n275), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(new_n322), .A3(new_n272), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT13), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n321), .A2(new_n325), .A3(new_n322), .A4(new_n272), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(new_n307), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n214), .A2(G20), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n329), .B1(new_n283), .B2(new_n225), .C1(new_n282), .C2(new_n223), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n289), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT11), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n286), .A2(new_n233), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n297), .A2(new_n291), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n207), .A2(G13), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT12), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  OR3_X1    g0136(.A1(new_n329), .A2(new_n335), .A3(KEYINPUT12), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n334), .A2(G68), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n324), .B2(new_n326), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n328), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n327), .A2(new_n343), .A3(G169), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT14), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n327), .A2(new_n343), .A3(new_n346), .A4(G169), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n345), .B(new_n347), .C1(new_n348), .C2(new_n327), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n342), .B1(new_n349), .B2(new_n339), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n260), .A2(G232), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n259), .B(new_n351), .C1(new_n215), .C2(new_n260), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n352), .B(new_n266), .C1(G107), .C2(new_n259), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(new_n272), .C1(new_n226), .C2(new_n276), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n301), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n334), .A2(G77), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT15), .B(G87), .Z(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n283), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n284), .A2(new_n282), .B1(new_n208), .B2(new_n225), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n333), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n356), .B(new_n361), .C1(G77), .C2(new_n290), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT70), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n354), .A2(G179), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT70), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n355), .A2(new_n366), .A3(new_n362), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n354), .A2(new_n307), .ZN(new_n370));
  AOI211_X1 g0170(.A(new_n362), .B(new_n370), .C1(G200), .C2(new_n354), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n257), .A2(new_n208), .A3(new_n258), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n258), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n214), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n228), .A2(new_n214), .ZN(new_n379));
  NOR2_X1   g0179(.A1(G58), .A2(G68), .ZN(new_n380));
  OAI21_X1  g0180(.A(G20), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n281), .A2(G159), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n373), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT74), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n376), .A2(KEYINPUT73), .A3(new_n377), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n377), .A2(KEYINPUT73), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(G68), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n383), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT74), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(new_n373), .C1(new_n378), .C2(new_n383), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n385), .A2(new_n390), .A3(new_n333), .A4(new_n392), .ZN(new_n393));
  OR3_X1    g0193(.A1(new_n297), .A2(new_n284), .A3(KEYINPUT75), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT75), .B1(new_n297), .B2(new_n284), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n293), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n284), .A2(new_n291), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n265), .A2(G232), .A3(new_n268), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n272), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n262), .A2(new_n260), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n224), .A2(G1698), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n316), .C2(new_n317), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n265), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(G200), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n401), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n404), .A2(new_n405), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n266), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(G190), .A3(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n393), .A2(new_n399), .A3(new_n407), .A4(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT17), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n393), .A2(new_n399), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n410), .A2(new_n348), .A3(new_n272), .A4(new_n400), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT76), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT76), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n408), .A2(new_n418), .A3(new_n348), .A4(new_n410), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n301), .B1(new_n401), .B2(new_n406), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n415), .A2(KEYINPUT18), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT18), .B1(new_n415), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n414), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n314), .A2(new_n350), .A3(new_n372), .A4(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT23), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n208), .B2(G107), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G116), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n208), .B(G87), .C1(new_n316), .C2(new_n317), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT87), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT22), .ZN(new_n436));
  OAI221_X1 g0236(.A(new_n432), .B1(new_n433), .B2(new_n283), .C1(new_n434), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n435), .A2(KEYINPUT22), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n434), .A2(new_n439), .A3(new_n436), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(KEYINPUT24), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT24), .ZN(new_n442));
  INV_X1    g0242(.A(new_n440), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n437), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n333), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(KEYINPUT88), .B(KEYINPUT25), .C1(new_n290), .C2(G107), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n256), .B2(G1), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n207), .A2(KEYINPUT78), .A3(G33), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n290), .B(new_n450), .C1(new_n287), .C2(new_n288), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G107), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n445), .A2(new_n446), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n207), .A2(G45), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(G274), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n459));
  OR2_X1    g0259(.A1(KEYINPUT5), .A2(G41), .ZN(new_n460));
  NAND2_X1  g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT80), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(G274), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n218), .A2(G1698), .ZN(new_n466));
  OAI221_X1 g0266(.A(new_n466), .B1(G250), .B2(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G294), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n266), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n462), .A2(new_n266), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G264), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n465), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT89), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n465), .A2(new_n470), .A3(KEYINPUT89), .A4(new_n472), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n307), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n340), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OR2_X1    g0279(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n480));
  NAND2_X1  g0280(.A1(KEYINPUT88), .A2(KEYINPUT25), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n291), .A2(new_n203), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n454), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n445), .A2(new_n482), .A3(new_n446), .A4(new_n453), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n301), .B1(new_n475), .B2(new_n476), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n473), .A2(new_n348), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n333), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n450), .A2(new_n489), .A3(G116), .A4(new_n290), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n207), .A2(new_n433), .A3(G13), .A4(G20), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n286), .A2(new_n233), .B1(G20), .B2(new_n433), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G283), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n493), .B(new_n208), .C1(G33), .C2(new_n202), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n492), .A2(KEYINPUT20), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT20), .B1(new_n492), .B2(new_n494), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n490), .B(new_n491), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n471), .A2(G270), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G264), .A2(G1698), .ZN(new_n499));
  OAI221_X1 g0299(.A(new_n499), .B1(new_n218), .B2(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(new_n266), .C1(G303), .C2(new_n259), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n465), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n497), .B1(new_n502), .B2(G190), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n465), .A2(new_n498), .A3(new_n501), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G200), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(KEYINPUT86), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT86), .ZN(new_n507));
  INV_X1    g0307(.A(new_n505), .ZN(new_n508));
  INV_X1    g0308(.A(new_n497), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n504), .B2(new_n307), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n504), .A2(G169), .A3(new_n497), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n504), .A2(KEYINPUT21), .A3(G169), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n465), .A2(G179), .A3(new_n498), .A4(new_n501), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT85), .B1(new_n518), .B2(new_n497), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT85), .ZN(new_n520));
  AOI211_X1 g0320(.A(new_n520), .B(new_n509), .C1(new_n516), .C2(new_n517), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n512), .B(new_n515), .C1(new_n519), .C2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n458), .A2(KEYINPUT80), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n463), .B1(new_n462), .B2(G274), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n455), .A2(new_n457), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n265), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n524), .A2(new_n525), .B1(new_n527), .B2(new_n218), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT81), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n465), .B(KEYINPUT81), .C1(new_n218), .C2(new_n527), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n260), .A2(KEYINPUT4), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n259), .A2(G244), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n316), .A2(new_n317), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n226), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n493), .B(new_n533), .C1(new_n535), .C2(KEYINPUT4), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n259), .A2(G250), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n260), .B1(new_n537), .B2(KEYINPUT4), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n266), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n530), .A2(new_n531), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G200), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n459), .A2(new_n464), .B1(new_n471), .B2(G257), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G190), .ZN(new_n544));
  NAND2_X1  g0344(.A1(KEYINPUT6), .A2(G97), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT77), .B1(new_n545), .B2(G107), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT77), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n547), .A2(new_n203), .A3(KEYINPUT6), .A4(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G97), .A2(G107), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT6), .B1(new_n204), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI22_X1  g0352(.A1(new_n552), .A2(new_n208), .B1(new_n225), .B2(new_n282), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n203), .B1(new_n376), .B2(new_n377), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n333), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n291), .A2(G97), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n451), .B2(G97), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(KEYINPUT79), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT79), .ZN(new_n559));
  AOI211_X1 g0359(.A(new_n559), .B(new_n556), .C1(new_n451), .C2(G97), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n541), .A2(new_n544), .A3(new_n555), .A4(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n530), .A2(new_n531), .A3(new_n348), .A4(new_n539), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n539), .A2(new_n542), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n301), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n555), .B1(new_n558), .B2(new_n560), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT84), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n226), .A2(G1698), .ZN(new_n570));
  OAI221_X1 g0370(.A(new_n570), .B1(G238), .B2(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G116), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n265), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(G274), .B1(KEYINPUT82), .B2(G250), .ZN(new_n574));
  OR2_X1    g0374(.A1(new_n574), .A2(new_n456), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT82), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n456), .A2(new_n576), .A3(G250), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n266), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n569), .B1(new_n579), .B2(G190), .ZN(new_n580));
  NOR4_X1   g0380(.A1(new_n573), .A2(new_n578), .A3(KEYINPUT84), .A4(new_n307), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n283), .B2(new_n202), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT83), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n259), .A2(new_n208), .A3(G68), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n208), .B1(new_n319), .B2(new_n583), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G87), .B2(new_n204), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT83), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n589), .B(new_n583), .C1(new_n283), .C2(new_n202), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n585), .A2(new_n586), .A3(new_n588), .A4(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n591), .A2(new_n333), .B1(new_n291), .B2(new_n358), .ZN(new_n592));
  OAI21_X1  g0392(.A(G200), .B1(new_n573), .B2(new_n578), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n452), .A2(G87), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n452), .A2(new_n357), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n575), .A2(new_n577), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n265), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n571), .A2(new_n572), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(new_n265), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n592), .A2(new_n596), .B1(new_n600), .B2(new_n301), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n579), .A2(new_n348), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n582), .A2(new_n595), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n568), .A2(new_n604), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n428), .A2(new_n488), .A3(new_n523), .A4(new_n605), .ZN(G372));
  NAND2_X1  g0406(.A1(new_n312), .A2(new_n313), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n412), .B(KEYINPUT17), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n349), .A2(new_n339), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n368), .A2(KEYINPUT91), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT91), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n364), .A2(new_n612), .A3(new_n365), .A4(new_n367), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n342), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n608), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n424), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n415), .A2(KEYINPUT18), .A3(new_n422), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n607), .B1(new_n619), .B2(KEYINPUT92), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT92), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n615), .B2(new_n618), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n303), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n625));
  XOR2_X1   g0425(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n603), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT26), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n592), .A2(new_n596), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n600), .A2(new_n301), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n602), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n579), .A2(G190), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n628), .B1(new_n567), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n627), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n634), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n483), .A2(new_n567), .A3(new_n562), .A4(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n518), .A2(new_n497), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n515), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n475), .A2(new_n476), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G169), .ZN(new_n642));
  INV_X1    g0442(.A(new_n486), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n640), .B1(new_n644), .B2(new_n484), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n636), .B(new_n631), .C1(new_n638), .C2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n624), .B1(new_n427), .B2(new_n647), .ZN(G369));
  NAND3_X1  g0448(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(G343), .ZN(new_n653));
  XOR2_X1   g0453(.A(new_n653), .B(KEYINPUT93), .Z(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(new_n509), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n640), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n522), .B2(new_n655), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n483), .A2(new_n487), .ZN(new_n658));
  INV_X1    g0458(.A(new_n654), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n484), .ZN(new_n660));
  OAI22_X1  g0460(.A1(new_n658), .A2(new_n660), .B1(new_n487), .B2(new_n654), .ZN(new_n661));
  XNOR2_X1  g0461(.A(KEYINPUT94), .B(G330), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n657), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n515), .B1(new_n519), .B2(new_n521), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(new_n654), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n454), .A2(new_n482), .B1(new_n642), .B2(new_n643), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n666), .A2(new_n488), .B1(new_n667), .B2(new_n654), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT95), .Z(G399));
  INV_X1    g0470(.A(new_n211), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n237), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT29), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT99), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n665), .A2(new_n667), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n638), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n568), .A2(new_n634), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n487), .B(new_n515), .C1(new_n519), .C2(new_n521), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT99), .A4(new_n483), .ZN(new_n684));
  INV_X1    g0484(.A(new_n626), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n604), .B2(new_n567), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n637), .A2(new_n625), .A3(KEYINPUT26), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n686), .A2(new_n687), .B1(new_n602), .B2(new_n601), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n681), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n678), .B1(new_n689), .B2(new_n654), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT98), .B1(new_n646), .B2(new_n654), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n646), .A2(KEYINPUT98), .A3(new_n654), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n690), .B1(new_n678), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n523), .A2(new_n605), .A3(new_n488), .A4(new_n654), .ZN(new_n696));
  INV_X1    g0496(.A(new_n517), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n579), .A2(new_n470), .A3(new_n472), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n543), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT96), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n543), .A2(new_n697), .A3(new_n703), .A4(new_n698), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n540), .A2(new_n348), .A3(new_n473), .A4(new_n504), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n702), .B(new_n704), .C1(new_n579), .C2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT97), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n659), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT97), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n706), .A2(new_n712), .A3(KEYINPUT31), .A4(new_n659), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n696), .A2(new_n708), .A3(new_n711), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n662), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n695), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n677), .B1(new_n717), .B2(G1), .ZN(G364));
  NOR2_X1   g0518(.A1(G13), .A2(G33), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G20), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n657), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n671), .A2(new_n534), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT100), .Z(new_n725));
  AOI22_X1  g0525(.A1(new_n725), .A2(G355), .B1(new_n433), .B2(new_n671), .ZN(new_n726));
  XOR2_X1   g0526(.A(new_n726), .B(KEYINPUT101), .Z(new_n727));
  NOR2_X1   g0527(.A1(new_n671), .A2(new_n259), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G45), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(new_n238), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(new_n250), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n233), .B1(G20), .B2(new_n301), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n721), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G13), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G45), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n673), .A2(G1), .A3(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n208), .A2(new_n348), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(G317), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(KEYINPUT33), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n745), .A2(KEYINPUT33), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n743), .A2(new_n307), .ZN(new_n749));
  XOR2_X1   g0549(.A(KEYINPUT104), .B(G326), .Z(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G294), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n307), .A2(G200), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n208), .B1(new_n753), .B2(new_n348), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n748), .B(new_n751), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT102), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n742), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(KEYINPUT102), .B1(new_n208), .B2(new_n348), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G190), .A2(G200), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT103), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n755), .B1(G311), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n208), .A2(G179), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n307), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(G283), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n534), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n763), .A2(new_n759), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n766), .B1(G329), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n762), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G303), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n757), .A2(new_n753), .A3(new_n758), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n770), .B1(new_n771), .B2(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n764), .A2(new_n203), .ZN(new_n776));
  INV_X1    g0576(.A(new_n772), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n777), .A2(G87), .ZN(new_n778));
  INV_X1    g0578(.A(new_n774), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n778), .B1(new_n779), .B2(G58), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n749), .A2(G50), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n754), .A2(new_n202), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n767), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n780), .A2(new_n781), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G68), .B2(new_n744), .ZN(new_n788));
  INV_X1    g0588(.A(new_n761), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n788), .B(new_n259), .C1(new_n225), .C2(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n775), .B1(new_n776), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n734), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n723), .A2(new_n736), .A3(new_n741), .A4(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n657), .A2(new_n662), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n657), .A2(new_n662), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n794), .A2(new_n795), .A3(new_n740), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n793), .A2(new_n796), .ZN(G396));
  NAND3_X1  g0597(.A1(new_n646), .A2(new_n372), .A3(new_n654), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n611), .A2(new_n362), .A3(new_n613), .A4(new_n659), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n659), .A2(new_n362), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n369), .B2(new_n371), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n798), .B1(new_n694), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(new_n715), .Z(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n740), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n259), .B1(new_n754), .B2(new_n228), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n761), .A2(G159), .B1(G150), .B2(new_n744), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  INV_X1    g0608(.A(new_n749), .ZN(new_n809));
  INV_X1    g0609(.A(G143), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n807), .B1(new_n808), .B2(new_n809), .C1(new_n810), .C2(new_n774), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n777), .A2(G50), .ZN(new_n813));
  INV_X1    g0613(.A(new_n764), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G68), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n806), .B(new_n816), .C1(G132), .C2(new_n768), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n534), .B1(new_n767), .B2(new_n818), .C1(new_n809), .C2(new_n771), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n782), .B(new_n819), .C1(G107), .C2(new_n777), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n761), .A2(G116), .B1(G87), .B2(new_n814), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(new_n752), .C2(new_n774), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G283), .B2(new_n744), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n734), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n734), .A2(new_n719), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n824), .B(new_n741), .C1(G77), .C2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT105), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n802), .A2(new_n720), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n805), .B1(new_n828), .B2(new_n829), .ZN(G384));
  NAND3_X1  g0630(.A1(new_n696), .A2(new_n711), .A3(new_n707), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n802), .ZN(new_n832));
  INV_X1    g0632(.A(new_n339), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n654), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  MUX2_X1   g0635(.A(new_n349), .B(new_n350), .S(new_n835), .Z(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT38), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT106), .ZN(new_n840));
  INV_X1    g0640(.A(new_n289), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n388), .A2(new_n389), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n842), .B2(new_n373), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n398), .B1(new_n843), .B2(new_n390), .ZN(new_n844));
  INV_X1    g0644(.A(new_n652), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n840), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n388), .A2(KEYINPUT16), .A3(new_n389), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT16), .B1(new_n388), .B2(new_n389), .ZN(new_n848));
  NOR3_X1   g0648(.A1(new_n847), .A2(new_n848), .A3(new_n841), .ZN(new_n849));
  OAI211_X1 g0649(.A(KEYINPUT106), .B(new_n652), .C1(new_n849), .C2(new_n398), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n618), .B2(new_n608), .ZN(new_n852));
  INV_X1    g0652(.A(new_n412), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n393), .A2(new_n399), .B1(new_n421), .B2(new_n845), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n853), .A2(KEYINPUT37), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n422), .B1(new_n849), .B2(new_n398), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n846), .A2(new_n850), .A3(new_n412), .A4(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n855), .B1(new_n857), .B2(KEYINPUT37), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n839), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n860));
  INV_X1    g0660(.A(new_n855), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n846), .A2(new_n850), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n414), .B2(new_n425), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n838), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT40), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n853), .A2(new_n854), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n415), .A2(new_n652), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n618), .B2(new_n608), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n839), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT108), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT108), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n876), .B(new_n839), .C1(new_n871), .C2(new_n873), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(new_n865), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(new_n838), .A3(KEYINPUT40), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n869), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n428), .A2(new_n831), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n880), .B(new_n881), .Z(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n662), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n852), .A2(new_n858), .A3(new_n839), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n862), .B2(new_n864), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT39), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT107), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n875), .A2(new_n888), .A3(new_n865), .A4(new_n877), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT107), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n866), .A2(new_n890), .A3(KEYINPUT39), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n887), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n609), .A2(new_n659), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n369), .A2(new_n654), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n798), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n836), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n884), .A2(new_n885), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n897), .A2(new_n898), .B1(new_n618), .B2(new_n652), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n883), .B(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n693), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n678), .B1(new_n903), .B2(new_n691), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n689), .A2(new_n654), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT29), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n427), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n623), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n902), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n207), .B2(new_n738), .ZN(new_n910));
  INV_X1    g0710(.A(new_n552), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n433), .B1(new_n911), .B2(KEYINPUT35), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(new_n235), .C1(KEYINPUT35), .C2(new_n911), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT36), .ZN(new_n914));
  OAI21_X1  g0714(.A(G77), .B1(new_n228), .B2(new_n214), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n237), .A2(new_n915), .B1(G50), .B2(new_n214), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(G1), .A3(new_n737), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n910), .A2(new_n914), .A3(new_n917), .ZN(G367));
  AND2_X1   g0718(.A1(new_n592), .A2(new_n594), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n654), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(new_n631), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n637), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT109), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n488), .A2(new_n665), .A3(new_n654), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n659), .A2(new_n566), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n562), .A2(new_n567), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT42), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n567), .B1(new_n931), .B2(new_n487), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n654), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT42), .ZN(new_n935));
  INV_X1    g0735(.A(new_n931), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n666), .A2(new_n935), .A3(new_n936), .A4(new_n488), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n932), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(KEYINPUT110), .A3(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT110), .B1(new_n938), .B2(new_n939), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n928), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n942), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n927), .A3(new_n940), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n931), .B1(new_n567), .B2(new_n654), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n663), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT111), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n943), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT112), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n947), .A2(KEYINPUT111), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT112), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n943), .A2(new_n945), .A3(new_n952), .A4(new_n948), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n950), .A2(new_n953), .ZN(new_n955));
  INV_X1    g0755(.A(new_n951), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n672), .B(KEYINPUT41), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n668), .A2(new_n946), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT44), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n668), .A2(new_n946), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT45), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n961), .A2(new_n963), .A3(new_n663), .ZN(new_n964));
  INV_X1    g0764(.A(new_n963), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n960), .B(KEYINPUT44), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n664), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n929), .B1(new_n661), .B2(new_n666), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n969), .A2(KEYINPUT113), .B1(new_n662), .B2(new_n657), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT113), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n929), .B(new_n971), .C1(new_n661), .C2(new_n666), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n663), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n973), .A2(new_n715), .A3(new_n906), .A4(new_n904), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT114), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT114), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n695), .A2(new_n976), .A3(new_n715), .A4(new_n973), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT115), .ZN(new_n978));
  AND3_X1   g0778(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(new_n975), .B2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n968), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n959), .B1(new_n981), .B2(new_n717), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n739), .A2(G1), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n954), .B(new_n957), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n534), .B1(new_n202), .B2(new_n764), .C1(new_n789), .C2(new_n765), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n809), .A2(new_n818), .B1(new_n203), .B2(new_n754), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT46), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n772), .B2(new_n433), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n745), .B2(new_n767), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n772), .A2(new_n987), .A3(new_n433), .ZN(new_n990));
  NOR4_X1   g0790(.A1(new_n985), .A2(new_n986), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n744), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n991), .B1(new_n752), .B2(new_n992), .C1(new_n771), .C2(new_n774), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n772), .A2(new_n228), .B1(new_n767), .B2(new_n808), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n764), .A2(new_n225), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n534), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT116), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n994), .B(new_n997), .C1(G150), .C2(new_n779), .ZN(new_n998));
  INV_X1    g0798(.A(new_n754), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n744), .A2(G159), .B1(new_n999), .B2(G68), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n998), .B(new_n1000), .C1(new_n810), .C2(new_n809), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n789), .A2(new_n223), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n993), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT47), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n734), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n921), .A2(new_n721), .A3(new_n922), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n735), .B1(new_n211), .B2(new_n358), .C1(new_n242), .C2(new_n729), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1005), .A2(new_n741), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n984), .A2(new_n1008), .ZN(G387));
  AOI22_X1  g0809(.A1(new_n761), .A2(G68), .B1(G97), .B2(new_n814), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n259), .B1(new_n767), .B2(new_n280), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n358), .A2(new_n754), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(new_n779), .C2(G50), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n772), .A2(new_n225), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n284), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1014), .B1(new_n1015), .B2(new_n744), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n749), .A2(G159), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1010), .A2(new_n1013), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT119), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n761), .A2(G303), .B1(G311), .B2(new_n744), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n745), .B2(new_n774), .C1(new_n773), .C2(new_n809), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT48), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n765), .B2(new_n754), .C1(new_n752), .C2(new_n772), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT49), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n814), .A2(G116), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n768), .A2(new_n750), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1025), .A2(new_n534), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1019), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n740), .B1(new_n1030), .B2(new_n734), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(KEYINPUT117), .B(KEYINPUT50), .ZN(new_n1032));
  OR3_X1    g0832(.A1(new_n284), .A2(new_n1032), .A3(G50), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(new_n284), .B2(G50), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1033), .A2(new_n730), .A3(new_n674), .A4(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n214), .A2(new_n225), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n728), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT118), .Z(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n730), .B2(new_n246), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n725), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1039), .B1(G107), .B2(new_n211), .C1(new_n674), .C2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n735), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1031), .B(new_n1042), .C1(new_n661), .C2(new_n722), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n973), .A2(new_n983), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n974), .A2(KEYINPUT114), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n974), .A2(KEYINPUT114), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n672), .B1(new_n717), .B2(new_n973), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1045), .A2(new_n1048), .ZN(G393));
  OR2_X1    g0849(.A1(new_n964), .A2(new_n967), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1047), .B2(new_n1046), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n981), .A2(new_n1051), .A3(new_n672), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n968), .A2(new_n983), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n946), .A2(new_n722), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n779), .A2(G159), .B1(G150), .B2(new_n749), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT51), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G68), .B2(new_n777), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n814), .A2(G87), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n761), .A2(new_n1015), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n754), .A2(new_n225), .B1(new_n767), .B2(new_n810), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n534), .B(new_n1060), .C1(G50), .C2(new_n744), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n992), .A2(new_n771), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n767), .A2(new_n773), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n776), .B(new_n1064), .C1(new_n761), .C2(G294), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n809), .A2(new_n745), .B1(new_n818), .B2(new_n774), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n777), .A2(G283), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n259), .B1(new_n999), .B2(G116), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1062), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n734), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n735), .B1(new_n202), .B2(new_n211), .C1(new_n729), .C2(new_n253), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1054), .A2(new_n741), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1052), .A2(new_n1053), .A3(new_n1074), .ZN(G390));
  INV_X1    g0875(.A(new_n893), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n897), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n887), .A2(new_n889), .A3(new_n1077), .A4(new_n891), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n689), .A2(new_n654), .A3(new_n802), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n895), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n836), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n1076), .A3(new_n878), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n714), .A2(new_n836), .A3(new_n662), .A4(new_n802), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1078), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n836), .A2(new_n831), .A3(G330), .A4(new_n802), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(G330), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n837), .B1(new_n832), .B2(new_n1089), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1090), .A2(new_n1083), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1080), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n802), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n837), .B1(new_n715), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n1086), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1091), .A2(new_n1092), .B1(new_n1095), .B2(new_n896), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n881), .A2(new_n1089), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n904), .A2(new_n906), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n428), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n624), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1084), .B(new_n1088), .C1(new_n1102), .C2(KEYINPUT120), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1088), .A2(new_n1084), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1095), .A2(new_n896), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1092), .A2(new_n1090), .A3(new_n1083), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n623), .A2(new_n907), .A3(new_n1097), .ZN(new_n1108));
  AOI21_X1  g0908(.A(KEYINPUT120), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1103), .A2(new_n1110), .A3(new_n672), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n983), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1104), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n534), .B1(new_n992), .B2(new_n203), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n778), .B(new_n1114), .C1(G283), .C2(new_n749), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n768), .A2(G294), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n779), .A2(G116), .B1(G77), .B2(new_n999), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n761), .A2(G97), .B1(G68), .B2(new_n814), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT54), .B(G143), .Z(new_n1120));
  NAND2_X1  g0920(.A1(new_n761), .A2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n744), .A2(G137), .B1(new_n999), .B2(G159), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n749), .A2(G128), .B1(new_n814), .B2(G50), .ZN(new_n1123));
  INV_X1    g0923(.A(G125), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n259), .B1(new_n767), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n779), .B2(G132), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n777), .A2(G150), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1119), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n734), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n741), .B(new_n1131), .C1(new_n892), .C2(new_n720), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n284), .B2(new_n825), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1113), .A2(new_n1133), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1111), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(G378));
  NAND3_X1  g0936(.A1(new_n869), .A2(G330), .A3(new_n879), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n300), .A2(new_n652), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n314), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n314), .A2(new_n1143), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1139), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n314), .A2(new_n1143), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n894), .B2(new_n900), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n899), .B(new_n1150), .C1(new_n892), .C2(new_n893), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1137), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n890), .B1(new_n866), .B2(KEYINPUT39), .ZN(new_n1155));
  AOI211_X1 g0955(.A(KEYINPUT107), .B(new_n888), .C1(new_n859), .C2(new_n865), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1076), .B1(new_n1157), .B2(new_n889), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1150), .B1(new_n1158), .B2(new_n899), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1137), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n894), .A2(new_n900), .A3(new_n1151), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1088), .A2(new_n1084), .A3(new_n1107), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1154), .A2(new_n1162), .B1(new_n1108), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n673), .B1(new_n1164), .B2(KEYINPUT57), .ZN(new_n1165));
  OAI21_X1  g0965(.A(KEYINPUT123), .B1(new_n1164), .B2(KEYINPUT57), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1108), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1152), .A2(new_n1153), .A3(new_n1137), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1160), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT123), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1165), .A2(new_n1166), .A3(new_n1173), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1151), .A2(new_n720), .B1(G50), .B2(new_n826), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n749), .A2(G116), .B1(G283), .B2(new_n768), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n202), .B2(new_n992), .C1(new_n203), .C2(new_n774), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n357), .B2(new_n761), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n764), .A2(new_n228), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1014), .A2(new_n1179), .A3(G41), .A4(new_n259), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(new_n214), .C2(new_n754), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT58), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n223), .B1(new_n316), .B2(G41), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n761), .A2(G137), .B1(new_n777), .B2(new_n1120), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n744), .A2(G132), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n749), .A2(G125), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n779), .A2(G128), .B1(G150), .B2(new_n999), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  AOI21_X1  g0989(.A(G41), .B1(new_n1188), .B2(KEYINPUT59), .ZN(new_n1190));
  AOI21_X1  g0990(.A(G33), .B1(new_n768), .B2(G124), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n784), .C2(new_n764), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1182), .B(new_n1183), .C1(new_n1189), .C2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n740), .B(new_n1175), .C1(new_n734), .C2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1154), .A2(new_n1162), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n983), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1174), .A2(new_n1196), .ZN(G375));
  NAND2_X1  g0997(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n1199), .A3(new_n958), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n789), .A2(new_n280), .B1(new_n223), .B2(new_n754), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT124), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1179), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n259), .B1(new_n772), .B2(new_n784), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n768), .A2(G128), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G132), .C2(new_n749), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n779), .A2(G137), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1204), .A2(new_n1205), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1203), .B(new_n1210), .C1(new_n744), .C2(new_n1120), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n992), .A2(new_n433), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1012), .B(new_n1212), .C1(G294), .C2(new_n749), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n779), .A2(G283), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n761), .A2(G107), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n259), .B(new_n995), .C1(G303), .C2(new_n768), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G97), .B2(new_n777), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n734), .B1(new_n1211), .B2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n741), .B(new_n1219), .C1(new_n836), .C2(new_n720), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n214), .B2(new_n825), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1107), .B2(new_n983), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1200), .A2(new_n1222), .ZN(G381));
  NOR2_X1   g1023(.A1(G375), .A2(G378), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1052), .A2(new_n1053), .A3(new_n1074), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n984), .A2(new_n1225), .A3(new_n1008), .ZN(new_n1226));
  INV_X1    g1026(.A(G396), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1045), .A2(new_n1227), .A3(new_n1048), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1226), .A2(G384), .A3(G381), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1224), .A2(new_n1229), .ZN(G407));
  INV_X1    g1030(.A(G343), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1224), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(G213), .ZN(G409));
  NAND2_X1  g1033(.A1(new_n957), .A2(new_n954), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT115), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n975), .A2(new_n977), .A3(new_n978), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1050), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n958), .B1(new_n1237), .B2(new_n716), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1234), .B1(new_n1238), .B2(new_n1112), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1008), .ZN(new_n1240));
  OAI21_X1  g1040(.A(G390), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT126), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1228), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1227), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1244), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(KEYINPUT126), .A3(new_n1228), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1241), .A2(new_n1248), .A3(new_n1226), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1243), .A2(new_n1242), .A3(new_n1244), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1241), .B2(new_n1226), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1135), .B1(new_n1174), .B2(new_n1196), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n672), .B(new_n1199), .C1(new_n1198), .C2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT60), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1222), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(G384), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G384), .B(new_n1222), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(G213), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(G343), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1164), .A2(new_n958), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1135), .A2(new_n1196), .A3(new_n1264), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1253), .A2(new_n1261), .A3(new_n1263), .A4(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1253), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT125), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1261), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1263), .A2(G2897), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1261), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1261), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT125), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n1266), .A2(new_n1267), .B1(new_n1268), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1263), .B1(G375), .B2(G378), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1265), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(new_n1267), .A3(new_n1276), .A4(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT61), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1252), .B1(new_n1279), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1283), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(new_n1266), .B2(KEYINPUT63), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G375), .A2(G378), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1263), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1281), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1288), .B1(new_n1289), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1287), .B1(new_n1293), .B2(new_n1266), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1285), .A2(new_n1294), .ZN(G405));
  INV_X1    g1095(.A(KEYINPUT127), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  OR3_X1    g1098(.A1(new_n1224), .A2(new_n1276), .A3(new_n1253), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1276), .B1(new_n1224), .B2(new_n1253), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1298), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1241), .A2(new_n1248), .A3(new_n1226), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1241), .A2(new_n1226), .ZN(new_n1304));
  OAI211_X1 g1104(.A(KEYINPUT127), .B(new_n1303), .C1(new_n1304), .C2(new_n1250), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1297), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1301), .B1(new_n1302), .B2(new_n1306), .ZN(G402));
endmodule


