//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1106,
    new_n1107;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT66), .B(KEYINPUT67), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(G137), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT69), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n464), .A2(new_n475), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n463), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(G160));
  INV_X1    g055(.A(new_n464), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n463), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n463), .C2(G112), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n481), .B2(G2105), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n464), .A2(KEYINPUT70), .A3(new_n459), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n483), .B(new_n484), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n490), .B(new_n491), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT73), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n459), .B2(G114), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT73), .A3(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G102), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n459), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n494), .A2(new_n496), .A3(G2104), .A4(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n470), .A2(new_n472), .A3(G126), .A4(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(KEYINPUT74), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n463), .A2(new_n464), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n463), .A2(new_n464), .A3(new_n506), .A4(new_n503), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n501), .B1(new_n505), .B2(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(G543), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(G88), .B1(G50), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT75), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n510), .A2(new_n512), .A3(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(G651), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT76), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n522), .A2(KEYINPUT76), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n514), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n515), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n531), .A2(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G651), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n515), .A2(new_n542), .B1(new_n529), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n510), .A2(new_n512), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XOR2_X1   g127(.A(KEYINPUT79), .B(G43), .Z(new_n553));
  AOI22_X1  g128(.A1(new_n516), .A2(G81), .B1(new_n517), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  AOI211_X1 g137(.A(KEYINPUT80), .B(KEYINPUT9), .C1(new_n517), .C2(G53), .ZN(new_n563));
  XOR2_X1   g138(.A(KEYINPUT80), .B(KEYINPUT9), .Z(new_n564));
  AND3_X1   g139(.A1(new_n517), .A2(G53), .A3(new_n564), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G91), .ZN(new_n568));
  OAI22_X1  g143(.A1(new_n567), .A2(new_n540), .B1(new_n515), .B2(new_n568), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n566), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  XNOR2_X1  g146(.A(G168), .B(KEYINPUT81), .ZN(G286));
  NAND2_X1  g147(.A1(new_n516), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n517), .A2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  AOI22_X1  g151(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n540), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  INV_X1    g154(.A(G48), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n515), .A2(new_n579), .B1(new_n529), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n516), .A2(G85), .B1(G47), .B2(new_n517), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n540), .B2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n513), .A2(G92), .A3(new_n514), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n547), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(G651), .A2(new_n592), .B1(new_n517), .B2(G54), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT82), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n587), .B1(new_n595), .B2(G868), .ZN(G284));
  OAI21_X1  g171(.A(new_n587), .B1(new_n595), .B2(G868), .ZN(G321));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G299), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G297));
  XNOR2_X1  g175(.A(G297), .B(KEYINPUT83), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n595), .A2(new_n602), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n605), .A2(KEYINPUT84), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT84), .B1(new_n605), .B2(new_n606), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n607), .B(new_n608), .C1(G868), .C2(new_n556), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n464), .A2(new_n467), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n482), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n463), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  OAI221_X1 g193(.A(new_n615), .B1(new_n616), .B2(new_n617), .C1(new_n488), .C2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(G2096), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n614), .A2(new_n620), .ZN(G156));
  INV_X1    g196(.A(KEYINPUT14), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT15), .B(G2435), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2438), .ZN(new_n624));
  XOR2_X1   g199(.A(G2427), .B(G2430), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT85), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n622), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n624), .B2(new_n626), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2451), .B(G2454), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT16), .B(G1341), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  AND2_X1   g209(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(G14), .B1(new_n628), .B2(new_n634), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n635), .A2(new_n636), .ZN(G401));
  XOR2_X1   g212(.A(G2072), .B(G2078), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT17), .ZN(new_n639));
  XOR2_X1   g214(.A(G2067), .B(G2678), .Z(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT86), .Z(new_n643));
  INV_X1    g218(.A(new_n638), .ZN(new_n644));
  INV_X1    g219(.A(new_n640), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(new_n645), .A3(new_n641), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT18), .Z(new_n647));
  AOI21_X1  g222(.A(new_n641), .B1(new_n638), .B2(new_n640), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n639), .B2(new_n640), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n643), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2096), .B(G2100), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1956), .B(G2474), .Z(new_n653));
  XOR2_X1   g228(.A(G1961), .B(G1966), .Z(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n656), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n656), .A2(new_n660), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n664));
  OAI221_X1 g239(.A(new_n661), .B1(new_n660), .B2(new_n658), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n664), .B2(new_n663), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G1991), .ZN(new_n667));
  INV_X1    g242(.A(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G6), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n582), .B2(new_n674), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT89), .Z(new_n677));
  XOR2_X1   g252(.A(KEYINPUT32), .B(G1981), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NOR2_X1   g255(.A1(G16), .A2(G23), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT90), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G288), .B2(new_n674), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT33), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n674), .A2(G22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT91), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G303), .B2(G16), .ZN(new_n688));
  INV_X1    g263(.A(G1971), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR4_X1   g266(.A1(new_n679), .A2(new_n680), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT34), .ZN(new_n693));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G25), .ZN(new_n695));
  NOR2_X1   g270(.A1(G95), .A2(G2105), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT87), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT88), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n482), .A2(G119), .ZN(new_n700));
  INV_X1    g275(.A(G131), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n488), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n695), .B1(new_n703), .B2(new_n694), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT35), .B(G1991), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n708));
  MUX2_X1   g283(.A(G24), .B(G290), .S(G16), .Z(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G1986), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G1986), .B2(new_n709), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n693), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G29), .A2(G35), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G162), .B2(G29), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(G2090), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n694), .A2(G26), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n482), .A2(G128), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT93), .Z(new_n724));
  INV_X1    g299(.A(new_n488), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G140), .ZN(new_n726));
  OAI221_X1 g301(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n463), .C2(G116), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n724), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n722), .B1(new_n728), .B2(G29), .ZN(new_n729));
  MUX2_X1   g304(.A(new_n722), .B(new_n729), .S(KEYINPUT28), .Z(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT94), .B(G2067), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n720), .A2(G2090), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n721), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n674), .A2(G20), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT23), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT23), .B1(new_n599), .B2(new_n674), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(new_n735), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1956), .ZN(new_n740));
  INV_X1    g315(.A(G28), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT30), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n741), .B2(KEYINPUT30), .ZN(new_n743));
  OR2_X1    g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  NAND2_X1  g319(.A1(KEYINPUT31), .A2(G11), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n742), .A2(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n619), .B2(new_n694), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n674), .A2(G21), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G168), .B2(new_n674), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT97), .B(G1966), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G5), .A2(G16), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G171), .B2(G16), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n747), .B(new_n751), .C1(G1961), .C2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT98), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n694), .A2(G27), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G164), .B2(new_n694), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(G2078), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(G2078), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n759), .B(new_n760), .C1(G1961), .C2(new_n753), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n754), .B2(new_n755), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n674), .A2(G4), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n595), .B2(new_n674), .ZN(new_n764));
  INV_X1    g339(.A(G1348), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n740), .A2(new_n756), .A3(new_n762), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n482), .A2(G129), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT26), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n771), .A2(new_n772), .B1(G105), .B2(new_n467), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n725), .B2(G141), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G29), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT96), .Z(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G29), .B2(G32), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT27), .B(G1996), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT24), .ZN(new_n781));
  INV_X1    g356(.A(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(G29), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n781), .B2(new_n782), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G160), .B2(new_n694), .ZN(new_n785));
  INV_X1    g360(.A(G2084), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n674), .A2(G19), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n556), .B2(new_n674), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1341), .Z(new_n790));
  NAND3_X1  g365(.A1(new_n780), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n694), .A2(G33), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT25), .Z(new_n794));
  INV_X1    g369(.A(G139), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n488), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT95), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(new_n463), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n792), .B1(new_n800), .B2(new_n694), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2072), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n734), .A2(new_n767), .A3(new_n791), .A4(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n712), .A2(new_n713), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n715), .A2(new_n804), .A3(new_n805), .ZN(G311));
  INV_X1    g381(.A(G311), .ZN(G150));
  XNOR2_X1  g382(.A(KEYINPUT101), .B(G55), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n529), .A2(new_n808), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n540), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n809), .B(new_n811), .C1(G93), .C2(new_n516), .ZN(new_n812));
  INV_X1    g387(.A(G860), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT37), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n595), .A2(G559), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT39), .Z(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n812), .B(new_n555), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n813), .B1(new_n818), .B2(new_n821), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n815), .B1(new_n822), .B2(new_n823), .ZN(G145));
  XNOR2_X1  g399(.A(new_n619), .B(G160), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G162), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n827));
  INV_X1    g402(.A(new_n507), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n499), .A2(KEYINPUT102), .A3(new_n500), .ZN(new_n829));
  AOI21_X1  g404(.A(KEYINPUT102), .B1(new_n499), .B2(new_n500), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n827), .A2(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n826), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n612), .B(KEYINPUT103), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(new_n775), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n703), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n800), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n482), .A2(G130), .ZN(new_n838));
  OAI221_X1 g413(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n463), .C2(G118), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G142), .B2(new_n725), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n728), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n837), .B(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(G37), .B1(new_n835), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n843), .B2(new_n835), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(G395));
  XOR2_X1   g422(.A(G288), .B(KEYINPUT106), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G290), .ZN(new_n849));
  XNOR2_X1  g424(.A(G303), .B(G305), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(KEYINPUT42), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT107), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n851), .B(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n852), .B1(new_n854), .B2(KEYINPUT42), .ZN(new_n855));
  INV_X1    g430(.A(new_n594), .ZN(new_n856));
  OR3_X1    g431(.A1(G299), .A2(KEYINPUT105), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT105), .B1(G299), .B2(new_n856), .ZN(new_n858));
  NAND2_X1  g433(.A1(G299), .A2(new_n856), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n604), .B(new_n819), .ZN(new_n863));
  MUX2_X1   g438(.A(new_n860), .B(new_n862), .S(new_n863), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n855), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G868), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(G868), .B2(new_n812), .ZN(G295));
  XOR2_X1   g442(.A(G295), .B(KEYINPUT108), .Z(G331));
  MUX2_X1   g443(.A(G168), .B(G286), .S(G171), .Z(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(new_n819), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n819), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT109), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n871), .A2(KEYINPUT109), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n862), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT110), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n862), .B(KEYINPUT110), .C1(new_n873), .C2(new_n872), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n870), .A2(new_n860), .A3(new_n871), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n876), .A2(new_n854), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n879), .A2(KEYINPUT111), .ZN(new_n880));
  AOI21_X1  g455(.A(G37), .B1(new_n879), .B2(KEYINPUT111), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT43), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n884));
  INV_X1    g459(.A(new_n854), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n872), .A2(new_n873), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n888), .A2(new_n860), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n870), .A2(new_n871), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n862), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n885), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g468(.A(KEYINPUT44), .B(new_n887), .C1(new_n893), .C2(new_n883), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n880), .A2(new_n881), .A3(new_n886), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT43), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n880), .A2(new_n881), .A3(new_n883), .A4(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT112), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT112), .ZN(new_n901));
  AOI211_X1 g476(.A(new_n901), .B(KEYINPUT44), .C1(new_n896), .C2(new_n897), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n894), .B1(new_n900), .B2(new_n902), .ZN(G397));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n501), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n499), .A2(KEYINPUT102), .A3(new_n500), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n505), .A2(new_n507), .ZN(new_n908));
  AOI21_X1  g483(.A(G1384), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(G160), .A2(G40), .ZN(new_n910));
  XNOR2_X1  g485(.A(KEYINPUT113), .B(KEYINPUT45), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n728), .B(G2067), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n775), .B(new_n668), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n915), .B(KEYINPUT114), .Z(new_n916));
  NOR2_X1   g491(.A1(new_n836), .A2(new_n705), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n728), .A2(G2067), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n912), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n913), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n775), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n912), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n912), .A2(new_n668), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT46), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n924), .A2(KEYINPUT46), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT47), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n706), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n912), .B1(new_n917), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n916), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(G290), .A2(G1986), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n912), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n933), .B(KEYINPUT48), .Z(new_n934));
  OAI211_X1 g509(.A(new_n920), .B(new_n928), .C1(new_n931), .C2(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n935), .B(KEYINPUT127), .Z(new_n936));
  INV_X1    g511(.A(G1384), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n831), .A2(G40), .A3(G160), .A4(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G8), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n582), .B(G1981), .Z(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT49), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n941), .ZN(new_n945));
  INV_X1    g520(.A(G1976), .ZN(new_n946));
  INV_X1    g521(.A(G288), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OR2_X1    g523(.A1(G305), .A2(G1981), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n942), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n951));
  INV_X1    g526(.A(G40), .ZN(new_n952));
  AOI211_X1 g527(.A(new_n952), .B(new_n469), .C1(new_n479), .C2(new_n478), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n831), .A2(new_n955), .A3(new_n937), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n957), .A2(G2090), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT115), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n910), .B1(new_n909), .B2(KEYINPUT45), .ZN(new_n960));
  NOR2_X1   g535(.A1(G164), .A2(G1384), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n961), .A2(new_n911), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n958), .A2(new_n959), .B1(new_n689), .B2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n959), .B2(new_n958), .ZN(new_n965));
  NAND2_X1  g540(.A1(G303), .A2(G8), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT55), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(G8), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n942), .B1(G1976), .B2(new_n947), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n945), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT52), .B1(G288), .B2(new_n946), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n950), .B1(new_n970), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n975), .A2(new_n969), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n953), .B1(new_n909), .B2(new_n955), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n961), .A2(new_n955), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n983), .A2(G2090), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n963), .A2(new_n689), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n940), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n977), .B1(new_n968), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(G160), .A2(KEYINPUT45), .A3(G40), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n938), .A2(KEYINPUT117), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n961), .A2(new_n911), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT117), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n992), .B(new_n953), .C1(new_n909), .C2(KEYINPUT45), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1966), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AND4_X1   g571(.A1(new_n786), .A2(new_n956), .A3(new_n953), .A4(new_n951), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n940), .B(G286), .C1(new_n996), .C2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT63), .B1(new_n988), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n965), .A2(G8), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n967), .ZN(new_n1002));
  AND4_X1   g577(.A1(KEYINPUT63), .A2(new_n977), .A3(new_n999), .A4(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n976), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT125), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G168), .A2(new_n940), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT123), .B1(new_n996), .B2(new_n998), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT123), .ZN(new_n1009));
  AOI211_X1 g584(.A(new_n1009), .B(new_n997), .C1(new_n994), .C2(new_n995), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1008), .A2(new_n1010), .A3(new_n940), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT124), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1007), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n996), .A2(new_n998), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n1009), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n996), .A2(KEYINPUT123), .A3(new_n998), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1015), .A2(new_n1012), .A3(new_n1016), .A4(G8), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT51), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT51), .B(new_n1006), .C1(new_n1014), .C2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1008), .A2(new_n1010), .A3(new_n1007), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1005), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1015), .A2(G8), .A3(new_n1016), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT124), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n1017), .A3(new_n1007), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1020), .B1(new_n1028), .B2(KEYINPUT51), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1029), .A2(KEYINPUT125), .A3(new_n1023), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT62), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1022), .A2(new_n1005), .A3(new_n1024), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT125), .B1(new_n1029), .B2(new_n1023), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT62), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n963), .B2(G2078), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n954), .A2(new_n956), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(G1961), .B2(new_n1038), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n994), .A2(G2078), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1040), .A2(KEYINPUT126), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1036), .B1(new_n1040), .B2(KEYINPUT126), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(G301), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1031), .A2(new_n1035), .A3(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(G171), .B(KEYINPUT54), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1036), .A2(G2078), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n960), .B(new_n1047), .C1(new_n909), .C2(new_n911), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1046), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1043), .A2(new_n1046), .B1(new_n1039), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT56), .B(G2072), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n960), .A2(new_n962), .A3(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1052), .B(KEYINPUT118), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(G299), .B(KEYINPUT57), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1956), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n983), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT61), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1058), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1055), .B1(new_n1063), .B2(new_n1053), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1054), .A2(KEYINPUT119), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1059), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(KEYINPUT120), .A3(new_n1055), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1067), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1066), .B1(new_n1072), .B2(new_n1062), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n938), .A2(G2067), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n957), .B2(new_n765), .ZN(new_n1075));
  INV_X1    g650(.A(new_n595), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT122), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1077), .A2(new_n1082), .A3(new_n1079), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1081), .A2(KEYINPUT60), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT60), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n960), .A2(new_n668), .A3(new_n962), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  NAND2_X1  g662(.A1(new_n938), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n555), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1090));
  XOR2_X1   g665(.A(new_n1089), .B(new_n1090), .Z(new_n1091));
  NOR3_X1   g666(.A1(new_n1084), .A2(new_n1085), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1073), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n1077), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1050), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1045), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1004), .B1(new_n1099), .B2(new_n988), .ZN(new_n1100));
  AND2_X1   g675(.A1(G290), .A2(G1986), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n912), .B1(new_n1101), .B2(new_n932), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n916), .A2(new_n930), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n936), .B1(new_n1100), .B2(new_n1103), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g679(.A(G319), .B1(new_n635), .B2(new_n636), .ZN(new_n1106));
  NOR3_X1   g680(.A1(G229), .A2(G227), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g681(.A1(new_n898), .A2(new_n845), .A3(new_n1107), .ZN(G225));
  INV_X1    g682(.A(G225), .ZN(G308));
endmodule


