

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U548 ( .A1(n589), .A2(n710), .ZN(n664) );
  XOR2_X1 U549 ( .A(KEYINPUT64), .B(n541), .Z(n792) );
  NOR2_X1 U550 ( .A1(G651), .A2(n570), .ZN(n786) );
  XNOR2_X2 U551 ( .A(n529), .B(n528), .ZN(G164) );
  NOR2_X2 U552 ( .A1(G2105), .A2(n522), .ZN(n878) );
  NOR2_X2 U553 ( .A1(G164), .A2(G1384), .ZN(n710) );
  INV_X1 U554 ( .A(KEYINPUT17), .ZN(n517) );
  NOR2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XNOR2_X1 U556 ( .A(n678), .B(KEYINPUT99), .ZN(n680) );
  NOR2_X1 U557 ( .A1(n536), .A2(n535), .ZN(G160) );
  AND2_X1 U558 ( .A1(n681), .A2(n679), .ZN(n514) );
  AND2_X1 U559 ( .A1(n618), .A2(n617), .ZN(n515) );
  XOR2_X1 U560 ( .A(n637), .B(KEYINPUT28), .Z(n516) );
  INV_X1 U561 ( .A(G2105), .ZN(n523) );
  INV_X1 U562 ( .A(n656), .ZN(n646) );
  AND2_X1 U563 ( .A1(n619), .A2(n515), .ZN(n620) );
  OR2_X1 U564 ( .A1(n654), .A2(n647), .ZN(n648) );
  INV_X1 U565 ( .A(KEYINPUT97), .ZN(n659) );
  XNOR2_X1 U566 ( .A(n660), .B(n659), .ZN(n673) );
  NAND2_X1 U567 ( .A1(n879), .A2(G138), .ZN(n520) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n523), .ZN(n883) );
  INV_X1 U569 ( .A(KEYINPUT40), .ZN(n748) );
  XNOR2_X2 U570 ( .A(n518), .B(n517), .ZN(n879) );
  INV_X1 U571 ( .A(G2104), .ZN(n522) );
  NAND2_X1 U572 ( .A1(G102), .A2(n878), .ZN(n519) );
  NAND2_X1 U573 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U574 ( .A(n521), .B(KEYINPUT86), .ZN(n527) );
  NOR2_X1 U575 ( .A1(n522), .A2(n523), .ZN(n882) );
  NAND2_X1 U576 ( .A1(G114), .A2(n882), .ZN(n525) );
  NAND2_X1 U577 ( .A1(G126), .A2(n883), .ZN(n524) );
  NAND2_X1 U578 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n529) );
  INV_X1 U580 ( .A(KEYINPUT87), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n879), .A2(G137), .ZN(n532) );
  NAND2_X1 U582 ( .A1(G101), .A2(n878), .ZN(n530) );
  XOR2_X1 U583 ( .A(KEYINPUT23), .B(n530), .Z(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n536) );
  NAND2_X1 U585 ( .A1(G113), .A2(n882), .ZN(n534) );
  NAND2_X1 U586 ( .A1(G125), .A2(n883), .ZN(n533) );
  NAND2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n535) );
  INV_X1 U588 ( .A(G651), .ZN(n540) );
  NOR2_X1 U589 ( .A1(G543), .A2(n540), .ZN(n537) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n537), .Z(n785) );
  NAND2_X1 U591 ( .A1(G64), .A2(n785), .ZN(n539) );
  XOR2_X1 U592 ( .A(KEYINPUT0), .B(G543), .Z(n570) );
  NAND2_X1 U593 ( .A1(G52), .A2(n786), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n546) );
  NOR2_X1 U595 ( .A1(G651), .A2(G543), .ZN(n788) );
  NAND2_X1 U596 ( .A1(G90), .A2(n788), .ZN(n543) );
  OR2_X1 U597 ( .A1(n540), .A2(n570), .ZN(n541) );
  NAND2_X1 U598 ( .A1(G77), .A2(n792), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n544), .Z(n545) );
  NOR2_X1 U601 ( .A1(n546), .A2(n545), .ZN(G171) );
  NAND2_X1 U602 ( .A1(n788), .A2(G89), .ZN(n547) );
  XNOR2_X1 U603 ( .A(n547), .B(KEYINPUT4), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G76), .A2(n792), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n550), .B(KEYINPUT5), .ZN(n555) );
  NAND2_X1 U607 ( .A1(G63), .A2(n785), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G51), .A2(n786), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U610 ( .A(KEYINPUT6), .B(n553), .Z(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U612 ( .A(n556), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U613 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U614 ( .A1(G75), .A2(n792), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n785), .A2(G62), .ZN(n557) );
  XOR2_X1 U616 ( .A(KEYINPUT83), .B(n557), .Z(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G88), .A2(n788), .ZN(n561) );
  NAND2_X1 U619 ( .A1(G50), .A2(n786), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U621 ( .A1(n563), .A2(n562), .ZN(G166) );
  INV_X1 U622 ( .A(G166), .ZN(G303) );
  NAND2_X1 U623 ( .A1(G651), .A2(G74), .ZN(n564) );
  XNOR2_X1 U624 ( .A(KEYINPUT79), .B(n564), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n786), .A2(G49), .ZN(n565) );
  XOR2_X1 U626 ( .A(KEYINPUT78), .B(n565), .Z(n566) );
  NOR2_X1 U627 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U628 ( .A(KEYINPUT80), .B(n568), .Z(n569) );
  NOR2_X1 U629 ( .A1(n785), .A2(n569), .ZN(n572) );
  NAND2_X1 U630 ( .A1(n570), .A2(G87), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(G288) );
  NAND2_X1 U632 ( .A1(G73), .A2(n792), .ZN(n574) );
  XNOR2_X1 U633 ( .A(KEYINPUT82), .B(KEYINPUT2), .ZN(n573) );
  XNOR2_X1 U634 ( .A(n574), .B(n573), .ZN(n581) );
  NAND2_X1 U635 ( .A1(G86), .A2(n788), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G48), .A2(n786), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U638 ( .A1(G61), .A2(n785), .ZN(n577) );
  XNOR2_X1 U639 ( .A(KEYINPUT81), .B(n577), .ZN(n578) );
  NOR2_X1 U640 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U641 ( .A1(n581), .A2(n580), .ZN(G305) );
  NAND2_X1 U642 ( .A1(G60), .A2(n785), .ZN(n583) );
  NAND2_X1 U643 ( .A1(G85), .A2(n788), .ZN(n582) );
  NAND2_X1 U644 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U645 ( .A1(G47), .A2(n786), .ZN(n584) );
  XNOR2_X1 U646 ( .A(KEYINPUT65), .B(n584), .ZN(n585) );
  NOR2_X1 U647 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U648 ( .A1(G72), .A2(n792), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n588), .A2(n587), .ZN(G290) );
  NAND2_X1 U650 ( .A1(G160), .A2(G40), .ZN(n711) );
  INV_X1 U651 ( .A(n711), .ZN(n589) );
  INV_X2 U652 ( .A(n664), .ZN(n641) );
  NAND2_X1 U653 ( .A1(n641), .A2(G2067), .ZN(n591) );
  NAND2_X1 U654 ( .A1(G1348), .A2(n664), .ZN(n590) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT95), .B(n592), .Z(n622) );
  NAND2_X1 U657 ( .A1(G66), .A2(n785), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G92), .A2(n788), .ZN(n593) );
  NAND2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n600) );
  NAND2_X1 U660 ( .A1(n786), .A2(G54), .ZN(n595) );
  XOR2_X1 U661 ( .A(KEYINPUT69), .B(n595), .Z(n597) );
  NAND2_X1 U662 ( .A1(G79), .A2(n792), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U664 ( .A(KEYINPUT70), .B(n598), .ZN(n599) );
  NOR2_X1 U665 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U666 ( .A(n601), .B(KEYINPUT15), .ZN(n972) );
  NAND2_X1 U667 ( .A1(n622), .A2(n972), .ZN(n621) );
  NAND2_X1 U668 ( .A1(n785), .A2(G56), .ZN(n602) );
  XNOR2_X1 U669 ( .A(n602), .B(KEYINPUT14), .ZN(n609) );
  NAND2_X1 U670 ( .A1(G68), .A2(n792), .ZN(n605) );
  NAND2_X1 U671 ( .A1(n788), .A2(G81), .ZN(n603) );
  XNOR2_X1 U672 ( .A(n603), .B(KEYINPUT12), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n607) );
  XNOR2_X1 U674 ( .A(KEYINPUT13), .B(KEYINPUT66), .ZN(n606) );
  XNOR2_X1 U675 ( .A(n607), .B(n606), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U677 ( .A(n610), .B(KEYINPUT67), .ZN(n612) );
  NAND2_X1 U678 ( .A1(G43), .A2(n786), .ZN(n611) );
  NAND2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n968) );
  XNOR2_X1 U680 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n615) );
  NOR2_X1 U681 ( .A1(G1996), .A2(n615), .ZN(n613) );
  NOR2_X1 U682 ( .A1(n968), .A2(n613), .ZN(n619) );
  INV_X1 U683 ( .A(G1341), .ZN(n967) );
  NAND2_X1 U684 ( .A1(n967), .A2(n615), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n614), .A2(n664), .ZN(n618) );
  AND2_X1 U686 ( .A1(n641), .A2(G1996), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n617) );
  NAND2_X1 U688 ( .A1(n621), .A2(n620), .ZN(n635) );
  NOR2_X1 U689 ( .A1(n622), .A2(n972), .ZN(n633) );
  NAND2_X1 U690 ( .A1(n641), .A2(G2072), .ZN(n623) );
  XNOR2_X1 U691 ( .A(n623), .B(KEYINPUT27), .ZN(n625) );
  INV_X1 U692 ( .A(G1956), .ZN(n989) );
  NOR2_X1 U693 ( .A1(n989), .A2(n641), .ZN(n624) );
  NOR2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n636) );
  NAND2_X1 U695 ( .A1(G65), .A2(n785), .ZN(n627) );
  NAND2_X1 U696 ( .A1(G91), .A2(n788), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U698 ( .A1(n786), .A2(G53), .ZN(n629) );
  NAND2_X1 U699 ( .A1(G78), .A2(n792), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n801) );
  AND2_X1 U702 ( .A1(n636), .A2(n801), .ZN(n632) );
  NOR2_X1 U703 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n638) );
  NOR2_X1 U705 ( .A1(n636), .A2(n801), .ZN(n637) );
  NAND2_X1 U706 ( .A1(n638), .A2(n516), .ZN(n640) );
  XOR2_X1 U707 ( .A(KEYINPUT96), .B(KEYINPUT29), .Z(n639) );
  XNOR2_X1 U708 ( .A(n640), .B(n639), .ZN(n645) );
  OR2_X1 U709 ( .A1(n641), .A2(G1961), .ZN(n643) );
  XNOR2_X1 U710 ( .A(G2078), .B(KEYINPUT25), .ZN(n944) );
  NAND2_X1 U711 ( .A1(n641), .A2(n944), .ZN(n642) );
  NAND2_X1 U712 ( .A1(n643), .A2(n642), .ZN(n650) );
  NAND2_X1 U713 ( .A1(n650), .A2(G171), .ZN(n644) );
  NAND2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n662) );
  NAND2_X1 U715 ( .A1(G8), .A2(n664), .ZN(n693) );
  NOR2_X1 U716 ( .A1(G1966), .A2(n693), .ZN(n654) );
  NOR2_X1 U717 ( .A1(G2084), .A2(n664), .ZN(n656) );
  NAND2_X1 U718 ( .A1(n646), .A2(G8), .ZN(n647) );
  XNOR2_X1 U719 ( .A(KEYINPUT30), .B(n648), .ZN(n649) );
  NOR2_X1 U720 ( .A1(G168), .A2(n649), .ZN(n652) );
  NOR2_X1 U721 ( .A1(G171), .A2(n650), .ZN(n651) );
  NOR2_X1 U722 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U723 ( .A(KEYINPUT31), .B(n653), .Z(n661) );
  AND2_X1 U724 ( .A1(n662), .A2(n661), .ZN(n655) );
  NOR2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U726 ( .A1(G8), .A2(n656), .ZN(n657) );
  NAND2_X1 U727 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U729 ( .A1(G286), .A2(n663), .ZN(n669) );
  NOR2_X1 U730 ( .A1(G1971), .A2(n693), .ZN(n666) );
  NOR2_X1 U731 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U733 ( .A1(n667), .A2(G303), .ZN(n668) );
  NAND2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U735 ( .A1(n670), .A2(G8), .ZN(n671) );
  XNOR2_X1 U736 ( .A(n671), .B(KEYINPUT32), .ZN(n672) );
  NAND2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U738 ( .A(n674), .B(KEYINPUT98), .ZN(n688) );
  NOR2_X1 U739 ( .A1(G1971), .A2(G303), .ZN(n675) );
  NOR2_X1 U740 ( .A1(G1976), .A2(G288), .ZN(n958) );
  NOR2_X1 U741 ( .A1(n675), .A2(n958), .ZN(n676) );
  NAND2_X1 U742 ( .A1(n688), .A2(n676), .ZN(n677) );
  NAND2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n959) );
  NAND2_X1 U744 ( .A1(n677), .A2(n959), .ZN(n678) );
  INV_X1 U745 ( .A(n693), .ZN(n681) );
  INV_X1 U746 ( .A(KEYINPUT33), .ZN(n679) );
  NAND2_X1 U747 ( .A1(n680), .A2(n514), .ZN(n684) );
  NAND2_X1 U748 ( .A1(n958), .A2(n681), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n682), .A2(KEYINPUT33), .ZN(n683) );
  NAND2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U751 ( .A(n685), .B(KEYINPUT100), .ZN(n686) );
  XOR2_X1 U752 ( .A(G1981), .B(G305), .Z(n978) );
  AND2_X1 U753 ( .A1(n686), .A2(n978), .ZN(n698) );
  NOR2_X1 U754 ( .A1(G2090), .A2(G303), .ZN(n687) );
  NAND2_X1 U755 ( .A1(G8), .A2(n687), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U757 ( .A1(n690), .A2(n693), .ZN(n696) );
  NOR2_X1 U758 ( .A1(G1981), .A2(G305), .ZN(n691) );
  XNOR2_X1 U759 ( .A(n691), .B(KEYINPUT93), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n692), .B(KEYINPUT24), .ZN(n694) );
  OR2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n732) );
  XOR2_X1 U764 ( .A(G1986), .B(G290), .Z(n970) );
  XOR2_X1 U765 ( .A(G2067), .B(KEYINPUT37), .Z(n699) );
  XNOR2_X1 U766 ( .A(KEYINPUT88), .B(n699), .ZN(n740) );
  NAND2_X1 U767 ( .A1(G116), .A2(n882), .ZN(n701) );
  NAND2_X1 U768 ( .A1(G128), .A2(n883), .ZN(n700) );
  NAND2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n702), .B(KEYINPUT35), .ZN(n707) );
  NAND2_X1 U771 ( .A1(G104), .A2(n878), .ZN(n704) );
  NAND2_X1 U772 ( .A1(G140), .A2(n879), .ZN(n703) );
  NAND2_X1 U773 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U774 ( .A(KEYINPUT34), .B(n705), .Z(n706) );
  NAND2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U776 ( .A(n708), .B(KEYINPUT36), .ZN(n892) );
  NAND2_X1 U777 ( .A1(n740), .A2(n892), .ZN(n709) );
  XOR2_X1 U778 ( .A(KEYINPUT89), .B(n709), .Z(n909) );
  NAND2_X1 U779 ( .A1(n970), .A2(n909), .ZN(n712) );
  NOR2_X1 U780 ( .A1(n710), .A2(n711), .ZN(n743) );
  NAND2_X1 U781 ( .A1(n712), .A2(n743), .ZN(n730) );
  NAND2_X1 U782 ( .A1(G95), .A2(n878), .ZN(n714) );
  NAND2_X1 U783 ( .A1(G131), .A2(n879), .ZN(n713) );
  NAND2_X1 U784 ( .A1(n714), .A2(n713), .ZN(n719) );
  NAND2_X1 U785 ( .A1(G107), .A2(n882), .ZN(n716) );
  NAND2_X1 U786 ( .A1(G119), .A2(n883), .ZN(n715) );
  NAND2_X1 U787 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U788 ( .A(KEYINPUT90), .B(n717), .ZN(n718) );
  NOR2_X1 U789 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U790 ( .A(n720), .B(KEYINPUT91), .ZN(n873) );
  XNOR2_X1 U791 ( .A(KEYINPUT92), .B(G1991), .ZN(n939) );
  NAND2_X1 U792 ( .A1(n873), .A2(n939), .ZN(n729) );
  NAND2_X1 U793 ( .A1(G141), .A2(n879), .ZN(n722) );
  NAND2_X1 U794 ( .A1(G129), .A2(n883), .ZN(n721) );
  NAND2_X1 U795 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U796 ( .A1(n878), .A2(G105), .ZN(n723) );
  XOR2_X1 U797 ( .A(KEYINPUT38), .B(n723), .Z(n724) );
  NOR2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n727) );
  NAND2_X1 U799 ( .A1(n882), .A2(G117), .ZN(n726) );
  NAND2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n874) );
  NAND2_X1 U801 ( .A1(G1996), .A2(n874), .ZN(n728) );
  NAND2_X1 U802 ( .A1(n729), .A2(n728), .ZN(n927) );
  NAND2_X1 U803 ( .A1(n743), .A2(n927), .ZN(n733) );
  NAND2_X1 U804 ( .A1(n730), .A2(n733), .ZN(n731) );
  NOR2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n747) );
  NOR2_X1 U806 ( .A1(G1996), .A2(n874), .ZN(n920) );
  INV_X1 U807 ( .A(n733), .ZN(n736) );
  NOR2_X1 U808 ( .A1(G1986), .A2(G290), .ZN(n734) );
  NOR2_X1 U809 ( .A1(n939), .A2(n873), .ZN(n923) );
  NOR2_X1 U810 ( .A1(n734), .A2(n923), .ZN(n735) );
  NOR2_X1 U811 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U812 ( .A1(n920), .A2(n737), .ZN(n738) );
  XNOR2_X1 U813 ( .A(KEYINPUT39), .B(n738), .ZN(n739) );
  NAND2_X1 U814 ( .A1(n909), .A2(n739), .ZN(n742) );
  NOR2_X1 U815 ( .A1(n740), .A2(n892), .ZN(n741) );
  XNOR2_X1 U816 ( .A(n741), .B(KEYINPUT101), .ZN(n908) );
  NAND2_X1 U817 ( .A1(n742), .A2(n908), .ZN(n744) );
  NAND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U819 ( .A(KEYINPUT102), .B(n745), .Z(n746) );
  NOR2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n749) );
  XNOR2_X1 U821 ( .A(n749), .B(n748), .ZN(G329) );
  XOR2_X1 U822 ( .A(G2430), .B(G2443), .Z(n751) );
  XNOR2_X1 U823 ( .A(KEYINPUT103), .B(G2451), .ZN(n750) );
  XNOR2_X1 U824 ( .A(n751), .B(n750), .ZN(n758) );
  XOR2_X1 U825 ( .A(G2435), .B(G2427), .Z(n753) );
  XNOR2_X1 U826 ( .A(G2446), .B(G2454), .ZN(n752) );
  XNOR2_X1 U827 ( .A(n753), .B(n752), .ZN(n754) );
  XOR2_X1 U828 ( .A(n754), .B(G2438), .Z(n756) );
  XNOR2_X1 U829 ( .A(G1348), .B(G1341), .ZN(n755) );
  XNOR2_X1 U830 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U831 ( .A(n758), .B(n757), .ZN(n759) );
  AND2_X1 U832 ( .A1(n759), .A2(G14), .ZN(G401) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U834 ( .A(G57), .ZN(G237) );
  INV_X1 U835 ( .A(G132), .ZN(G219) );
  INV_X1 U836 ( .A(G82), .ZN(G220) );
  INV_X1 U837 ( .A(n801), .ZN(G299) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n760) );
  XNOR2_X1 U839 ( .A(n760), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U840 ( .A(G223), .ZN(n823) );
  NAND2_X1 U841 ( .A1(n823), .A2(G567), .ZN(n761) );
  XOR2_X1 U842 ( .A(KEYINPUT11), .B(n761), .Z(G234) );
  INV_X1 U843 ( .A(G860), .ZN(n830) );
  OR2_X1 U844 ( .A1(n968), .A2(n830), .ZN(G153) );
  INV_X1 U845 ( .A(G171), .ZN(G301) );
  NAND2_X1 U846 ( .A1(G301), .A2(G868), .ZN(n762) );
  XNOR2_X1 U847 ( .A(n762), .B(KEYINPUT68), .ZN(n764) );
  INV_X1 U848 ( .A(G868), .ZN(n808) );
  NAND2_X1 U849 ( .A1(n808), .A2(n972), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n764), .A2(n763), .ZN(G284) );
  NOR2_X1 U851 ( .A1(G286), .A2(n808), .ZN(n766) );
  NOR2_X1 U852 ( .A1(G868), .A2(G299), .ZN(n765) );
  NOR2_X1 U853 ( .A1(n766), .A2(n765), .ZN(G297) );
  NAND2_X1 U854 ( .A1(n830), .A2(G559), .ZN(n767) );
  INV_X1 U855 ( .A(n972), .ZN(n896) );
  NAND2_X1 U856 ( .A1(n767), .A2(n896), .ZN(n768) );
  XNOR2_X1 U857 ( .A(n768), .B(KEYINPUT71), .ZN(n769) );
  XOR2_X1 U858 ( .A(KEYINPUT16), .B(n769), .Z(G148) );
  NOR2_X1 U859 ( .A1(G868), .A2(n968), .ZN(n772) );
  NAND2_X1 U860 ( .A1(G868), .A2(n896), .ZN(n770) );
  NOR2_X1 U861 ( .A1(G559), .A2(n770), .ZN(n771) );
  NOR2_X1 U862 ( .A1(n772), .A2(n771), .ZN(G282) );
  NAND2_X1 U863 ( .A1(G123), .A2(n883), .ZN(n773) );
  XNOR2_X1 U864 ( .A(n773), .B(KEYINPUT18), .ZN(n774) );
  XNOR2_X1 U865 ( .A(n774), .B(KEYINPUT72), .ZN(n776) );
  NAND2_X1 U866 ( .A1(G99), .A2(n878), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G135), .A2(n879), .ZN(n778) );
  NAND2_X1 U869 ( .A1(G111), .A2(n882), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n918) );
  XNOR2_X1 U872 ( .A(n918), .B(G2096), .ZN(n782) );
  INV_X1 U873 ( .A(G2100), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(G156) );
  XNOR2_X1 U875 ( .A(n968), .B(KEYINPUT73), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n896), .A2(G559), .ZN(n783) );
  XNOR2_X1 U877 ( .A(n784), .B(n783), .ZN(n829) );
  NAND2_X1 U878 ( .A1(G67), .A2(n785), .ZN(n797) );
  NAND2_X1 U879 ( .A1(G55), .A2(n786), .ZN(n787) );
  XNOR2_X1 U880 ( .A(n787), .B(KEYINPUT76), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G93), .A2(n788), .ZN(n789) );
  XNOR2_X1 U882 ( .A(n789), .B(KEYINPUT74), .ZN(n790) );
  NAND2_X1 U883 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U884 ( .A1(G80), .A2(n792), .ZN(n793) );
  XNOR2_X1 U885 ( .A(KEYINPUT75), .B(n793), .ZN(n794) );
  NOR2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U888 ( .A(n798), .B(KEYINPUT77), .Z(n831) );
  XOR2_X1 U889 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n799) );
  XNOR2_X1 U890 ( .A(G305), .B(n799), .ZN(n800) );
  XNOR2_X1 U891 ( .A(G290), .B(n800), .ZN(n803) );
  XNOR2_X1 U892 ( .A(G166), .B(n801), .ZN(n802) );
  XNOR2_X1 U893 ( .A(n803), .B(n802), .ZN(n804) );
  XOR2_X1 U894 ( .A(n831), .B(n804), .Z(n805) );
  XNOR2_X1 U895 ( .A(n805), .B(G288), .ZN(n899) );
  XNOR2_X1 U896 ( .A(n829), .B(n899), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n806), .A2(G868), .ZN(n807) );
  XOR2_X1 U898 ( .A(KEYINPUT85), .B(n807), .Z(n810) );
  NAND2_X1 U899 ( .A1(n831), .A2(n808), .ZN(n809) );
  NAND2_X1 U900 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n811) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n811), .Z(n812) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n812), .ZN(n813) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n813), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n814), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U907 ( .A1(G220), .A2(G219), .ZN(n815) );
  XOR2_X1 U908 ( .A(KEYINPUT22), .B(n815), .Z(n816) );
  NOR2_X1 U909 ( .A1(G218), .A2(n816), .ZN(n817) );
  NAND2_X1 U910 ( .A1(G96), .A2(n817), .ZN(n827) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n827), .ZN(n821) );
  NAND2_X1 U912 ( .A1(G69), .A2(G120), .ZN(n818) );
  NOR2_X1 U913 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U914 ( .A1(G108), .A2(n819), .ZN(n828) );
  NAND2_X1 U915 ( .A1(G567), .A2(n828), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n833) );
  NAND2_X1 U917 ( .A1(G483), .A2(G661), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n833), .A2(n822), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U922 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U924 ( .A1(n826), .A2(n825), .ZN(G188) );
  XOR2_X1 U925 ( .A(G96), .B(KEYINPUT104), .Z(G221) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  INV_X1 U928 ( .A(G69), .ZN(G235) );
  NOR2_X1 U929 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  NAND2_X1 U931 ( .A1(n830), .A2(n829), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(G145) );
  XNOR2_X1 U933 ( .A(KEYINPUT105), .B(n833), .ZN(G319) );
  XOR2_X1 U934 ( .A(KEYINPUT43), .B(KEYINPUT42), .Z(n835) );
  XNOR2_X1 U935 ( .A(G2090), .B(KEYINPUT106), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U937 ( .A(n836), .B(G2100), .Z(n838) );
  XNOR2_X1 U938 ( .A(G2072), .B(G2067), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U940 ( .A(G2096), .B(G2678), .Z(n840) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U944 ( .A(G1981), .B(G1971), .Z(n844) );
  XNOR2_X1 U945 ( .A(G1966), .B(G1961), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U947 ( .A(G1991), .B(G1976), .Z(n846) );
  XNOR2_X1 U948 ( .A(G1956), .B(G1996), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U950 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U951 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U953 ( .A(G1986), .B(G2474), .Z(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U955 ( .A1(G124), .A2(n883), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n853), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U957 ( .A1(G100), .A2(n878), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n854), .B(KEYINPUT108), .ZN(n855) );
  NAND2_X1 U959 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G136), .A2(n879), .ZN(n858) );
  NAND2_X1 U961 ( .A1(G112), .A2(n882), .ZN(n857) );
  NAND2_X1 U962 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U963 ( .A1(n860), .A2(n859), .ZN(G162) );
  NAND2_X1 U964 ( .A1(G118), .A2(n882), .ZN(n862) );
  NAND2_X1 U965 ( .A1(G130), .A2(n883), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G106), .A2(n878), .ZN(n864) );
  NAND2_X1 U968 ( .A1(G142), .A2(n879), .ZN(n863) );
  NAND2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U970 ( .A(KEYINPUT45), .B(n865), .Z(n866) );
  NOR2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U972 ( .A(n918), .B(n868), .ZN(n872) );
  XOR2_X1 U973 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n870) );
  XNOR2_X1 U974 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n869) );
  XNOR2_X1 U975 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U976 ( .A(n872), .B(n871), .ZN(n877) );
  XNOR2_X1 U977 ( .A(G160), .B(n873), .ZN(n875) );
  XNOR2_X1 U978 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U979 ( .A(n877), .B(n876), .Z(n891) );
  NAND2_X1 U980 ( .A1(G103), .A2(n878), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G139), .A2(n879), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n889) );
  NAND2_X1 U983 ( .A1(G115), .A2(n882), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G127), .A2(n883), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U986 ( .A(KEYINPUT109), .B(n886), .ZN(n887) );
  XNOR2_X1 U987 ( .A(KEYINPUT47), .B(n887), .ZN(n888) );
  NOR2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n910) );
  XNOR2_X1 U989 ( .A(n910), .B(G162), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n892), .B(G164), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U993 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U994 ( .A(n968), .B(G286), .ZN(n898) );
  XNOR2_X1 U995 ( .A(G171), .B(n896), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U998 ( .A1(G37), .A2(n901), .ZN(G397) );
  NOR2_X1 U999 ( .A1(G227), .A2(G229), .ZN(n902) );
  XOR2_X1 U1000 ( .A(KEYINPUT49), .B(n902), .Z(n903) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n903), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(G401), .A2(n904), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(KEYINPUT112), .B(n905), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1008 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1022) );
  INV_X1 U1009 ( .A(KEYINPUT55), .ZN(n953) );
  NAND2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(G2072), .B(n910), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(G164), .B(G2078), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1014 ( .A(KEYINPUT113), .B(n913), .Z(n914) );
  XNOR2_X1 U1015 ( .A(KEYINPUT50), .B(n914), .ZN(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n929) );
  XOR2_X1 U1017 ( .A(G2084), .B(G160), .Z(n917) );
  NOR2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n925) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(n921), .B(KEYINPUT51), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(KEYINPUT52), .B(n930), .ZN(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT114), .B(n931), .Z(n932) );
  NAND2_X1 U1028 ( .A1(n953), .A2(n932), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n933), .A2(G29), .ZN(n1020) );
  XNOR2_X1 U1030 ( .A(KEYINPUT115), .B(G2090), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(n934), .B(G35), .ZN(n951) );
  XNOR2_X1 U1032 ( .A(G2084), .B(G34), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(n935), .B(KEYINPUT54), .ZN(n949) );
  XNOR2_X1 U1034 ( .A(G2072), .B(G33), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n943) );
  XOR2_X1 U1037 ( .A(G32), .B(G1996), .Z(n938) );
  NAND2_X1 U1038 ( .A1(n938), .A2(G28), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(G25), .B(n939), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n946) );
  XOR2_X1 U1042 ( .A(G27), .B(n944), .Z(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(n947), .B(KEYINPUT53), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(n953), .B(n952), .ZN(n955) );
  INV_X1 U1048 ( .A(G29), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(G11), .A2(n956), .ZN(n1018) );
  INV_X1 U1051 ( .A(G16), .ZN(n1014) );
  XOR2_X1 U1052 ( .A(KEYINPUT56), .B(KEYINPUT116), .Z(n957) );
  XNOR2_X1 U1053 ( .A(n1014), .B(n957), .ZN(n987) );
  XNOR2_X1 U1054 ( .A(G299), .B(n989), .ZN(n965) );
  XNOR2_X1 U1055 ( .A(KEYINPUT119), .B(n958), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1057 ( .A(G1971), .B(G166), .Z(n961) );
  XNOR2_X1 U1058 ( .A(KEYINPUT120), .B(n961), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n966), .B(KEYINPUT121), .ZN(n985) );
  XNOR2_X1 U1062 ( .A(KEYINPUT122), .B(n967), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(n968), .ZN(n977) );
  XNOR2_X1 U1064 ( .A(G171), .B(G1961), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(G1348), .B(n972), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(KEYINPUT118), .B(n973), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n983) );
  XNOR2_X1 U1070 ( .A(G1966), .B(G168), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n980), .B(KEYINPUT117), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(n981), .B(KEYINPUT57), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n1016) );
  XNOR2_X1 U1077 ( .A(KEYINPUT123), .B(G1961), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(n988), .B(G5), .ZN(n1003) );
  XNOR2_X1 U1079 ( .A(n989), .B(G20), .ZN(n997) );
  XOR2_X1 U1080 ( .A(G1981), .B(G6), .Z(n992) );
  XOR2_X1 U1081 ( .A(KEYINPUT124), .B(G19), .Z(n990) );
  XNOR2_X1 U1082 ( .A(G1341), .B(n990), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n995) );
  XOR2_X1 U1084 ( .A(KEYINPUT59), .B(G1348), .Z(n993) );
  XNOR2_X1 U1085 ( .A(G4), .B(n993), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(n998), .B(KEYINPUT60), .ZN(n999) );
  XOR2_X1 U1089 ( .A(KEYINPUT125), .B(n999), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G21), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1011) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(G24), .B(G1986), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1008) );
  XOR2_X1 U1096 ( .A(G1976), .B(KEYINPUT126), .Z(n1006) );
  XNOR2_X1 U1097 ( .A(G23), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT58), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(KEYINPUT61), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1022), .B(n1021), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

