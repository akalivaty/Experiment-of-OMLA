//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1214, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1286, new_n1287,
    new_n1288;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AND2_X1   g0006(.A1(G68), .A2(G238), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n207), .B(new_n212), .C1(G107), .C2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G116), .A2(G270), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n203), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G68), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n221), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n206), .B(new_n225), .C1(new_n228), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT64), .B(G250), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G257), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NAND2_X1  g0049(.A1(G33), .A2(G97), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n222), .A2(G1698), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G226), .B2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n250), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT65), .B(G41), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n263), .B(G274), .C1(new_n264), .C2(G45), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n260), .A2(G238), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n262), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT13), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT13), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  OR3_X1    g0074(.A1(new_n273), .A2(KEYINPUT14), .A3(new_n274), .ZN(new_n275));
  OR3_X1    g0075(.A1(new_n269), .A2(KEYINPUT69), .A3(new_n271), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n269), .B1(KEYINPUT69), .B2(new_n271), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G179), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT14), .B1(new_n273), .B2(new_n274), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n227), .A2(G33), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n281), .A2(new_n218), .B1(new_n227), .B2(G68), .ZN(new_n282));
  XOR2_X1   g0082(.A(new_n282), .B(KEYINPUT70), .Z(new_n283));
  NAND2_X1  g0083(.A1(new_n227), .A2(new_n253), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n216), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT66), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT66), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n288), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n287), .A2(new_n226), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT11), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT11), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n285), .A2(new_n293), .A3(new_n290), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT12), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n296), .B1(new_n298), .B2(new_n229), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n297), .A2(KEYINPUT12), .A3(G68), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n263), .A2(G20), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n287), .A2(new_n289), .A3(new_n226), .A4(new_n301), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n299), .A2(new_n300), .B1(new_n302), .B2(new_n229), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n295), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n280), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G20), .A2(G77), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT8), .B(G58), .ZN(new_n308));
  XOR2_X1   g0108(.A(KEYINPUT15), .B(G87), .Z(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n307), .B1(new_n284), .B2(new_n308), .C1(new_n310), .C2(new_n281), .ZN(new_n311));
  INV_X1    g0111(.A(new_n302), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n311), .A2(new_n290), .B1(G77), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n298), .A2(new_n218), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT3), .B(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G238), .A2(G1698), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(new_n317), .C1(new_n222), .C2(G1698), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(new_n261), .C1(G107), .C2(new_n316), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n260), .A2(new_n266), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n319), .B(new_n265), .C1(new_n219), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n274), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n315), .B(new_n322), .C1(G179), .C2(new_n321), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n306), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n308), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n302), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT72), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n308), .A2(new_n297), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n326), .B2(new_n328), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n290), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT7), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n316), .B2(G20), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT71), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G58), .A2(G68), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n227), .B1(new_n230), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G159), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n284), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n337), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(G58), .A2(G68), .ZN(new_n343));
  NOR2_X1   g0143(.A1(G58), .A2(G68), .ZN(new_n344));
  OAI21_X1  g0144(.A(G20), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(KEYINPUT71), .C1(new_n340), .C2(new_n284), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n336), .A2(G68), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n332), .B1(new_n347), .B2(KEYINPUT16), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n229), .B1(new_n334), .B2(new_n335), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n345), .B1(new_n340), .B2(new_n284), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n331), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G1698), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n254), .A2(new_n256), .A3(G223), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT73), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT73), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n316), .A2(new_n357), .A3(G223), .A4(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G87), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n316), .A2(G226), .A3(G1698), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n356), .A2(new_n358), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n261), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT74), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n260), .A2(G232), .A3(new_n266), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n265), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n363), .B1(new_n265), .B2(new_n364), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n362), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n265), .A2(new_n364), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(new_n361), .B2(new_n261), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n368), .A2(G190), .B1(G200), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n353), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT17), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n353), .A2(new_n371), .A3(KEYINPUT17), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n370), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n369), .A2(KEYINPUT74), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(new_n365), .B1(new_n261), .B2(new_n361), .ZN(new_n379));
  INV_X1    g0179(.A(G179), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n274), .A2(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n316), .A2(new_n333), .A3(G20), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT7), .B1(new_n257), .B2(new_n227), .ZN(new_n383));
  OAI21_X1  g0183(.A(G68), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n342), .A2(new_n346), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT16), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(new_n352), .A3(new_n290), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n329), .A2(new_n330), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n381), .A2(KEYINPUT18), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT18), .B1(new_n381), .B2(new_n389), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n324), .A2(new_n376), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n276), .A2(G190), .A3(new_n277), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n270), .A2(G200), .A3(new_n272), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n394), .A2(new_n295), .A3(new_n304), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n227), .B1(new_n344), .B2(new_n216), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT67), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G150), .ZN(new_n401));
  OAI221_X1 g0201(.A(new_n400), .B1(new_n401), .B2(new_n284), .C1(new_n308), .C2(new_n281), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(new_n290), .B1(G50), .B2(new_n312), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n298), .A2(new_n216), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT68), .A3(KEYINPUT9), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT68), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT9), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n407), .A2(new_n408), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n403), .A2(new_n404), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n406), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n354), .A2(G222), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G223), .A2(G1698), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n316), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(new_n261), .C1(G77), .C2(new_n316), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(new_n265), .C1(new_n217), .C2(new_n320), .ZN(new_n418));
  INV_X1    g0218(.A(G190), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(G200), .B2(new_n418), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT10), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT10), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n413), .A2(new_n424), .A3(new_n421), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n418), .A2(new_n274), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n405), .B(new_n427), .C1(G179), .C2(new_n418), .ZN(new_n428));
  INV_X1    g0228(.A(new_n315), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n321), .A2(G200), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(new_n430), .C1(new_n419), .C2(new_n321), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n397), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G41), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT65), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT65), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G41), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT5), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(KEYINPUT5), .ZN(new_n440));
  INV_X1    g0240(.A(G45), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(G1), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(G264), .A3(new_n260), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n209), .A2(new_n354), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n211), .A2(G1698), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n254), .A3(new_n256), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G294), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n261), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n440), .A2(KEYINPUT75), .ZN(new_n451));
  INV_X1    g0251(.A(G274), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n440), .B2(KEYINPUT75), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n451), .A2(new_n453), .A3(new_n439), .A4(new_n442), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n444), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT82), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n444), .A2(new_n450), .A3(KEYINPUT82), .A4(new_n454), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n419), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G200), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT80), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n254), .A2(new_n256), .A3(new_n227), .A4(G87), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT22), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT22), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n316), .A2(new_n466), .A3(new_n227), .A4(G87), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT79), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n227), .A2(G107), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(KEYINPUT78), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT23), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n470), .B2(new_n469), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n469), .B(new_n472), .C1(new_n470), .C2(KEYINPUT78), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G116), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT77), .B1(new_n476), .B2(G20), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT77), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n478), .A2(new_n227), .A3(G33), .A4(G116), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n474), .A2(new_n475), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n463), .B1(new_n468), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n465), .A2(new_n467), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n471), .A2(new_n473), .B1(new_n477), .B2(new_n479), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT80), .A4(new_n475), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n482), .A2(KEYINPUT24), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT24), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n463), .B(new_n487), .C1(new_n468), .C2(new_n481), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n290), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n253), .A2(G1), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n298), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n332), .A2(G107), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT25), .B1(new_n297), .B2(G107), .ZN(new_n493));
  OR3_X1    g0293(.A1(new_n297), .A2(KEYINPUT25), .A3(G107), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n495), .B(KEYINPUT81), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n462), .A2(new_n489), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n457), .A2(new_n458), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G169), .ZN(new_n499));
  INV_X1    g0299(.A(new_n455), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G179), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n496), .A2(new_n489), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n254), .A2(new_n256), .A3(G244), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G283), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n505), .A2(G1698), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n508), .A2(new_n254), .A3(new_n256), .A4(G244), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n254), .A2(new_n256), .A3(G250), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n354), .B1(new_n511), .B2(KEYINPUT4), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n261), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n443), .A2(G257), .A3(new_n260), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n454), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G200), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n513), .A2(G190), .A3(new_n454), .A4(new_n514), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n297), .A2(G97), .ZN(new_n518));
  OAI21_X1  g0318(.A(G107), .B1(new_n382), .B2(new_n383), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n284), .A2(new_n218), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT6), .ZN(new_n521));
  AND2_X1   g0321(.A1(G97), .A2(G107), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G97), .A2(G107), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G107), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(KEYINPUT6), .A3(G97), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n520), .B1(new_n527), .B2(G20), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n519), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n518), .B1(new_n529), .B2(new_n290), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n332), .A2(G97), .A3(new_n491), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n516), .A2(new_n517), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n515), .A2(new_n274), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n524), .A2(new_n526), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n534), .A2(new_n227), .B1(new_n218), .B2(new_n284), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n525), .B1(new_n334), .B2(new_n335), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n290), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n518), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n531), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n513), .A2(new_n380), .A3(new_n454), .A4(new_n514), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n533), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n442), .A2(new_n452), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n209), .B1(new_n441), .B2(G1), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n260), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(G238), .A2(G1698), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n219), .B2(G1698), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(new_n316), .B1(G33), .B2(G116), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n544), .B1(new_n547), .B2(new_n260), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G200), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n523), .A2(new_n208), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n250), .A2(new_n227), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n550), .A2(KEYINPUT19), .A3(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n254), .A2(new_n256), .A3(new_n227), .A4(G68), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT19), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n250), .B2(G20), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n290), .B1(new_n298), .B2(new_n310), .ZN(new_n557));
  OAI211_X1 g0357(.A(G190), .B(new_n544), .C1(new_n547), .C2(new_n260), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n332), .A2(G87), .A3(new_n491), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n549), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n548), .A2(new_n274), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(new_n290), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n332), .A2(new_n491), .A3(new_n309), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n310), .A2(new_n298), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n380), .B(new_n544), .C1(new_n547), .C2(new_n260), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n561), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n532), .A2(new_n541), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n443), .A2(G270), .A3(new_n260), .ZN(new_n570));
  INV_X1    g0370(.A(G303), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n255), .A2(G33), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n354), .A2(G257), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G264), .A2(G1698), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n254), .A2(new_n256), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  AND4_X1   g0377(.A1(KEYINPUT76), .A2(new_n574), .A3(new_n261), .A4(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n260), .B1(new_n257), .B2(new_n571), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT76), .B1(new_n579), .B2(new_n577), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n454), .B(new_n570), .C1(new_n578), .C2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(G116), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G20), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n507), .B(new_n227), .C1(G33), .C2(new_n210), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n290), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT20), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n332), .A2(G116), .A3(new_n491), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT20), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n290), .A2(new_n588), .A3(new_n583), .A4(new_n584), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n298), .A2(new_n582), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n586), .A2(new_n587), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n581), .A2(G169), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n578), .A2(new_n580), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n570), .A2(new_n454), .ZN(new_n596));
  OAI21_X1  g0396(.A(G200), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n591), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n570), .A2(new_n454), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT76), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n261), .B1(new_n316), .B2(G303), .ZN(new_n601));
  INV_X1    g0401(.A(new_n577), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n579), .A2(KEYINPUT76), .A3(new_n577), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n599), .A2(G190), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n597), .A2(new_n598), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n581), .A2(new_n591), .A3(KEYINPUT21), .A4(G169), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n591), .A2(new_n599), .A3(G179), .A4(new_n605), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n594), .A2(new_n607), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n569), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n433), .A2(new_n503), .A3(new_n611), .ZN(G372));
  INV_X1    g0412(.A(new_n376), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n324), .A2(new_n613), .A3(new_n396), .ZN(new_n614));
  INV_X1    g0414(.A(new_n392), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n426), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n428), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n433), .ZN(new_n620));
  INV_X1    g0420(.A(new_n541), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n621), .A2(KEYINPUT26), .A3(new_n560), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n489), .A2(new_n496), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n499), .A2(new_n501), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n594), .A2(new_n608), .A3(new_n609), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n489), .A2(new_n496), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n625), .A2(new_n626), .B1(new_n627), .B2(new_n462), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n560), .B(new_n532), .C1(new_n628), .C2(new_n621), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n622), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n567), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n619), .B1(new_n620), .B2(new_n633), .ZN(G369));
  XOR2_X1   g0434(.A(new_n610), .B(KEYINPUT83), .Z(new_n635));
  INV_X1    g0435(.A(G13), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(G20), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n263), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G343), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n591), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n635), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n594), .A2(new_n608), .A3(new_n609), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(new_n645), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(G330), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n503), .B1(new_n627), .B2(new_n643), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n625), .B2(new_n643), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g0454(.A(new_n643), .B(KEYINPUT84), .Z(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n502), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n647), .A2(new_n643), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n503), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n654), .A2(new_n657), .A3(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n204), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n264), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n523), .A2(new_n208), .A3(new_n582), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n663), .A2(new_n263), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n665), .B1(new_n232), .B2(new_n663), .ZN(new_n666));
  XOR2_X1   g0466(.A(new_n666), .B(KEYINPUT28), .Z(new_n667));
  INV_X1    g0467(.A(KEYINPUT89), .ZN(new_n668));
  OR3_X1    g0468(.A1(new_n633), .A2(KEYINPUT29), .A3(new_n655), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT29), .B1(new_n633), .B2(new_n644), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n515), .A2(new_n380), .A3(new_n581), .A4(new_n548), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n500), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n581), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT85), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n444), .A2(new_n450), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n548), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n675), .B(G179), .C1(new_n676), .C2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n544), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n546), .A2(new_n316), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n476), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n680), .B1(new_n682), .B2(new_n261), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n676), .A3(new_n450), .A4(new_n444), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n454), .A3(new_n514), .A4(new_n513), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n679), .A2(new_n685), .A3(KEYINPUT30), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n599), .A2(G179), .A3(new_n605), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n683), .A2(new_n450), .A3(new_n444), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n688), .B1(KEYINPUT85), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n515), .B1(new_n676), .B2(new_n678), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n674), .B1(new_n686), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT86), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n693), .A2(KEYINPUT86), .A3(KEYINPUT31), .A4(new_n655), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT87), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n532), .A2(new_n541), .A3(new_n568), .ZN(new_n700));
  INV_X1    g0500(.A(new_n610), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n462), .A2(new_n489), .A3(new_n496), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n625), .A2(new_n703), .A3(new_n656), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n699), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n503), .A2(KEYINPUT87), .A3(new_n611), .A4(new_n656), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT31), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT30), .B1(new_n679), .B2(new_n685), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n690), .A2(new_n687), .A3(new_n691), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n673), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n707), .B1(new_n710), .B2(new_n643), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n705), .A2(new_n706), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(G330), .B1(new_n698), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT88), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT88), .ZN(new_n715));
  OAI211_X1 g0515(.A(new_n715), .B(G330), .C1(new_n698), .C2(new_n712), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n668), .B1(new_n671), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n717), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(KEYINPUT89), .A3(new_n670), .A4(new_n669), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n667), .B1(new_n721), .B2(G1), .ZN(G364));
  AOI21_X1  g0522(.A(new_n226), .B1(G20), .B2(new_n274), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n227), .A2(G179), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G190), .A2(G200), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n726), .A2(KEYINPUT32), .A3(new_n340), .ZN(new_n727));
  INV_X1    g0527(.A(new_n724), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n728), .A2(G190), .A3(new_n460), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n525), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n728), .A2(new_n419), .A3(new_n460), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n257), .B(new_n731), .C1(G87), .C2(new_n732), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT92), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT32), .B1(new_n726), .B2(new_n340), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n227), .A2(new_n380), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(G190), .A3(G200), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n216), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n460), .A2(G190), .ZN(new_n739));
  OAI21_X1  g0539(.A(G20), .B1(new_n739), .B2(G179), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(new_n725), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n741), .A2(new_n210), .B1(new_n218), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n736), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n745), .A2(G190), .A3(new_n460), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n734), .B(new_n744), .C1(new_n229), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n745), .A2(new_n739), .ZN(new_n749));
  AOI211_X1 g0549(.A(new_n727), .B(new_n748), .C1(G58), .C2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G311), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n742), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n730), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G283), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n732), .B(KEYINPUT93), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G303), .ZN(new_n757));
  INV_X1    g0557(.A(G326), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n737), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(KEYINPUT33), .B(G317), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n316), .B(new_n759), .C1(new_n746), .C2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n726), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n749), .A2(G322), .B1(new_n762), .B2(G329), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n754), .A2(new_n757), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n752), .B(new_n764), .C1(G294), .C2(new_n740), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n723), .B1(new_n750), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT90), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n245), .A2(G45), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n662), .A2(new_n316), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n441), .B2(new_n232), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n771), .A2(new_n774), .B1(new_n582), .B2(new_n662), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n316), .A2(G355), .A3(new_n204), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n723), .B(new_n770), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n663), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n637), .A2(G45), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n778), .A2(G1), .A3(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n777), .B(new_n780), .C1(new_n649), .C2(new_n770), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n766), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n780), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n651), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n649), .A2(new_n650), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  NOR2_X1   g0588(.A1(new_n323), .A2(new_n644), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n431), .B1(new_n429), .B2(new_n643), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(new_n790), .B2(new_n323), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n656), .B(new_n791), .C1(new_n631), .C2(new_n632), .ZN(new_n792));
  INV_X1    g0592(.A(new_n791), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n633), .B2(new_n655), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n792), .B(new_n794), .C1(new_n717), .C2(KEYINPUT95), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n717), .A2(KEYINPUT95), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n795), .B(new_n796), .Z(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n780), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n793), .A2(new_n768), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n723), .A2(new_n767), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n218), .ZN(new_n801));
  INV_X1    g0601(.A(G283), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n747), .A2(new_n802), .B1(new_n737), .B2(new_n571), .ZN(new_n803));
  INV_X1    g0603(.A(new_n742), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(G116), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT94), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n762), .A2(G311), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n749), .A2(G294), .B1(G97), .B2(new_n740), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n316), .B1(new_n753), .B2(G87), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n806), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n755), .A2(new_n525), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n746), .A2(G150), .B1(new_n749), .B2(G143), .ZN(new_n812));
  INV_X1    g0612(.A(G137), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n813), .B2(new_n737), .C1(new_n340), .C2(new_n742), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT34), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n814), .A2(new_n815), .B1(G132), .B2(new_n762), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n753), .A2(G68), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n756), .A2(G50), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n316), .B1(new_n741), .B2(new_n221), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n810), .A2(new_n811), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n723), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n799), .A2(new_n783), .A3(new_n801), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n798), .A2(new_n824), .ZN(G384));
  NAND3_X1  g0625(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n644), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n705), .A2(new_n706), .A3(new_n711), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n433), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n829));
  XNOR2_X1  g0629(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT37), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n641), .B1(new_n387), .B2(new_n388), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n371), .B2(new_n353), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n379), .A2(new_n380), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n377), .A2(new_n274), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n389), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n831), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n389), .A2(new_n642), .ZN(new_n838));
  AND4_X1   g0638(.A1(new_n831), .A2(new_n372), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT98), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n832), .B1(new_n392), .B2(new_n376), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n372), .A2(new_n836), .A3(new_n838), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT37), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n833), .A2(new_n831), .A3(new_n836), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT98), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n840), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n326), .A2(new_n328), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n386), .A2(new_n290), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n347), .A2(KEYINPUT16), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n642), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n392), .B2(new_n376), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n381), .A2(new_n853), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n372), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n855), .B1(new_n858), .B2(KEYINPUT97), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT97), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n857), .A2(new_n372), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n831), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(KEYINPUT38), .B(new_n856), .C1(new_n862), .C2(new_n839), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n849), .A2(new_n863), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n280), .A2(new_n305), .A3(new_n643), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n305), .A2(new_n644), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n305), .A2(new_n280), .B1(new_n866), .B2(new_n396), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n827), .A2(new_n791), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT40), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT99), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  OR2_X1    g0672(.A1(KEYINPUT99), .A2(KEYINPUT40), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n827), .A2(new_n791), .A3(new_n868), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n858), .A2(KEYINPUT97), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n861), .A3(new_n854), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n839), .B1(new_n876), .B2(KEYINPUT37), .ZN(new_n877));
  INV_X1    g0677(.A(new_n856), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n848), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n863), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n872), .A2(new_n874), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n870), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n830), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(G330), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n620), .B1(new_n669), .B2(new_n670), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(new_n618), .ZN(new_n886));
  INV_X1    g0686(.A(new_n789), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n792), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(new_n868), .A3(new_n880), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n849), .A2(new_n863), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n879), .A2(KEYINPUT39), .A3(new_n863), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n865), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n392), .A2(new_n641), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n889), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n886), .B(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n884), .B(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n263), .B2(new_n637), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n527), .B(KEYINPUT96), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n582), .B1(new_n900), .B2(KEYINPUT35), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n228), .C1(KEYINPUT35), .C2(new_n900), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT36), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n338), .A2(G77), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n231), .A2(new_n904), .B1(G50), .B2(new_n229), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(G1), .A3(new_n636), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n899), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT102), .Z(G367));
  NAND3_X1  g0708(.A1(new_n756), .A2(KEYINPUT46), .A3(G116), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT105), .Z(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT46), .B1(new_n732), .B2(G116), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT106), .ZN(new_n912));
  INV_X1    g0712(.A(G317), .ZN(new_n913));
  INV_X1    g0713(.A(G294), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n257), .B1(new_n726), .B2(new_n913), .C1(new_n747), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(G283), .B2(new_n804), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n729), .A2(G97), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n910), .A2(new_n912), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n737), .A2(new_n751), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n741), .A2(new_n525), .ZN(new_n920));
  INV_X1    g0720(.A(new_n749), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n571), .ZN(new_n922));
  NOR4_X1   g0722(.A1(new_n918), .A2(new_n919), .A3(new_n920), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n749), .A2(G150), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n732), .A2(G58), .B1(new_n740), .B2(G68), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n813), .B2(new_n726), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n746), .A2(G159), .B1(G50), .B2(new_n804), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT107), .ZN(new_n928));
  INV_X1    g0728(.A(G143), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n928), .B(new_n316), .C1(new_n929), .C2(new_n737), .ZN(new_n930));
  AOI211_X1 g0730(.A(new_n926), .B(new_n930), .C1(G77), .C2(new_n729), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n923), .B1(new_n924), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT47), .Z(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n723), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n557), .A2(new_n559), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n644), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n568), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n567), .B2(new_n936), .ZN(new_n938));
  INV_X1    g0738(.A(new_n770), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n770), .A2(new_n723), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n941), .B1(new_n204), .B2(new_n310), .C1(new_n241), .C2(new_n773), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n934), .A2(new_n783), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n779), .A2(G1), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n660), .A2(new_n657), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n655), .A2(new_n539), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n532), .A3(new_n541), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n621), .A2(new_n655), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT44), .Z(new_n953));
  NAND3_X1  g0753(.A1(new_n651), .A2(KEYINPUT104), .A3(new_n653), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n947), .A2(new_n951), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT45), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT104), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n654), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n957), .B(new_n959), .Z(new_n960));
  OAI21_X1  g0760(.A(new_n660), .B1(new_n653), .B2(new_n659), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n651), .B(new_n961), .Z(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n960), .A2(new_n963), .B1(new_n718), .B2(new_n720), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n663), .B(KEYINPUT41), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n946), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n654), .A2(new_n951), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n951), .A2(new_n660), .ZN(new_n970));
  XOR2_X1   g0770(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n541), .B1(new_n949), .B2(new_n625), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n973), .A2(new_n656), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n969), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n968), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n968), .A2(new_n975), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n944), .B1(new_n967), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(G387));
  NOR2_X1   g0782(.A1(new_n310), .A2(new_n741), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n316), .B1(new_n401), .B2(new_n726), .C1(new_n730), .C2(new_n210), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(G50), .C2(new_n749), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n804), .A2(G68), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n737), .A2(new_n340), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT109), .Z(new_n988));
  AOI22_X1  g0788(.A1(new_n325), .A2(new_n746), .B1(new_n732), .B2(G77), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n985), .A2(new_n986), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n746), .A2(G311), .B1(new_n749), .B2(G317), .ZN(new_n991));
  INV_X1    g0791(.A(G322), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n991), .B1(new_n571), .B2(new_n742), .C1(new_n992), .C2(new_n737), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT48), .ZN(new_n994));
  INV_X1    g0794(.A(new_n732), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n994), .B1(new_n802), .B2(new_n741), .C1(new_n914), .C2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT49), .Z(new_n997));
  INV_X1    g0797(.A(new_n729), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n257), .B1(new_n758), .B2(new_n726), .C1(new_n998), .C2(new_n582), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n990), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n723), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n653), .B2(new_n939), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n308), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n664), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(G68), .A2(G77), .ZN(new_n1005));
  OAI21_X1  g0805(.A(KEYINPUT50), .B1(new_n308), .B2(G50), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1004), .A2(new_n441), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n772), .B(new_n1007), .C1(new_n237), .C2(new_n441), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n316), .A2(new_n664), .A3(new_n204), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(G107), .B2(new_n204), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT108), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1002), .B1(new_n941), .B2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n945), .A2(new_n963), .B1(new_n1013), .B2(new_n783), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n718), .A2(new_n720), .A3(new_n962), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n663), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n962), .B1(new_n718), .B2(new_n720), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(G393));
  NOR2_X1   g0818(.A1(new_n995), .A2(new_n229), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n741), .A2(new_n218), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G50), .B2(new_n746), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n308), .B2(new_n742), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT110), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n921), .A2(new_n340), .B1(new_n401), .B2(new_n737), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT51), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n753), .A2(G87), .B1(G143), .B2(new_n762), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1023), .A2(new_n1025), .A3(new_n316), .A4(new_n1026), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1019), .B(new_n1027), .C1(KEYINPUT110), .C2(new_n1022), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n316), .B(new_n731), .C1(G322), .C2(new_n762), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n740), .A2(G116), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n921), .A2(new_n751), .B1(new_n913), .B2(new_n737), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT52), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n746), .A2(G303), .B1(G294), .B2(new_n804), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G283), .B2(new_n732), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n723), .B1(new_n1028), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n951), .A2(new_n770), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n941), .B1(new_n210), .B2(new_n204), .C1(new_n248), .C2(new_n773), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1036), .A2(new_n783), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n960), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n721), .A2(new_n963), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(new_n1040), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n663), .B1(new_n1017), .B2(new_n960), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1039), .B1(new_n946), .B2(new_n1040), .C1(new_n1042), .C2(new_n1043), .ZN(G390));
  NOR2_X1   g0844(.A1(new_n869), .A2(new_n650), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n793), .B1(new_n714), .B2(new_n716), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1046), .B1(new_n1047), .B2(new_n868), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n827), .A2(new_n791), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n868), .B1(new_n1049), .B2(G330), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1047), .B2(new_n868), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n790), .A2(new_n323), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n643), .B(new_n1052), .C1(new_n631), .C2(new_n632), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n887), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n888), .A2(new_n1048), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n828), .A2(new_n650), .ZN(new_n1057));
  OR3_X1    g0857(.A1(new_n885), .A2(new_n618), .A3(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n865), .B(KEYINPUT111), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n868), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n890), .B(new_n1060), .C1(new_n1055), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n892), .A2(new_n893), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n792), .B2(new_n887), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n865), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1047), .A2(new_n868), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n1062), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1046), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1056), .A2(new_n1058), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1048), .A2(new_n888), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1050), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1066), .A2(new_n1055), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1065), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n864), .B(new_n1059), .C1(new_n1054), .C2(new_n868), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1045), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1062), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n885), .A2(new_n1057), .A3(new_n618), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1073), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1069), .A2(new_n663), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1063), .A2(new_n768), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n800), .A2(new_n308), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n732), .A2(G150), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT113), .Z(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT53), .ZN(new_n1085));
  INV_X1    g0885(.A(G125), .ZN(new_n1086));
  XOR2_X1   g0886(.A(KEYINPUT54), .B(G143), .Z(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n316), .B1(new_n1086), .B2(new_n726), .C1(new_n1088), .C2(new_n742), .ZN(new_n1089));
  INV_X1    g0889(.A(G132), .ZN(new_n1090));
  INV_X1    g0890(.A(G128), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n921), .A2(new_n1090), .B1(new_n1091), .B2(new_n737), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT112), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1089), .B(new_n1093), .C1(G159), .C2(new_n740), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n813), .B2(new_n747), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1085), .B(new_n1095), .C1(G50), .C2(new_n729), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n726), .A2(new_n914), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n316), .B1(new_n756), .B2(G87), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n804), .A2(G97), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n737), .A2(new_n802), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1100), .B(new_n1020), .C1(G116), .C2(new_n749), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1098), .A2(new_n818), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1097), .B(new_n1102), .C1(G107), .C2(new_n746), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n723), .B1(new_n1096), .B2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1081), .A2(new_n783), .A3(new_n1082), .A4(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT114), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1076), .A2(new_n945), .A3(new_n1077), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n1080), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(G378));
  NAND2_X1  g0909(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1078), .B1(new_n1110), .B2(new_n1056), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n405), .A2(new_n642), .ZN(new_n1112));
  XOR2_X1   g0912(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n426), .B2(new_n428), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n413), .A2(new_n424), .A3(new_n421), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n424), .B1(new_n413), .B2(new_n421), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n428), .B(new_n1114), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1112), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n428), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n1113), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1122), .A2(new_n405), .A3(new_n642), .A4(new_n1118), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n882), .B2(G330), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n650), .B(new_n1124), .C1(new_n870), .C2(new_n881), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n896), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n869), .A2(new_n871), .B1(new_n879), .B2(new_n863), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n827), .A2(new_n791), .A3(new_n868), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n890), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n874), .A2(new_n1129), .B1(new_n1131), .B2(KEYINPUT40), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1124), .B1(new_n1132), .B2(new_n650), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n889), .A2(new_n894), .A3(new_n895), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n882), .A2(G330), .A3(new_n1125), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1128), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1111), .A2(KEYINPUT57), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT116), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n889), .A2(new_n894), .A3(KEYINPUT117), .A4(new_n895), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT117), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1136), .A2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1139), .B(new_n1141), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1147), .A2(new_n1111), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n663), .B(new_n1138), .C1(new_n1148), .C2(KEYINPUT57), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1125), .A2(new_n769), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n316), .B(new_n264), .C1(new_n749), .C2(G107), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n802), .B2(new_n726), .C1(new_n310), .C2(new_n742), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n741), .A2(new_n229), .B1(new_n582), .B2(new_n737), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1153), .A2(KEYINPUT115), .B1(G77), .B2(new_n732), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(KEYINPUT115), .B2(new_n1153), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n998), .A2(new_n221), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n747), .A2(new_n210), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(new_n1152), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT58), .Z(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n216), .B1(G33), .B2(G41), .C1(new_n316), .C2(new_n264), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n921), .A2(new_n1091), .B1(new_n742), .B2(new_n813), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n995), .A2(new_n1088), .B1(new_n401), .B2(new_n741), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(G132), .C2(new_n746), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1086), .B2(new_n737), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT59), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n762), .A2(G124), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n998), .B2(new_n340), .ZN(new_n1168));
  OR3_X1    g0968(.A1(new_n1168), .A2(G33), .A3(G41), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1161), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n723), .B1(new_n1160), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n800), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1173), .A2(G50), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1150), .A2(new_n780), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1147), .B2(new_n945), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1149), .A2(new_n1176), .ZN(G375));
  NAND2_X1  g0977(.A1(new_n749), .A2(G137), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n1090), .B2(new_n737), .C1(new_n747), .C2(new_n1088), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT120), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G159), .A2(new_n756), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n257), .B(new_n1156), .C1(G128), .C2(new_n762), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n1180), .C2(new_n1179), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n804), .A2(G150), .B1(G50), .B2(new_n740), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT121), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n983), .B1(new_n756), .B2(G97), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n257), .B1(new_n921), .B2(new_n802), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n753), .B2(G77), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n746), .A2(G116), .B1(G107), .B2(new_n804), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT119), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n762), .A2(G303), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1186), .A2(new_n1188), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n737), .A2(new_n914), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1183), .A2(new_n1185), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n780), .B1(new_n1194), .B2(new_n723), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(G68), .B2(new_n1173), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT122), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n767), .B2(new_n1061), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT118), .B1(new_n1056), .B2(new_n946), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT118), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1073), .A2(new_n1201), .A3(new_n945), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1199), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1073), .A2(new_n1078), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n965), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(G381));
  NOR2_X1   g1009(.A1(G375), .A2(G378), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n787), .B(new_n1014), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(G387), .A2(G390), .A3(G384), .A4(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1208), .A3(new_n1212), .ZN(G407));
  INV_X1    g1013(.A(G343), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(G407), .A2(G213), .A3(new_n1215), .ZN(G409));
  NAND3_X1  g1016(.A1(new_n1149), .A2(G378), .A3(new_n1176), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1147), .A2(new_n965), .A3(new_n1111), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT123), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n946), .B1(new_n1128), .B2(new_n1136), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1219), .B1(new_n1220), .B2(new_n1175), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1137), .A2(new_n945), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1175), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(KEYINPUT123), .A3(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1218), .A2(new_n1221), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1108), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT124), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT124), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1225), .A2(new_n1108), .A3(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1217), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n778), .B1(new_n1205), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1056), .A2(new_n1058), .A3(KEYINPUT60), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1206), .A3(new_n1233), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1234), .A2(G384), .A3(new_n1203), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G384), .B1(new_n1234), .B2(new_n1203), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1214), .A2(G213), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1230), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(KEYINPUT62), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1230), .A2(new_n1238), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1214), .A2(G213), .A3(G2897), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1234), .A2(new_n1203), .ZN(new_n1245));
  INV_X1    g1045(.A(G384), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1234), .A2(G384), .A3(new_n1203), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1242), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1241), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT62), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1230), .A2(new_n1254), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1240), .A2(new_n1252), .A3(new_n1253), .A4(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1211), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1041), .A2(new_n663), .A3(new_n1015), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n787), .B1(new_n1258), .B2(new_n1014), .ZN(new_n1259));
  OAI21_X1  g1059(.A(KEYINPUT125), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(new_n1262), .A3(new_n1211), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(KEYINPUT126), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n981), .A2(G390), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n981), .A2(G390), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1263), .A3(new_n1260), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1260), .A2(KEYINPUT126), .A3(new_n1263), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1268), .B1(new_n1269), .B2(new_n1267), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1266), .B1(new_n1270), .B2(new_n1265), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1256), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1250), .B1(new_n1230), .B2(new_n1238), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1239), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1271), .A2(KEYINPUT61), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT127), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1239), .B2(new_n1274), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1225), .A2(new_n1108), .A3(new_n1228), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1228), .B1(new_n1225), .B2(new_n1108), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1281), .A2(new_n1217), .B1(G213), .B2(new_n1214), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1282), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1237), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1275), .A2(new_n1276), .A3(new_n1278), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1272), .A2(new_n1284), .ZN(G405));
  NAND2_X1  g1085(.A1(G375), .A2(new_n1108), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1217), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1287), .B(new_n1237), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(new_n1271), .ZN(G402));
endmodule


