//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001;
  XOR2_X1   g000(.A(KEYINPUT80), .B(KEYINPUT5), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT78), .ZN(new_n203));
  AND2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT77), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT77), .ZN(new_n210));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G148gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT76), .B1(new_n214), .B2(G141gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT76), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(G148gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(G141gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n215), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n211), .A2(KEYINPUT2), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n203), .B1(new_n213), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n212), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n224), .A2(KEYINPUT78), .A3(new_n220), .A4(new_n221), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT74), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n204), .A2(new_n205), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(KEYINPUT74), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n217), .A2(G148gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n219), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n231), .A2(KEYINPUT75), .B1(KEYINPUT2), .B2(new_n211), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT75), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n219), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n229), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n226), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(G113gat), .B(G120gat), .Z(new_n238));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g039(.A(G127gat), .B(G134gat), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n238), .B(new_n239), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(G127gat), .B(G134gat), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n239), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G120gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n243), .B(new_n244), .C1(KEYINPUT1), .C2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n237), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n226), .A2(new_n236), .A3(new_n247), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n202), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n226), .A2(new_n255), .A3(new_n236), .A4(new_n247), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT79), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n235), .B1(new_n223), .B2(new_n225), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n259), .A2(KEYINPUT79), .A3(new_n255), .A4(new_n247), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n250), .A2(KEYINPUT4), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n248), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  AOI211_X1 g063(.A(KEYINPUT3), .B(new_n235), .C1(new_n223), .C2(new_n225), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n252), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n254), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n247), .B1(new_n237), .B2(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n259), .A2(new_n263), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n253), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n202), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(new_n261), .B2(new_n256), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G1gat), .B(G29gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT0), .ZN(new_n276));
  XNOR2_X1  g075(.A(G57gat), .B(G85gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n276), .B(new_n277), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT85), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT85), .ZN(new_n281));
  AOI211_X1 g080(.A(new_n281), .B(new_n278), .C1(new_n267), .C2(new_n273), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n274), .B2(new_n279), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n288), .A2(new_n254), .B1(new_n270), .B2(new_n272), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(new_n278), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n283), .A2(new_n286), .B1(KEYINPUT6), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292));
  INV_X1    g091(.A(G169gat), .ZN(new_n293));
  INV_X1    g092(.A(G176gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G183gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(KEYINPUT27), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT27), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(G183gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT67), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(G183gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n311));
  AOI21_X1  g110(.A(G190gat), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT27), .B(G183gat), .ZN(new_n316));
  INV_X1    g115(.A(G190gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(KEYINPUT28), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n304), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n295), .A2(KEYINPUT23), .A3(new_n297), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n300), .A2(KEYINPUT23), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n321), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT24), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n317), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n320), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT25), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n305), .A2(new_n317), .A3(KEYINPUT65), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT65), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(G183gat), .B2(G190gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n324), .A2(KEYINPUT64), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT64), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n303), .A2(new_n335), .A3(new_n323), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n333), .A2(new_n334), .A3(new_n325), .A4(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(KEYINPUT23), .B2(new_n300), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT23), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n248), .B1(new_n319), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G227gat), .ZN(new_n347));
  INV_X1    g146(.A(G233gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(KEYINPUT25), .A2(new_n328), .B1(new_n337), .B2(new_n343), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n298), .A2(new_n301), .B1(G183gat), .B2(G190gat), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT28), .B1(new_n309), .B2(new_n312), .ZN(new_n353));
  INV_X1    g152(.A(new_n318), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n355), .A3(new_n247), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n346), .A2(new_n350), .A3(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G15gat), .B(G43gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n350), .B1(new_n346), .B2(new_n356), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n346), .A2(new_n356), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT33), .B1(new_n368), .B2(new_n349), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT69), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n351), .A2(new_n355), .A3(new_n247), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n247), .B1(new_n351), .B2(new_n355), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n349), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n363), .B1(new_n373), .B2(KEYINPUT32), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT69), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT33), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n373), .A2(KEYINPUT32), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n363), .A2(new_n376), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n360), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  AOI211_X1 g183(.A(new_n382), .B(new_n359), .C1(new_n370), .C2(new_n378), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT22), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT73), .B(G211gat), .ZN(new_n388));
  INV_X1    g187(.A(G218gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G197gat), .B(G204gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G211gat), .B(G218gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT29), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n259), .B1(new_n399), .B2(new_n263), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n401));
  OAI211_X1 g200(.A(G228gat), .B(G233gat), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(G22gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n397), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n265), .B2(KEYINPUT29), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n399), .A2(new_n263), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n237), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n397), .B1(new_n269), .B2(new_n398), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n410), .A2(G22gat), .A3(new_n400), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n403), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G78gat), .B(G106gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT31), .B(G50gat), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n413), .B(new_n414), .Z(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(KEYINPUT82), .ZN(new_n416));
  OAI21_X1  g215(.A(G22gat), .B1(new_n410), .B2(new_n400), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n406), .A2(new_n404), .A3(new_n408), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(new_n402), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n412), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n415), .B(KEYINPUT82), .Z(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n412), .B2(new_n419), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n386), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G226gat), .A2(G233gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n351), .A2(new_n355), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n398), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n426), .B1(new_n351), .B2(new_n355), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n405), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n427), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT29), .B1(new_n351), .B2(new_n355), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n432), .B(new_n397), .C1(new_n427), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G8gat), .B(G36gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G64gat), .B(G92gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n431), .A2(new_n434), .A3(new_n438), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(KEYINPUT30), .A3(new_n441), .ZN(new_n442));
  OR3_X1    g241(.A1(new_n435), .A2(KEYINPUT30), .A3(new_n439), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR4_X1   g244(.A1(new_n291), .A2(new_n425), .A3(KEYINPUT35), .A4(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n425), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n386), .A2(new_n424), .A3(KEYINPUT88), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n226), .A2(new_n236), .A3(new_n247), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n247), .B1(new_n226), .B2(new_n236), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n253), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n271), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n270), .B2(new_n287), .ZN(new_n455));
  INV_X1    g254(.A(new_n273), .ZN(new_n456));
  OAI211_X1 g255(.A(KEYINPUT6), .B(new_n279), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n285), .B2(new_n290), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(new_n458), .A3(new_n444), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n446), .B1(new_n459), .B2(KEYINPUT35), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  OR3_X1    g260(.A1(new_n420), .A2(new_n423), .A3(KEYINPUT83), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT83), .B1(new_n420), .B2(new_n423), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n462), .A2(new_n463), .B1(new_n458), .B2(new_n444), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT86), .B(KEYINPUT37), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n431), .A2(new_n434), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n439), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n468), .B1(new_n431), .B2(new_n434), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT38), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n469), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n439), .A4(new_n466), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n457), .A2(new_n441), .A3(new_n470), .A4(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n283), .B2(new_n286), .ZN(new_n475));
  XNOR2_X1  g274(.A(KEYINPUT84), .B(KEYINPUT40), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n256), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n255), .B1(new_n259), .B2(new_n247), .ZN(new_n479));
  OAI22_X1  g278(.A1(new_n478), .A2(new_n479), .B1(new_n264), .B2(new_n265), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n253), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n278), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n237), .A2(KEYINPUT3), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n269), .A3(new_n248), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n261), .A2(new_n256), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n252), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT39), .B1(new_n251), .B2(new_n253), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n477), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n480), .A2(new_n253), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n451), .A2(new_n452), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n481), .B1(new_n492), .B2(new_n252), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n494), .A2(KEYINPUT40), .A3(new_n278), .A4(new_n482), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n490), .A2(new_n443), .A3(new_n442), .A4(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n281), .B1(new_n289), .B2(new_n278), .ZN(new_n497));
  OAI211_X1 g296(.A(KEYINPUT85), .B(new_n279), .C1(new_n455), .C2(new_n456), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n424), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT87), .B1(new_n475), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n470), .A2(new_n473), .A3(new_n441), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(new_n457), .C1(new_n499), .C2(new_n285), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n279), .B1(new_n487), .B2(new_n481), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n476), .B1(new_n504), .B2(new_n494), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(new_n444), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n506), .A2(new_n497), .A3(new_n498), .A4(new_n495), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT87), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n503), .A2(new_n507), .A3(new_n508), .A4(new_n424), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n464), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(new_n384), .B2(new_n385), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT72), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(KEYINPUT72), .B(new_n511), .C1(new_n384), .C2(new_n385), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n367), .A2(KEYINPUT69), .A3(new_n369), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n375), .B1(new_n374), .B2(new_n377), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n383), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n359), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n379), .A2(new_n383), .A3(new_n360), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(KEYINPUT36), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT71), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n520), .A2(KEYINPUT71), .A3(KEYINPUT36), .A4(new_n521), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n516), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n461), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G57gat), .B(G64gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G71gat), .B(G78gat), .ZN(new_n533));
  INV_X1    g332(.A(G57gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT91), .A3(G64gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n537), .B(KEYINPUT92), .Z(new_n538));
  INV_X1    g337(.A(KEYINPUT9), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  OAI22_X1  g339(.A1(new_n536), .A2(new_n538), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT21), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G127gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT89), .ZN(new_n548));
  INV_X1    g347(.A(G1gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(KEYINPUT89), .A3(G1gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT16), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(G8gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n541), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(KEYINPUT21), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n546), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT93), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G155gat), .ZN(new_n561));
  XOR2_X1   g360(.A(G183gat), .B(G211gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n558), .A2(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT41), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n568), .B(new_n571), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  OAI22_X1  g374(.A1(new_n575), .A2(KEYINPUT97), .B1(new_n570), .B2(new_n569), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT8), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(KEYINPUT95), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(KEYINPUT95), .B2(new_n578), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n581), .B(KEYINPUT7), .C1(G85gat), .C2(G92gat), .ZN(new_n582));
  INV_X1    g381(.A(G85gat), .ZN(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n581), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n580), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G99gat), .B(G106gat), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n590), .A2(new_n580), .A3(new_n585), .A4(new_n586), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(KEYINPUT96), .A3(new_n591), .ZN(new_n592));
  OR3_X1    g391(.A1(new_n587), .A2(KEYINPUT96), .A3(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT14), .ZN(new_n595));
  INV_X1    g394(.A(G29gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n598));
  AOI21_X1  g397(.A(G36gat), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G36gat), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n595), .A2(new_n600), .A3(G29gat), .ZN(new_n601));
  OR3_X1    g400(.A1(new_n599), .A2(KEYINPUT15), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT15), .B1(new_n599), .B2(new_n601), .ZN(new_n603));
  XNOR2_X1  g402(.A(G43gat), .B(G50gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n576), .B1(new_n594), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT17), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n605), .B2(new_n606), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n608), .B1(new_n613), .B2(new_n594), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n575), .A2(KEYINPUT97), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT98), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n614), .A2(new_n616), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n573), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n619), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n621), .A2(new_n572), .A3(new_n617), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(G230gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(new_n348), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n556), .B1(new_n593), .B2(new_n592), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n591), .A2(KEYINPUT99), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n589), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n587), .A2(KEYINPUT99), .A3(new_n588), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n541), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n627), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n594), .A2(KEYINPUT10), .A3(new_n556), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n626), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR4_X1   g434(.A1(new_n628), .A2(new_n632), .A3(new_n625), .A4(new_n348), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OR3_X1    g439(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n640), .B1(new_n635), .B2(new_n636), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n567), .A2(new_n624), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G113gat), .B(G141gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G197gat), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT11), .B(G169gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT12), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n555), .B1(new_n611), .B2(new_n612), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT90), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n652), .A2(new_n653), .B1(new_n555), .B2(new_n607), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT90), .B1(new_n613), .B2(new_n555), .ZN(new_n655));
  NAND2_X1  g454(.A1(G229gat), .A2(G233gat), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT18), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT18), .A4(new_n656), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n555), .B(new_n607), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n656), .B(KEYINPUT13), .Z(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND4_X1   g462(.A1(new_n651), .A2(new_n659), .A3(new_n660), .A4(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(new_n657), .B2(new_n658), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n651), .B1(new_n666), .B2(new_n660), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n645), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n529), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n458), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n549), .ZN(G1324gat));
  INV_X1    g471(.A(G8gat), .ZN(new_n673));
  INV_X1    g472(.A(new_n670), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(new_n674), .B2(new_n445), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT100), .B(KEYINPUT16), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n673), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n670), .A2(new_n444), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT42), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(KEYINPUT42), .B2(new_n678), .ZN(G1325gat));
  AOI21_X1  g479(.A(G15gat), .B1(new_n674), .B2(new_n386), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT101), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n516), .A2(new_n526), .A3(KEYINPUT102), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT102), .B1(new_n516), .B2(new_n526), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n686), .A2(G15gat), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n682), .B1(new_n687), .B2(new_n674), .ZN(G1326gat));
  NAND2_X1  g487(.A1(new_n462), .A2(new_n463), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n670), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  AOI21_X1  g492(.A(new_n624), .B1(new_n461), .B2(new_n528), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n567), .A2(new_n668), .A3(new_n643), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n458), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n596), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n527), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n516), .A2(new_n526), .A3(KEYINPUT102), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n510), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT103), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n685), .A2(new_n706), .A3(new_n510), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n460), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n700), .B1(new_n708), .B2(new_n624), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT44), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n709), .A2(new_n695), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(new_n697), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n699), .B1(new_n712), .B2(new_n596), .ZN(G1328gat));
  NAND3_X1  g512(.A1(new_n696), .A2(new_n600), .A3(new_n445), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT46), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n600), .B1(new_n711), .B2(new_n445), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n715), .A2(new_n716), .ZN(G1329gat));
  NAND2_X1  g516(.A1(new_n711), .A2(new_n686), .ZN(new_n718));
  INV_X1    g517(.A(new_n386), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(G43gat), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n718), .A2(G43gat), .B1(new_n696), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g521(.A(G50gat), .ZN(new_n723));
  INV_X1    g522(.A(new_n424), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n724), .A3(new_n695), .A4(new_n710), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n723), .B1(new_n725), .B2(KEYINPUT104), .ZN(new_n726));
  AOI211_X1 g525(.A(new_n700), .B(new_n624), .C1(new_n461), .C2(new_n528), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n706), .B1(new_n685), .B2(new_n510), .ZN(new_n728));
  AND4_X1   g527(.A1(new_n706), .A2(new_n510), .A3(new_n702), .A4(new_n703), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n461), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n623), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n727), .B1(new_n731), .B2(new_n700), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n732), .A2(new_n733), .A3(new_n724), .A4(new_n695), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n726), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n696), .A2(new_n723), .A3(new_n689), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT48), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n709), .A2(new_n689), .A3(new_n695), .A4(new_n710), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G50gat), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT48), .B1(new_n742), .B2(new_n736), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n739), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n737), .B1(new_n726), .B2(new_n734), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT105), .B1(new_n746), .B2(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1331gat));
  NAND4_X1  g547(.A1(new_n567), .A2(new_n668), .A3(new_n624), .A4(new_n643), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n708), .A2(new_n458), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n534), .ZN(G1332gat));
  OR3_X1    g550(.A1(new_n708), .A2(KEYINPUT106), .A3(new_n749), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT106), .B1(new_n708), .B2(new_n749), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n444), .B(KEYINPUT107), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT108), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1333gat));
  NOR4_X1   g558(.A1(new_n708), .A2(G71gat), .A3(new_n719), .A4(new_n749), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n752), .A2(new_n686), .A3(new_n753), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(G71gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g562(.A1(new_n752), .A2(new_n689), .A3(new_n753), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g564(.A1(new_n709), .A2(new_n710), .ZN(new_n766));
  INV_X1    g565(.A(new_n668), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n567), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n644), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n697), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G85gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n705), .A2(new_n707), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n624), .B1(new_n776), .B2(new_n461), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n775), .B1(new_n777), .B2(new_n768), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n730), .A2(new_n775), .A3(new_n623), .A4(new_n768), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n781), .A2(new_n583), .A3(new_n697), .A4(new_n643), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n774), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT109), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n774), .A2(new_n785), .A3(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1336gat));
  INV_X1    g586(.A(new_n754), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n732), .A2(new_n788), .A3(new_n770), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n584), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n754), .A2(G92gat), .A3(new_n644), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(new_n781), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n766), .A2(new_n444), .A3(new_n771), .ZN(new_n796));
  INV_X1    g595(.A(new_n793), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n730), .A2(new_n623), .A3(new_n768), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(KEYINPUT110), .A3(new_n775), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n775), .A2(KEYINPUT110), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n777), .A2(new_n768), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n797), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n796), .A2(new_n584), .B1(new_n802), .B2(KEYINPUT111), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n802), .A2(KEYINPUT111), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n795), .A2(new_n805), .ZN(G1337gat));
  INV_X1    g605(.A(G99gat), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n781), .A2(new_n807), .A3(new_n386), .A4(new_n643), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n766), .A2(new_n685), .A3(new_n771), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n807), .B2(new_n809), .ZN(G1338gat));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n798), .A2(KEYINPUT51), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n424), .A2(new_n644), .A3(G106gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n779), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n732), .A2(KEYINPUT113), .A3(new_n724), .A4(new_n770), .ZN(new_n817));
  INV_X1    g616(.A(G106gat), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n709), .A2(new_n724), .A3(new_n710), .A4(new_n770), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n816), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n799), .A2(new_n801), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n813), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n709), .A2(new_n689), .A3(new_n710), .A4(new_n770), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(G106gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n815), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n811), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n817), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n814), .A2(new_n815), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n826), .ZN(new_n832));
  INV_X1    g631(.A(new_n813), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n799), .B2(new_n801), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT53), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n831), .A2(KEYINPUT114), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n828), .A2(new_n836), .ZN(G1339gat));
  NOR2_X1   g636(.A1(new_n645), .A2(new_n767), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n666), .A2(new_n651), .A3(new_n660), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n656), .B1(new_n654), .B2(new_n655), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n661), .A2(new_n662), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n649), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n623), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n635), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n633), .A2(new_n626), .A3(new_n634), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n639), .B1(new_n635), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT55), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n641), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n844), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n643), .A3(new_n843), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n668), .B2(new_n854), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n855), .B1(new_n857), .B2(new_n624), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n566), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI211_X1 g659(.A(KEYINPUT115), .B(new_n855), .C1(new_n857), .C2(new_n624), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n839), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n788), .A2(new_n458), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n862), .A2(new_n690), .A3(new_n386), .A4(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(G113gat), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n864), .A2(new_n865), .A3(new_n668), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n857), .A2(new_n624), .ZN(new_n867));
  INV_X1    g666(.A(new_n855), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n567), .B1(new_n869), .B2(KEYINPUT115), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n858), .A2(new_n859), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n838), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n458), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n873), .A2(new_n450), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(new_n754), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n767), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n866), .B1(new_n876), .B2(new_n865), .ZN(G1340gat));
  INV_X1    g676(.A(G120gat), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n864), .A2(new_n878), .A3(new_n644), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n643), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n878), .ZN(G1341gat));
  INV_X1    g680(.A(G127gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n875), .A2(new_n882), .A3(new_n567), .ZN(new_n883));
  OAI21_X1  g682(.A(G127gat), .B1(new_n864), .B2(new_n566), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1342gat));
  INV_X1    g684(.A(G134gat), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n624), .A2(new_n445), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n874), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT116), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT56), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  OAI21_X1  g691(.A(G134gat), .B1(new_n864), .B2(new_n624), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(G1343gat));
  AND2_X1   g693(.A1(new_n685), .A2(new_n863), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n862), .A2(new_n724), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n838), .B1(new_n869), .B2(new_n566), .ZN(new_n900));
  OR3_X1    g699(.A1(new_n900), .A2(new_n898), .A3(new_n690), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n897), .B1(new_n896), .B2(new_n898), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n895), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G141gat), .B1(new_n904), .B2(new_n668), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n862), .A2(new_n697), .A3(new_n724), .A4(new_n685), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n907), .B(KEYINPUT119), .Z(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n754), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n767), .A2(new_n217), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n905), .B(new_n906), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n907), .A2(new_n788), .A3(new_n910), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n904), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(KEYINPUT118), .B(new_n895), .C1(new_n902), .C2(new_n903), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n767), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n912), .B1(new_n916), .B2(G141gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n911), .B1(new_n917), .B2(new_n906), .ZN(G1344gat));
  NAND3_X1  g717(.A1(new_n862), .A2(KEYINPUT57), .A3(new_n724), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n898), .B1(new_n900), .B2(new_n690), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n644), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(new_n895), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT59), .B1(new_n924), .B2(new_n214), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n914), .A2(new_n643), .A3(new_n915), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n214), .A2(KEYINPUT59), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n908), .A2(new_n214), .A3(new_n643), .A4(new_n754), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1345gat));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n931));
  OAI21_X1  g730(.A(G155gat), .B1(new_n931), .B2(new_n566), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n567), .A2(new_n207), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n909), .B2(new_n933), .ZN(G1346gat));
  OAI21_X1  g733(.A(G162gat), .B1(new_n931), .B2(new_n624), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n908), .A2(new_n208), .A3(new_n887), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1347gat));
  NOR2_X1   g736(.A1(new_n872), .A2(new_n697), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n450), .A3(new_n788), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n293), .A3(new_n767), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n697), .A2(new_n444), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n862), .A2(new_n690), .A3(new_n386), .A4(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT120), .ZN(new_n944));
  OAI21_X1  g743(.A(G169gat), .B1(new_n944), .B2(new_n668), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n945), .A2(KEYINPUT121), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n945), .A2(KEYINPUT121), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n941), .B1(new_n946), .B2(new_n947), .ZN(G1348gat));
  OAI21_X1  g747(.A(G176gat), .B1(new_n944), .B2(new_n644), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n940), .A2(new_n294), .A3(new_n643), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1349gat));
  OAI21_X1  g750(.A(G183gat), .B1(new_n944), .B2(new_n566), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n940), .A2(new_n316), .A3(new_n567), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n317), .A3(new_n623), .ZN(new_n956));
  OAI21_X1  g755(.A(G190gat), .B1(new_n944), .B2(new_n624), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n957), .A2(KEYINPUT61), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1351gat));
  NOR3_X1   g759(.A1(new_n686), .A2(new_n424), .A3(new_n754), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n938), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(G197gat), .B1(new_n962), .B2(new_n767), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n964), .B1(new_n685), .B2(new_n942), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n685), .A2(new_n964), .A3(new_n942), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT123), .Z(new_n969));
  AND3_X1   g768(.A1(new_n921), .A2(G197gat), .A3(new_n767), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(G1352gat));
  INV_X1    g770(.A(G204gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n962), .A2(new_n972), .A3(new_n643), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT62), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n972), .B1(new_n969), .B2(new_n923), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n975), .A2(KEYINPUT124), .A3(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n979), .B1(new_n974), .B2(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1353gat));
  INV_X1    g780(.A(KEYINPUT63), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n566), .B1(new_n966), .B2(new_n967), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n921), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(G211gat), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n984), .B1(new_n921), .B2(new_n983), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n982), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(new_n987), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n989), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n985), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n962), .A2(new_n388), .A3(new_n567), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n991), .A2(KEYINPUT126), .A3(new_n992), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(G1354gat));
  AOI21_X1  g796(.A(G218gat), .B1(new_n962), .B2(new_n623), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n623), .A2(G218gat), .ZN(new_n999));
  XOR2_X1   g798(.A(new_n999), .B(KEYINPUT127), .Z(new_n1000));
  NOR2_X1   g799(.A1(new_n922), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n998), .B1(new_n969), .B2(new_n1001), .ZN(G1355gat));
endmodule


