

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750;

  XNOR2_X1 U371 ( .A(n572), .B(KEYINPUT42), .ZN(n747) );
  BUF_X1 U372 ( .A(n650), .Z(n350) );
  XNOR2_X1 U373 ( .A(n349), .B(KEYINPUT109), .ZN(n648) );
  NAND2_X1 U374 ( .A1(n443), .A2(n600), .ZN(n349) );
  XNOR2_X1 U375 ( .A(n607), .B(n365), .ZN(n650) );
  XNOR2_X1 U376 ( .A(n447), .B(G119), .ZN(n464) );
  XNOR2_X2 U377 ( .A(n724), .B(n465), .ZN(n437) );
  XNOR2_X2 U378 ( .A(n438), .B(n464), .ZN(n724) );
  INV_X4 U379 ( .A(G116), .ZN(n369) );
  XNOR2_X1 U380 ( .A(n457), .B(G107), .ZN(n725) );
  INV_X2 U381 ( .A(n615), .ZN(n682) );
  NOR2_X1 U382 ( .A1(n619), .A2(n717), .ZN(n623) );
  NOR2_X2 U383 ( .A1(n592), .A2(n350), .ZN(n564) );
  XNOR2_X2 U384 ( .A(n492), .B(KEYINPUT10), .ZN(n493) );
  XNOR2_X1 U385 ( .A(n370), .B(KEYINPUT22), .ZN(n530) );
  INV_X4 U386 ( .A(KEYINPUT4), .ZN(n367) );
  INV_X1 U387 ( .A(G125), .ZN(n469) );
  NOR2_X1 U388 ( .A1(n705), .A2(n717), .ZN(n708) );
  NOR2_X1 U389 ( .A1(n695), .A2(n717), .ZN(n371) );
  NOR2_X1 U390 ( .A1(n615), .A2(n612), .ZN(n611) );
  NAND2_X1 U391 ( .A1(n529), .A2(n667), .ZN(n631) );
  NOR2_X1 U392 ( .A1(n576), .A2(n546), .ZN(n624) );
  XNOR2_X1 U393 ( .A(n386), .B(KEYINPUT86), .ZN(n546) );
  OR2_X1 U394 ( .A1(n530), .A2(n379), .ZN(n532) );
  XNOR2_X1 U395 ( .A(n581), .B(n476), .ZN(n584) );
  AND2_X1 U396 ( .A1(n658), .A2(n659), .ZN(n662) );
  XNOR2_X1 U397 ( .A(n568), .B(n358), .ZN(n579) );
  XNOR2_X1 U398 ( .A(n456), .B(n455), .ZN(n733) );
  XNOR2_X1 U399 ( .A(n410), .B(n467), .ZN(n409) );
  XNOR2_X1 U400 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U401 ( .A(G104), .B(G110), .ZN(n457) );
  NAND2_X1 U402 ( .A1(n584), .A2(n484), .ZN(n412) );
  XNOR2_X1 U403 ( .A(n412), .B(n411), .ZN(n351) );
  INV_X1 U404 ( .A(n607), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n412), .B(n411), .ZN(n510) );
  INV_X2 U406 ( .A(n563), .ZN(n607) );
  NOR2_X2 U407 ( .A1(n535), .A2(n744), .ZN(n390) );
  OR2_X1 U408 ( .A1(n530), .A2(n418), .ZN(n417) );
  XNOR2_X2 U409 ( .A(n403), .B(n355), .ZN(n543) );
  NAND2_X1 U410 ( .A1(n428), .A2(n427), .ZN(n426) );
  NOR2_X1 U411 ( .A1(n538), .A2(n357), .ZN(n427) );
  INV_X1 U412 ( .A(n658), .ZN(n419) );
  XNOR2_X1 U413 ( .A(n528), .B(n361), .ZN(n568) );
  INV_X1 U414 ( .A(G472), .ZN(n361) );
  AND2_X1 U415 ( .A1(n426), .A2(n422), .ZN(n375) );
  NOR2_X1 U416 ( .A1(n543), .A2(n541), .ZN(n652) );
  XNOR2_X1 U417 ( .A(n354), .B(n391), .ZN(n454) );
  XNOR2_X1 U418 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n498) );
  XNOR2_X1 U419 ( .A(n466), .B(G134), .ZN(n500) );
  XNOR2_X1 U420 ( .A(n502), .B(n504), .ZN(n392) );
  INV_X1 U421 ( .A(KEYINPUT9), .ZN(n368) );
  NAND2_X1 U422 ( .A1(n398), .A2(n397), .ZN(n396) );
  INV_X1 U423 ( .A(n582), .ZN(n397) );
  INV_X1 U424 ( .A(n401), .ZN(n398) );
  XNOR2_X1 U425 ( .A(KEYINPUT111), .B(KEYINPUT36), .ZN(n582) );
  NAND2_X1 U426 ( .A1(n579), .A2(n357), .ZN(n431) );
  NAND2_X1 U427 ( .A1(n538), .A2(n357), .ZN(n430) );
  BUF_X1 U428 ( .A(n658), .Z(n377) );
  XNOR2_X1 U429 ( .A(n509), .B(n353), .ZN(n542) );
  NOR2_X1 U430 ( .A1(G902), .A2(n711), .ZN(n509) );
  INV_X1 U431 ( .A(G478), .ZN(n507) );
  AND2_X1 U432 ( .A1(n416), .A2(n419), .ZN(n415) );
  INV_X1 U433 ( .A(n568), .ZN(n667) );
  INV_X1 U434 ( .A(n377), .ZN(n576) );
  XNOR2_X1 U435 ( .A(n733), .B(n433), .ZN(n698) );
  XNOR2_X1 U436 ( .A(n465), .B(n461), .ZN(n433) );
  NOR2_X1 U437 ( .A1(n497), .A2(G952), .ZN(n717) );
  AND2_X1 U438 ( .A1(n485), .A2(G214), .ZN(n408) );
  XNOR2_X1 U439 ( .A(KEYINPUT12), .B(KEYINPUT96), .ZN(n407) );
  XNOR2_X1 U440 ( .A(G143), .B(G104), .ZN(n486) );
  NOR2_X1 U441 ( .A1(n749), .A2(n747), .ZN(n364) );
  NOR2_X1 U442 ( .A1(G902), .A2(G237), .ZN(n471) );
  XNOR2_X1 U443 ( .A(n372), .B(KEYINPUT70), .ZN(n491) );
  XNOR2_X1 U444 ( .A(KEYINPUT69), .B(G131), .ZN(n372) );
  XNOR2_X1 U445 ( .A(n406), .B(n404), .ZN(n490) );
  XNOR2_X1 U446 ( .A(n486), .B(n405), .ZN(n404) );
  XNOR2_X1 U447 ( .A(n408), .B(n407), .ZN(n406) );
  INV_X1 U448 ( .A(KEYINPUT97), .ZN(n405) );
  XNOR2_X1 U449 ( .A(G113), .B(G122), .ZN(n487) );
  XNOR2_X1 U450 ( .A(G137), .B(KEYINPUT5), .ZN(n448) );
  XOR2_X1 U451 ( .A(KEYINPUT94), .B(KEYINPUT76), .Z(n449) );
  XNOR2_X1 U452 ( .A(n451), .B(n369), .ZN(n391) );
  INV_X1 U453 ( .A(KEYINPUT48), .ZN(n363) );
  XNOR2_X1 U454 ( .A(G113), .B(KEYINPUT3), .ZN(n447) );
  XNOR2_X1 U455 ( .A(n470), .B(n468), .ZN(n410) );
  XOR2_X1 U456 ( .A(KEYINPUT88), .B(KEYINPUT17), .Z(n444) );
  INV_X1 U457 ( .A(KEYINPUT84), .ZN(n385) );
  NAND2_X1 U458 ( .A1(G234), .A2(G237), .ZN(n477) );
  INV_X1 U459 ( .A(KEYINPUT38), .ZN(n365) );
  XNOR2_X1 U460 ( .A(KEYINPUT15), .B(G902), .ZN(n612) );
  INV_X1 U461 ( .A(KEYINPUT0), .ZN(n411) );
  XOR2_X1 U462 ( .A(G137), .B(G140), .Z(n518) );
  XNOR2_X1 U463 ( .A(n366), .B(n387), .ZN(n516) );
  XNOR2_X1 U464 ( .A(n513), .B(KEYINPUT24), .ZN(n387) );
  XNOR2_X1 U465 ( .A(n514), .B(n515), .ZN(n366) );
  XNOR2_X1 U466 ( .A(G128), .B(G119), .ZN(n513) );
  XNOR2_X1 U467 ( .A(n458), .B(KEYINPUT73), .ZN(n439) );
  INV_X1 U468 ( .A(KEYINPUT41), .ZN(n440) );
  AND2_X1 U469 ( .A1(n383), .A2(n420), .ZN(n389) );
  OR2_X1 U470 ( .A1(n700), .A2(G902), .ZN(n403) );
  NAND2_X1 U471 ( .A1(n542), .A2(n543), .ZN(n577) );
  XNOR2_X1 U472 ( .A(n527), .B(KEYINPUT62), .ZN(n618) );
  XNOR2_X1 U473 ( .A(n392), .B(n503), .ZN(n505) );
  AND2_X1 U474 ( .A1(n661), .A2(n396), .ZN(n395) );
  NOR2_X1 U475 ( .A1(n414), .A2(n413), .ZN(n529) );
  NAND2_X1 U476 ( .A1(n417), .A2(n415), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n577), .B(KEYINPUT104), .ZN(n639) );
  OR2_X1 U478 ( .A1(n378), .A2(n530), .ZN(n386) );
  NAND2_X1 U479 ( .A1(n579), .A2(n583), .ZN(n378) );
  XNOR2_X1 U480 ( .A(n696), .B(n388), .ZN(n699) );
  XNOR2_X1 U481 ( .A(n698), .B(n697), .ZN(n388) );
  XOR2_X1 U482 ( .A(n508), .B(n507), .Z(n353) );
  XOR2_X1 U483 ( .A(n464), .B(n450), .Z(n354) );
  XOR2_X1 U484 ( .A(KEYINPUT13), .B(G475), .Z(n355) );
  INV_X1 U485 ( .A(n429), .ZN(n424) );
  AND2_X1 U486 ( .A1(n646), .A2(n610), .ZN(n356) );
  XOR2_X1 U487 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n357) );
  XOR2_X1 U488 ( .A(KEYINPUT101), .B(KEYINPUT6), .Z(n358) );
  INV_X1 U489 ( .A(KEYINPUT34), .ZN(n432) );
  XOR2_X1 U490 ( .A(KEYINPUT65), .B(n614), .Z(n359) );
  XOR2_X1 U491 ( .A(n693), .B(n692), .Z(n360) );
  INV_X1 U492 ( .A(n500), .ZN(n434) );
  XNOR2_X2 U493 ( .A(n526), .B(n525), .ZN(n658) );
  AND2_X2 U494 ( .A1(n362), .A2(n356), .ZN(n736) );
  XNOR2_X1 U495 ( .A(n599), .B(n363), .ZN(n362) );
  XNOR2_X1 U496 ( .A(n364), .B(KEYINPUT46), .ZN(n435) );
  XNOR2_X2 U497 ( .A(n493), .B(KEYINPUT68), .ZN(n732) );
  XNOR2_X2 U498 ( .A(n367), .B(G101), .ZN(n458) );
  XNOR2_X1 U499 ( .A(n501), .B(n368), .ZN(n502) );
  XNOR2_X2 U500 ( .A(n369), .B(G122), .ZN(n501) );
  NAND2_X1 U501 ( .A1(n373), .A2(n510), .ZN(n370) );
  XNOR2_X1 U502 ( .A(n371), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X2 U503 ( .A(n534), .B(KEYINPUT35), .ZN(n744) );
  INV_X1 U504 ( .A(n539), .ZN(n425) );
  NAND2_X1 U505 ( .A1(n435), .A2(n436), .ZN(n599) );
  XNOR2_X1 U506 ( .A(n453), .B(n454), .ZN(n527) );
  NOR2_X4 U507 ( .A1(n616), .A2(n684), .ZN(n709) );
  NOR2_X2 U508 ( .A1(n713), .A2(G902), .ZN(n526) );
  XNOR2_X1 U509 ( .A(n380), .B(n521), .ZN(n713) );
  INV_X2 U510 ( .A(n552), .ZN(n497) );
  AND2_X1 U511 ( .A1(n652), .A2(n659), .ZN(n373) );
  NAND2_X1 U512 ( .A1(n550), .A2(n549), .ZN(n376) );
  NAND2_X1 U513 ( .A1(n563), .A2(n600), .ZN(n581) );
  XNOR2_X2 U514 ( .A(n474), .B(n445), .ZN(n563) );
  INV_X1 U515 ( .A(n351), .ZN(n539) );
  AND2_X1 U516 ( .A1(n351), .A2(KEYINPUT34), .ZN(n422) );
  NAND2_X1 U517 ( .A1(n374), .A2(n590), .ZN(n534) );
  NAND2_X1 U518 ( .A1(n389), .A2(n423), .ZN(n374) );
  NOR2_X2 U519 ( .A1(n586), .A2(n674), .ZN(n572) );
  NAND2_X1 U520 ( .A1(n375), .A2(n424), .ZN(n383) );
  XNOR2_X2 U521 ( .A(n376), .B(KEYINPUT45), .ZN(n718) );
  XNOR2_X2 U522 ( .A(KEYINPUT32), .B(n532), .ZN(n745) );
  NAND2_X1 U523 ( .A1(n691), .A2(n612), .ZN(n474) );
  NOR2_X2 U524 ( .A1(G902), .A2(n698), .ZN(n462) );
  NAND2_X1 U525 ( .A1(n421), .A2(n432), .ZN(n420) );
  NAND2_X1 U526 ( .A1(n531), .A2(n579), .ZN(n379) );
  XNOR2_X1 U527 ( .A(n732), .B(n516), .ZN(n380) );
  NAND2_X1 U528 ( .A1(n381), .A2(n596), .ZN(n597) );
  NAND2_X1 U529 ( .A1(n595), .A2(KEYINPUT47), .ZN(n381) );
  NOR2_X2 U530 ( .A1(n586), .A2(n585), .ZN(n636) );
  AND2_X1 U531 ( .A1(n589), .A2(n446), .ZN(n436) );
  XNOR2_X2 U532 ( .A(n382), .B(KEYINPUT77), .ZN(n684) );
  NAND2_X1 U533 ( .A1(n682), .A2(KEYINPUT2), .ZN(n382) );
  AND2_X2 U534 ( .A1(n384), .A2(n359), .ZN(n616) );
  XNOR2_X1 U535 ( .A(n611), .B(n385), .ZN(n384) );
  XNOR2_X1 U536 ( .A(n390), .B(KEYINPUT44), .ZN(n550) );
  XNOR2_X2 U537 ( .A(G143), .B(G128), .ZN(n466) );
  NOR2_X1 U538 ( .A1(n394), .A2(n393), .ZN(n644) );
  NOR2_X1 U539 ( .A1(n402), .A2(n582), .ZN(n393) );
  NAND2_X1 U540 ( .A1(n399), .A2(n395), .ZN(n394) );
  NAND2_X1 U541 ( .A1(n402), .A2(n400), .ZN(n399) );
  AND2_X1 U542 ( .A1(n401), .A2(n582), .ZN(n400) );
  INV_X1 U543 ( .A(n581), .ZN(n401) );
  XNOR2_X1 U544 ( .A(n601), .B(KEYINPUT110), .ZN(n402) );
  INV_X1 U545 ( .A(n542), .ZN(n541) );
  XNOR2_X2 U546 ( .A(n437), .B(n409), .ZN(n691) );
  AND2_X1 U547 ( .A1(n530), .A2(KEYINPUT102), .ZN(n413) );
  NAND2_X1 U548 ( .A1(n661), .A2(KEYINPUT102), .ZN(n416) );
  OR2_X1 U549 ( .A1(n661), .A2(KEYINPUT102), .ZN(n418) );
  XNOR2_X2 U550 ( .A(KEYINPUT64), .B(G953), .ZN(n552) );
  NAND2_X1 U551 ( .A1(n426), .A2(n425), .ZN(n421) );
  NAND2_X1 U552 ( .A1(n429), .A2(n432), .ZN(n423) );
  NAND2_X1 U553 ( .A1(n424), .A2(n426), .ZN(n657) );
  INV_X1 U554 ( .A(n579), .ZN(n428) );
  NAND2_X1 U555 ( .A1(n431), .A2(n430), .ZN(n429) );
  XNOR2_X2 U556 ( .A(n434), .B(n491), .ZN(n456) );
  XNOR2_X2 U557 ( .A(n501), .B(KEYINPUT16), .ZN(n438) );
  XNOR2_X2 U558 ( .A(n439), .B(n725), .ZN(n465) );
  XNOR2_X2 U559 ( .A(n441), .B(n440), .ZN(n674) );
  NAND2_X1 U560 ( .A1(n648), .A2(n652), .ZN(n441) );
  INV_X1 U561 ( .A(n650), .ZN(n443) );
  BUF_X1 U562 ( .A(n709), .Z(n714) );
  NAND2_X1 U563 ( .A1(n718), .A2(n736), .ZN(n615) );
  XNOR2_X2 U564 ( .A(n570), .B(KEYINPUT1), .ZN(n661) );
  XNOR2_X2 U565 ( .A(n463), .B(n462), .ZN(n570) );
  XNOR2_X1 U566 ( .A(n473), .B(n472), .ZN(n445) );
  XNOR2_X1 U567 ( .A(KEYINPUT82), .B(n598), .ZN(n446) );
  XNOR2_X1 U568 ( .A(n492), .B(n444), .ZN(n470) );
  INV_X1 U569 ( .A(n750), .ZN(n610) );
  XNOR2_X1 U570 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U571 ( .A(n702), .B(n701), .ZN(n703) );
  INV_X1 U572 ( .A(KEYINPUT87), .ZN(n620) );
  INV_X1 U573 ( .A(n639), .ZN(n637) );
  XNOR2_X1 U574 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U575 ( .A(n449), .B(n448), .ZN(n450) );
  NOR2_X1 U576 ( .A1(G953), .A2(G237), .ZN(n485) );
  NAND2_X1 U577 ( .A1(n485), .A2(G210), .ZN(n451) );
  XNOR2_X1 U578 ( .A(n458), .B(G146), .ZN(n452) );
  XNOR2_X1 U579 ( .A(n456), .B(n452), .ZN(n453) );
  XNOR2_X1 U580 ( .A(KEYINPUT71), .B(G469), .ZN(n463) );
  INV_X1 U581 ( .A(n518), .ZN(n455) );
  XOR2_X1 U582 ( .A(G146), .B(KEYINPUT80), .Z(n460) );
  NAND2_X1 U583 ( .A1(G227), .A2(n497), .ZN(n459) );
  XNOR2_X1 U584 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U585 ( .A(KEYINPUT79), .B(KEYINPUT19), .Z(n476) );
  XNOR2_X1 U586 ( .A(n466), .B(KEYINPUT18), .ZN(n468) );
  NAND2_X1 U587 ( .A1(G224), .A2(n497), .ZN(n467) );
  XNOR2_X2 U588 ( .A(n469), .B(G146), .ZN(n492) );
  XOR2_X1 U589 ( .A(KEYINPUT81), .B(KEYINPUT89), .Z(n473) );
  XNOR2_X1 U590 ( .A(n471), .B(KEYINPUT75), .ZN(n475) );
  NAND2_X1 U591 ( .A1(G210), .A2(n475), .ZN(n472) );
  NAND2_X1 U592 ( .A1(G214), .A2(n475), .ZN(n600) );
  INV_X1 U593 ( .A(G953), .ZN(n719) );
  NOR2_X1 U594 ( .A1(G898), .A2(n719), .ZN(n729) );
  XNOR2_X1 U595 ( .A(n477), .B(KEYINPUT90), .ZN(n478) );
  XNOR2_X1 U596 ( .A(KEYINPUT14), .B(n478), .ZN(n480) );
  NAND2_X1 U597 ( .A1(G902), .A2(n480), .ZN(n551) );
  INV_X1 U598 ( .A(n551), .ZN(n479) );
  NAND2_X1 U599 ( .A1(n729), .A2(n479), .ZN(n483) );
  NAND2_X1 U600 ( .A1(n480), .A2(G952), .ZN(n481) );
  XOR2_X1 U601 ( .A(KEYINPUT91), .B(n481), .Z(n681) );
  NOR2_X1 U602 ( .A1(G953), .A2(n681), .ZN(n556) );
  INV_X1 U603 ( .A(n556), .ZN(n482) );
  NAND2_X1 U604 ( .A1(n483), .A2(n482), .ZN(n484) );
  XOR2_X1 U605 ( .A(KEYINPUT11), .B(G140), .Z(n488) );
  XNOR2_X1 U606 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U607 ( .A(n490), .B(n489), .Z(n496) );
  INV_X1 U608 ( .A(n491), .ZN(n494) );
  XOR2_X1 U609 ( .A(n494), .B(n732), .Z(n495) );
  XNOR2_X1 U610 ( .A(n496), .B(n495), .ZN(n700) );
  NAND2_X1 U611 ( .A1(n497), .A2(G234), .ZN(n499) );
  XNOR2_X1 U612 ( .A(n499), .B(n498), .ZN(n517) );
  NAND2_X1 U613 ( .A1(n517), .A2(G217), .ZN(n506) );
  XNOR2_X1 U614 ( .A(n500), .B(G107), .ZN(n503) );
  XOR2_X1 U615 ( .A(KEYINPUT7), .B(KEYINPUT98), .Z(n504) );
  XOR2_X1 U616 ( .A(n506), .B(n505), .Z(n711) );
  INV_X1 U617 ( .A(KEYINPUT99), .ZN(n508) );
  NAND2_X1 U618 ( .A1(G234), .A2(n612), .ZN(n511) );
  XNOR2_X1 U619 ( .A(KEYINPUT20), .B(n511), .ZN(n522) );
  NAND2_X1 U620 ( .A1(G221), .A2(n522), .ZN(n512) );
  XOR2_X1 U621 ( .A(n512), .B(KEYINPUT21), .Z(n659) );
  INV_X1 U622 ( .A(n659), .ZN(n574) );
  XOR2_X1 U623 ( .A(KEYINPUT72), .B(G110), .Z(n514) );
  INV_X1 U624 ( .A(KEYINPUT92), .ZN(n515) );
  NAND2_X1 U625 ( .A1(n517), .A2(G221), .ZN(n520) );
  XNOR2_X1 U626 ( .A(n518), .B(KEYINPUT23), .ZN(n519) );
  NAND2_X1 U627 ( .A1(G217), .A2(n522), .ZN(n524) );
  XOR2_X1 U628 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n523) );
  NOR2_X1 U629 ( .A1(G902), .A2(n527), .ZN(n528) );
  INV_X1 U630 ( .A(n661), .ZN(n583) );
  NOR2_X1 U631 ( .A1(n377), .A2(n583), .ZN(n531) );
  NAND2_X1 U632 ( .A1(n631), .A2(n745), .ZN(n535) );
  NAND2_X1 U633 ( .A1(n661), .A2(n662), .ZN(n538) );
  NAND2_X1 U634 ( .A1(n541), .A2(n543), .ZN(n533) );
  XNOR2_X1 U635 ( .A(n533), .B(KEYINPUT103), .ZN(n590) );
  NAND2_X1 U636 ( .A1(n570), .A2(n662), .ZN(n557) );
  NOR2_X1 U637 ( .A1(n539), .A2(n557), .ZN(n536) );
  NAND2_X1 U638 ( .A1(n667), .A2(n536), .ZN(n537) );
  XOR2_X1 U639 ( .A(KEYINPUT95), .B(n537), .Z(n628) );
  OR2_X1 U640 ( .A1(n667), .A2(n538), .ZN(n670) );
  NOR2_X1 U641 ( .A1(n670), .A2(n539), .ZN(n540) );
  XNOR2_X1 U642 ( .A(n540), .B(KEYINPUT31), .ZN(n641) );
  NAND2_X1 U643 ( .A1(n628), .A2(n641), .ZN(n544) );
  NOR2_X1 U644 ( .A1(n543), .A2(n542), .ZN(n632) );
  INV_X1 U645 ( .A(n632), .ZN(n642) );
  NAND2_X1 U646 ( .A1(n642), .A2(n577), .ZN(n649) );
  NAND2_X1 U647 ( .A1(n544), .A2(n649), .ZN(n545) );
  XNOR2_X1 U648 ( .A(n545), .B(KEYINPUT100), .ZN(n548) );
  INV_X1 U649 ( .A(n624), .ZN(n547) );
  AND2_X1 U650 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U651 ( .A1(G900), .A2(n551), .ZN(n553) );
  NAND2_X1 U652 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U653 ( .A(KEYINPUT105), .B(n554), .ZN(n555) );
  NOR2_X1 U654 ( .A1(n556), .A2(n555), .ZN(n573) );
  NOR2_X2 U655 ( .A1(n557), .A2(n573), .ZN(n558) );
  XNOR2_X1 U656 ( .A(n558), .B(KEYINPUT78), .ZN(n562) );
  XOR2_X1 U657 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n560) );
  NAND2_X1 U658 ( .A1(n568), .A2(n600), .ZN(n559) );
  XNOR2_X1 U659 ( .A(n560), .B(n559), .ZN(n561) );
  NAND2_X1 U660 ( .A1(n562), .A2(n561), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n564), .B(KEYINPUT39), .ZN(n608) );
  NOR2_X1 U662 ( .A1(n577), .A2(n608), .ZN(n565) );
  XNOR2_X1 U663 ( .A(n565), .B(KEYINPUT40), .ZN(n749) );
  NAND2_X1 U664 ( .A1(n419), .A2(n659), .ZN(n566) );
  NOR2_X1 U665 ( .A1(n573), .A2(n566), .ZN(n567) );
  AND2_X1 U666 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U667 ( .A(KEYINPUT28), .B(n569), .ZN(n571) );
  NAND2_X1 U668 ( .A1(n571), .A2(n570), .ZN(n586) );
  INV_X1 U669 ( .A(n600), .ZN(n651) );
  NOR2_X1 U670 ( .A1(n574), .A2(n573), .ZN(n575) );
  AND2_X1 U671 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U672 ( .A1(n578), .A2(n637), .ZN(n580) );
  NOR2_X1 U673 ( .A1(n580), .A2(n579), .ZN(n601) );
  INV_X1 U674 ( .A(n584), .ZN(n585) );
  NAND2_X1 U675 ( .A1(n649), .A2(n636), .ZN(n587) );
  NOR2_X1 U676 ( .A1(KEYINPUT47), .A2(n587), .ZN(n588) );
  NOR2_X1 U677 ( .A1(n644), .A2(n588), .ZN(n589) );
  NAND2_X1 U678 ( .A1(n352), .A2(n590), .ZN(n591) );
  NOR2_X1 U679 ( .A1(n592), .A2(n591), .ZN(n635) );
  INV_X1 U680 ( .A(n649), .ZN(n593) );
  NAND2_X1 U681 ( .A1(n593), .A2(KEYINPUT47), .ZN(n594) );
  XOR2_X1 U682 ( .A(n594), .B(KEYINPUT83), .Z(n596) );
  INV_X1 U683 ( .A(n636), .ZN(n595) );
  NOR2_X1 U684 ( .A1(n635), .A2(n597), .ZN(n598) );
  NAND2_X1 U685 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U686 ( .A(KEYINPUT106), .B(n602), .ZN(n603) );
  NOR2_X1 U687 ( .A1(n661), .A2(n603), .ZN(n605) );
  XNOR2_X1 U688 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n604) );
  XNOR2_X1 U689 ( .A(n605), .B(n604), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n646) );
  OR2_X1 U691 ( .A1(n642), .A2(n608), .ZN(n609) );
  XOR2_X1 U692 ( .A(KEYINPUT112), .B(n609), .Z(n750) );
  XNOR2_X1 U693 ( .A(KEYINPUT85), .B(n612), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n613), .A2(KEYINPUT2), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n709), .A2(G472), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U697 ( .A(KEYINPUT113), .B(KEYINPUT63), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n623), .B(n622), .ZN(G57) );
  XOR2_X1 U699 ( .A(n624), .B(G101), .Z(G3) );
  NOR2_X1 U700 ( .A1(n639), .A2(n628), .ZN(n625) );
  XOR2_X1 U701 ( .A(G104), .B(n625), .Z(G6) );
  XOR2_X1 U702 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n627) );
  XNOR2_X1 U703 ( .A(G107), .B(KEYINPUT114), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n627), .B(n626), .ZN(n630) );
  NOR2_X1 U705 ( .A1(n642), .A2(n628), .ZN(n629) );
  XOR2_X1 U706 ( .A(n630), .B(n629), .Z(G9) );
  XNOR2_X1 U707 ( .A(n631), .B(G110), .ZN(G12) );
  XOR2_X1 U708 ( .A(G128), .B(KEYINPUT29), .Z(n634) );
  NAND2_X1 U709 ( .A1(n636), .A2(n632), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n634), .B(n633), .ZN(G30) );
  XOR2_X1 U711 ( .A(G143), .B(n635), .Z(G45) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U713 ( .A(n638), .B(G146), .ZN(G48) );
  NOR2_X1 U714 ( .A1(n639), .A2(n641), .ZN(n640) );
  XOR2_X1 U715 ( .A(G113), .B(n640), .Z(G15) );
  NOR2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U717 ( .A(G116), .B(n643), .Z(G18) );
  XNOR2_X1 U718 ( .A(n644), .B(G125), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n645), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U720 ( .A(G140), .B(n646), .ZN(G42) );
  NOR2_X1 U721 ( .A1(n657), .A2(n674), .ZN(n647) );
  NOR2_X1 U722 ( .A1(G953), .A2(n647), .ZN(n688) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n651), .A2(n350), .ZN(n653) );
  NAND2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n654) );
  AND2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n677) );
  NOR2_X1 U728 ( .A1(n659), .A2(n377), .ZN(n660) );
  XOR2_X1 U729 ( .A(KEYINPUT49), .B(n660), .Z(n666) );
  OR2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n663), .B(KEYINPUT50), .ZN(n664) );
  XNOR2_X1 U732 ( .A(KEYINPUT115), .B(n664), .ZN(n665) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n668) );
  NAND2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n669), .B(KEYINPUT116), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n673) );
  XOR2_X1 U737 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n672) );
  XNOR2_X1 U738 ( .A(n673), .B(n672), .ZN(n675) );
  NOR2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U740 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U741 ( .A(n678), .B(KEYINPUT118), .ZN(n679) );
  XNOR2_X1 U742 ( .A(KEYINPUT52), .B(n679), .ZN(n680) );
  NOR2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n686) );
  NOR2_X1 U744 ( .A1(n682), .A2(KEYINPUT2), .ZN(n683) );
  NOR2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U748 ( .A(n689), .B(KEYINPUT53), .ZN(n690) );
  XNOR2_X1 U749 ( .A(KEYINPUT119), .B(n690), .ZN(G75) );
  NAND2_X1 U750 ( .A1(n709), .A2(G210), .ZN(n694) );
  XOR2_X1 U751 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n693) );
  XNOR2_X1 U752 ( .A(n691), .B(KEYINPUT55), .ZN(n692) );
  XNOR2_X1 U753 ( .A(n694), .B(n360), .ZN(n695) );
  XOR2_X1 U754 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n697) );
  NAND2_X1 U755 ( .A1(n714), .A2(G469), .ZN(n696) );
  NOR2_X1 U756 ( .A1(n717), .A2(n699), .ZN(G54) );
  NAND2_X1 U757 ( .A1(n709), .A2(G475), .ZN(n704) );
  INV_X1 U758 ( .A(n700), .ZN(n702) );
  XOR2_X1 U759 ( .A(KEYINPUT59), .B(KEYINPUT121), .Z(n701) );
  XNOR2_X1 U760 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U761 ( .A(KEYINPUT66), .B(KEYINPUT122), .ZN(n706) );
  XNOR2_X1 U762 ( .A(n706), .B(KEYINPUT60), .ZN(n707) );
  XNOR2_X1 U763 ( .A(n708), .B(n707), .ZN(G60) );
  NAND2_X1 U764 ( .A1(G478), .A2(n714), .ZN(n710) );
  XNOR2_X1 U765 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n717), .A2(n712), .ZN(G63) );
  NAND2_X1 U767 ( .A1(G217), .A2(n714), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n713), .B(n715), .ZN(n716) );
  NOR2_X1 U769 ( .A1(n717), .A2(n716), .ZN(G66) );
  NAND2_X1 U770 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U771 ( .A1(G953), .A2(G224), .ZN(n720) );
  XNOR2_X1 U772 ( .A(KEYINPUT61), .B(n720), .ZN(n721) );
  NAND2_X1 U773 ( .A1(n721), .A2(G898), .ZN(n722) );
  NAND2_X1 U774 ( .A1(n723), .A2(n722), .ZN(n731) );
  XNOR2_X1 U775 ( .A(n724), .B(n725), .ZN(n726) );
  XNOR2_X1 U776 ( .A(n726), .B(KEYINPUT123), .ZN(n727) );
  XNOR2_X1 U777 ( .A(n727), .B(G101), .ZN(n728) );
  NOR2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U779 ( .A(n731), .B(n730), .ZN(G69) );
  XNOR2_X1 U780 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U781 ( .A(n734), .B(KEYINPUT124), .ZN(n735) );
  XNOR2_X1 U782 ( .A(KEYINPUT4), .B(n735), .ZN(n738) );
  XOR2_X1 U783 ( .A(n736), .B(n738), .Z(n737) );
  NAND2_X1 U784 ( .A1(n737), .A2(n497), .ZN(n743) );
  XNOR2_X1 U785 ( .A(G227), .B(n738), .ZN(n739) );
  NAND2_X1 U786 ( .A1(n739), .A2(G900), .ZN(n740) );
  XOR2_X1 U787 ( .A(KEYINPUT125), .B(n740), .Z(n741) );
  NAND2_X1 U788 ( .A1(G953), .A2(n741), .ZN(n742) );
  NAND2_X1 U789 ( .A1(n743), .A2(n742), .ZN(G72) );
  XOR2_X1 U790 ( .A(n744), .B(G122), .Z(G24) );
  XNOR2_X1 U791 ( .A(n745), .B(G119), .ZN(n746) );
  XNOR2_X1 U792 ( .A(n746), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U793 ( .A(G137), .B(KEYINPUT127), .ZN(n748) );
  XNOR2_X1 U794 ( .A(n748), .B(n747), .ZN(G39) );
  XOR2_X1 U795 ( .A(n749), .B(G131), .Z(G33) );
  XOR2_X1 U796 ( .A(G134), .B(n750), .Z(G36) );
endmodule

