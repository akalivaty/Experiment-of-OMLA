

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U326 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U327 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n431) );
  XNOR2_X1 U328 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U329 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U330 ( .A(n429), .B(KEYINPUT48), .ZN(n543) );
  NOR2_X1 U331 ( .A1(n528), .A2(n453), .ZN(n563) );
  XNOR2_X1 U332 ( .A(n455), .B(KEYINPUT122), .ZN(n456) );
  XNOR2_X1 U333 ( .A(n457), .B(n456), .ZN(G1350GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n295) );
  XNOR2_X1 U335 ( .A(G8GAT), .B(KEYINPUT15), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n309) );
  XOR2_X1 U337 ( .A(G64GAT), .B(G127GAT), .Z(n297) );
  NAND2_X1 U338 ( .A1(G231GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n299) );
  XNOR2_X1 U340 ( .A(G183GAT), .B(G211GAT), .ZN(n298) );
  XNOR2_X1 U341 ( .A(n298), .B(KEYINPUT81), .ZN(n358) );
  XOR2_X1 U342 ( .A(n299), .B(n358), .Z(n303) );
  XNOR2_X1 U343 ( .A(G15GAT), .B(G1GAT), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n300), .B(KEYINPUT71), .ZN(n390) );
  XNOR2_X1 U345 ( .A(G71GAT), .B(G57GAT), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n301), .B(KEYINPUT13), .ZN(n401) );
  XNOR2_X1 U347 ( .A(n390), .B(n401), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U349 ( .A(n304), .B(KEYINPUT12), .Z(n307) );
  XNOR2_X1 U350 ( .A(G22GAT), .B(G155GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n305), .B(G78GAT), .ZN(n436) );
  XNOR2_X1 U352 ( .A(n436), .B(KEYINPUT14), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n578) );
  XNOR2_X1 U355 ( .A(KEYINPUT113), .B(n578), .ZN(n535) );
  XOR2_X1 U356 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n311) );
  XNOR2_X1 U357 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U359 ( .A(n312), .B(G127GAT), .Z(n314) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(G120GAT), .ZN(n313) );
  XNOR2_X1 U361 ( .A(n314), .B(n313), .ZN(n349) );
  XOR2_X1 U362 ( .A(G71GAT), .B(G176GAT), .Z(n316) );
  XNOR2_X1 U363 ( .A(G169GAT), .B(G183GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n349), .B(n317), .ZN(n330) );
  XOR2_X1 U366 ( .A(KEYINPUT91), .B(G190GAT), .Z(n319) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G99GAT), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n328) );
  XNOR2_X1 U369 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n320), .B(KEYINPUT17), .ZN(n359) );
  XOR2_X1 U371 ( .A(n359), .B(G15GAT), .Z(n322) );
  NAND2_X1 U372 ( .A1(G227GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U374 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n324) );
  XNOR2_X1 U375 ( .A(KEYINPUT90), .B(KEYINPUT20), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U377 ( .A(n326), .B(n325), .Z(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n528) );
  XOR2_X1 U380 ( .A(KEYINPUT96), .B(KEYINPUT1), .Z(n332) );
  XNOR2_X1 U381 ( .A(G1GAT), .B(G57GAT), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U383 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n334) );
  XNOR2_X1 U384 ( .A(G155GAT), .B(G148GAT), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n347) );
  XOR2_X1 U387 ( .A(KEYINPUT4), .B(KEYINPUT97), .Z(n338) );
  NAND2_X1 U388 ( .A1(G225GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U390 ( .A(n339), .B(G85GAT), .Z(n345) );
  XNOR2_X1 U391 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n340), .B(KEYINPUT94), .ZN(n341) );
  XOR2_X1 U393 ( .A(n341), .B(KEYINPUT93), .Z(n343) );
  XNOR2_X1 U394 ( .A(G141GAT), .B(G162GAT), .ZN(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n441) );
  XNOR2_X1 U396 ( .A(G29GAT), .B(n441), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n349), .B(n348), .ZN(n515) );
  XOR2_X1 U400 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n351) );
  NAND2_X1 U401 ( .A1(G226GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U403 ( .A(n352), .B(KEYINPUT98), .Z(n357) );
  XNOR2_X1 U404 ( .A(G169GAT), .B(G36GAT), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n353), .B(G8GAT), .ZN(n386) );
  XOR2_X1 U406 ( .A(G64GAT), .B(G92GAT), .Z(n355) );
  XNOR2_X1 U407 ( .A(G176GAT), .B(G204GAT), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n398) );
  XNOR2_X1 U409 ( .A(n386), .B(n398), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n363) );
  XOR2_X1 U411 ( .A(G190GAT), .B(G218GAT), .Z(n366) );
  XOR2_X1 U412 ( .A(n358), .B(n366), .Z(n361) );
  XOR2_X1 U413 ( .A(G197GAT), .B(KEYINPUT21), .Z(n437) );
  XNOR2_X1 U414 ( .A(n359), .B(n437), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n517) );
  XOR2_X1 U417 ( .A(KEYINPUT119), .B(n517), .Z(n430) );
  XOR2_X1 U418 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n365) );
  XNOR2_X1 U419 ( .A(KEYINPUT11), .B(KEYINPUT80), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n367) );
  XOR2_X1 U421 ( .A(n367), .B(n366), .Z(n369) );
  XNOR2_X1 U422 ( .A(G36GAT), .B(G92GAT), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n374) );
  XNOR2_X1 U424 ( .A(G99GAT), .B(G106GAT), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n370), .B(G85GAT), .ZN(n399) );
  XOR2_X1 U426 ( .A(KEYINPUT66), .B(n399), .Z(n372) );
  NAND2_X1 U427 ( .A1(G232GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U429 ( .A(n374), .B(n373), .Z(n383) );
  XNOR2_X1 U430 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n375), .B(G29GAT), .ZN(n376) );
  XOR2_X1 U432 ( .A(n376), .B(KEYINPUT7), .Z(n378) );
  XNOR2_X1 U433 ( .A(G50GAT), .B(KEYINPUT70), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n395) );
  XOR2_X1 U435 ( .A(KEYINPUT9), .B(KEYINPUT78), .Z(n380) );
  XNOR2_X1 U436 ( .A(G134GAT), .B(G162GAT), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n395), .B(n381), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n562) );
  XOR2_X1 U440 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n389) );
  XOR2_X1 U441 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n385) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(G141GAT), .ZN(n384) );
  XNOR2_X1 U443 ( .A(n385), .B(n384), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n394) );
  XOR2_X1 U446 ( .A(G22GAT), .B(n390), .Z(n392) );
  NAND2_X1 U447 ( .A1(G229GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U449 ( .A(n394), .B(n393), .Z(n397) );
  XNOR2_X1 U450 ( .A(n395), .B(G113GAT), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n571) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n417) );
  XOR2_X1 U453 ( .A(KEYINPUT76), .B(G148GAT), .Z(n445) );
  INV_X1 U454 ( .A(n445), .ZN(n400) );
  NAND2_X1 U455 ( .A1(n401), .A2(n400), .ZN(n404) );
  INV_X1 U456 ( .A(n401), .ZN(n402) );
  NAND2_X1 U457 ( .A1(n402), .A2(n445), .ZN(n403) );
  NAND2_X1 U458 ( .A1(n404), .A2(n403), .ZN(n406) );
  XNOR2_X1 U459 ( .A(G120GAT), .B(G78GAT), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n415) );
  XOR2_X1 U461 ( .A(KEYINPUT31), .B(KEYINPUT73), .Z(n408) );
  XNOR2_X1 U462 ( .A(KEYINPUT77), .B(KEYINPUT33), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n409), .B(KEYINPUT74), .ZN(n413) );
  XOR2_X1 U465 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n411) );
  NAND2_X1 U466 ( .A1(G230GAT), .A2(G233GAT), .ZN(n410) );
  XOR2_X1 U467 ( .A(n411), .B(n410), .Z(n412) );
  XNOR2_X1 U468 ( .A(n417), .B(n416), .ZN(n574) );
  XNOR2_X1 U469 ( .A(n574), .B(KEYINPUT64), .ZN(n418) );
  XNOR2_X1 U470 ( .A(n418), .B(KEYINPUT41), .ZN(n557) );
  NAND2_X1 U471 ( .A1(n571), .A2(n557), .ZN(n419) );
  XNOR2_X1 U472 ( .A(KEYINPUT46), .B(n419), .ZN(n420) );
  NAND2_X1 U473 ( .A1(n420), .A2(n535), .ZN(n421) );
  NOR2_X1 U474 ( .A1(n562), .A2(n421), .ZN(n422) );
  XNOR2_X1 U475 ( .A(n422), .B(KEYINPUT47), .ZN(n428) );
  XNOR2_X1 U476 ( .A(n571), .B(KEYINPUT72), .ZN(n555) );
  XOR2_X1 U477 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n424) );
  XNOR2_X1 U478 ( .A(KEYINPUT36), .B(n562), .ZN(n582) );
  NAND2_X1 U479 ( .A1(n578), .A2(n582), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  NOR2_X1 U481 ( .A1(n555), .A2(n425), .ZN(n426) );
  NAND2_X1 U482 ( .A1(n574), .A2(n426), .ZN(n427) );
  NAND2_X1 U483 ( .A1(n428), .A2(n427), .ZN(n429) );
  NAND2_X1 U484 ( .A1(n430), .A2(n543), .ZN(n432) );
  NOR2_X1 U485 ( .A1(n515), .A2(n433), .ZN(n568) );
  XOR2_X1 U486 ( .A(G204GAT), .B(KEYINPUT22), .Z(n435) );
  XNOR2_X1 U487 ( .A(KEYINPUT95), .B(KEYINPUT23), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n451) );
  XOR2_X1 U489 ( .A(n437), .B(n436), .Z(n439) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n449) );
  XOR2_X1 U493 ( .A(G211GAT), .B(KEYINPUT24), .Z(n443) );
  XNOR2_X1 U494 ( .A(G106GAT), .B(KEYINPUT92), .ZN(n442) );
  XNOR2_X1 U495 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U496 ( .A(n444), .B(G218GAT), .Z(n447) );
  XNOR2_X1 U497 ( .A(G50GAT), .B(n445), .ZN(n446) );
  XNOR2_X1 U498 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U500 ( .A(n451), .B(n450), .ZN(n467) );
  NAND2_X1 U501 ( .A1(n568), .A2(n467), .ZN(n452) );
  XOR2_X1 U502 ( .A(n452), .B(KEYINPUT55), .Z(n453) );
  INV_X1 U503 ( .A(n563), .ZN(n454) );
  NOR2_X1 U504 ( .A1(n535), .A2(n454), .ZN(n457) );
  INV_X1 U505 ( .A(G183GAT), .ZN(n455) );
  NAND2_X1 U506 ( .A1(n574), .A2(n555), .ZN(n491) );
  INV_X1 U507 ( .A(n562), .ZN(n458) );
  NAND2_X1 U508 ( .A1(n458), .A2(n578), .ZN(n461) );
  XNOR2_X1 U509 ( .A(KEYINPUT16), .B(KEYINPUT85), .ZN(n459) );
  XNOR2_X1 U510 ( .A(n459), .B(KEYINPUT84), .ZN(n460) );
  XNOR2_X1 U511 ( .A(n461), .B(n460), .ZN(n476) );
  INV_X1 U512 ( .A(n528), .ZN(n519) );
  XNOR2_X1 U513 ( .A(n517), .B(KEYINPUT27), .ZN(n469) );
  NAND2_X1 U514 ( .A1(n469), .A2(n515), .ZN(n545) );
  XNOR2_X1 U515 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n462), .B(n467), .ZN(n522) );
  NOR2_X1 U517 ( .A1(n545), .A2(n522), .ZN(n527) );
  XNOR2_X1 U518 ( .A(KEYINPUT101), .B(n527), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n519), .A2(n463), .ZN(n474) );
  NAND2_X1 U520 ( .A1(n517), .A2(n519), .ZN(n464) );
  NAND2_X1 U521 ( .A1(n464), .A2(n467), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n465), .B(KEYINPUT102), .ZN(n466) );
  XNOR2_X1 U523 ( .A(KEYINPUT25), .B(n466), .ZN(n471) );
  NOR2_X1 U524 ( .A1(n467), .A2(n519), .ZN(n468) );
  XNOR2_X1 U525 ( .A(n468), .B(KEYINPUT26), .ZN(n569) );
  AND2_X1 U526 ( .A1(n569), .A2(n469), .ZN(n470) );
  NOR2_X1 U527 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U528 ( .A1(n515), .A2(n472), .ZN(n473) );
  NOR2_X1 U529 ( .A1(n474), .A2(n473), .ZN(n486) );
  INV_X1 U530 ( .A(n486), .ZN(n475) );
  NAND2_X1 U531 ( .A1(n476), .A2(n475), .ZN(n503) );
  NOR2_X1 U532 ( .A1(n491), .A2(n503), .ZN(n477) );
  XOR2_X1 U533 ( .A(KEYINPUT103), .B(n477), .Z(n483) );
  NAND2_X1 U534 ( .A1(n515), .A2(n483), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n478), .B(KEYINPUT34), .ZN(n479) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n479), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n517), .A2(n483), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .Z(n482) );
  NAND2_X1 U540 ( .A1(n483), .A2(n519), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(G1326GAT) );
  NAND2_X1 U542 ( .A1(n522), .A2(n483), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(KEYINPUT104), .ZN(n485) );
  XNOR2_X1 U544 ( .A(G22GAT), .B(n485), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT106), .B(KEYINPUT37), .Z(n490) );
  NOR2_X1 U546 ( .A1(n486), .A2(n578), .ZN(n487) );
  XOR2_X1 U547 ( .A(KEYINPUT105), .B(n487), .Z(n488) );
  NAND2_X1 U548 ( .A1(n488), .A2(n582), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(n512) );
  NOR2_X1 U550 ( .A1(n512), .A2(n491), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n492), .B(KEYINPUT38), .ZN(n498) );
  NAND2_X1 U552 ( .A1(n515), .A2(n498), .ZN(n494) );
  XOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n498), .A2(n517), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n498), .A2(n519), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  XOR2_X1 U560 ( .A(G50GAT), .B(KEYINPUT107), .Z(n500) );
  NAND2_X1 U561 ( .A1(n498), .A2(n522), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(G1331GAT) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n506) );
  INV_X1 U564 ( .A(n571), .ZN(n501) );
  NAND2_X1 U565 ( .A1(n501), .A2(n557), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(KEYINPUT108), .ZN(n513) );
  NOR2_X1 U567 ( .A1(n513), .A2(n503), .ZN(n504) );
  XOR2_X1 U568 ( .A(KEYINPUT109), .B(n504), .Z(n509) );
  NAND2_X1 U569 ( .A1(n509), .A2(n515), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n517), .A2(n509), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n509), .A2(n519), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U576 ( .A1(n509), .A2(n522), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NOR2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(KEYINPUT110), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n515), .A2(n523), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n523), .A2(n517), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U584 ( .A(G99GAT), .B(KEYINPUT111), .Z(n521) );
  NAND2_X1 U585 ( .A1(n519), .A2(n523), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1338GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n525) );
  NAND2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U590 ( .A(G106GAT), .B(n526), .Z(G1339GAT) );
  NAND2_X1 U591 ( .A1(n543), .A2(n527), .ZN(n529) );
  NOR2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n530), .B(KEYINPUT114), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n539), .A2(n555), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U597 ( .A1(n557), .A2(n539), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XNOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n537) );
  INV_X1 U600 ( .A(n539), .ZN(n534) );
  NOR2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n541) );
  NAND2_X1 U605 ( .A1(n562), .A2(n539), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U608 ( .A1(n543), .A2(n569), .ZN(n544) );
  NOR2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n552), .A2(n571), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  NAND2_X1 U613 ( .A1(n552), .A2(n557), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U616 ( .A(G155GAT), .B(KEYINPUT117), .Z(n551) );
  NAND2_X1 U617 ( .A1(n552), .A2(n578), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n562), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT118), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n563), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U625 ( .A1(n563), .A2(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT56), .Z(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(KEYINPUT60), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT59), .B(n567), .Z(n573) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT123), .ZN(n583) );
  NAND2_X1 U637 ( .A1(n583), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U640 ( .A(n574), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n583), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n580) );
  NAND2_X1 U644 ( .A1(n583), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n585) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

