//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT91), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT11), .B(G169gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  OR3_X1    g006(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT92), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT93), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  OAI22_X1  g015(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n212), .A2(KEYINPUT92), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(KEYINPUT92), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT93), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n208), .B(new_n211), .C1(new_n217), .C2(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n210), .A2(KEYINPUT94), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(new_n208), .ZN(new_n223));
  INV_X1    g022(.A(new_n209), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n224), .A2(new_n225), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n210), .A2(KEYINPUT94), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n222), .A2(new_n223), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT17), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT16), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(G1gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G1gat), .B2(new_n231), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(G8gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n229), .A2(new_n235), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n237), .A2(KEYINPUT18), .A3(new_n240), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n229), .B(new_n235), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n239), .B(KEYINPUT13), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n207), .B1(new_n244), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT96), .ZN(new_n251));
  INV_X1    g050(.A(new_n207), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n243), .A2(new_n245), .A3(new_n248), .A4(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(KEYINPUT96), .B(new_n207), .C1(new_n244), .C2(new_n249), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n257), .A2(KEYINPUT72), .ZN(new_n258));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259));
  INV_X1    g058(.A(G211gat), .ZN(new_n260));
  INV_X1    g059(.A(G218gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n259), .B1(KEYINPUT22), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n258), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(KEYINPUT73), .Z(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT25), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT24), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(G183gat), .A3(G190gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G183gat), .B(G190gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n270), .B1(new_n271), .B2(new_n269), .ZN(new_n272));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT23), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(G169gat), .B2(G176gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n268), .B1(new_n272), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(KEYINPUT64), .B(new_n268), .C1(new_n272), .C2(new_n278), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n268), .B1(new_n273), .B2(KEYINPUT23), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(G169gat), .A3(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n275), .A2(KEYINPUT65), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n283), .A2(new_n285), .A3(new_n277), .A4(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT66), .B1(new_n287), .B2(new_n272), .ZN(new_n288));
  INV_X1    g087(.A(new_n270), .ZN(new_n289));
  XOR2_X1   g088(.A(G183gat), .B(G190gat), .Z(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(KEYINPUT24), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n286), .A2(new_n277), .A3(new_n285), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n283), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n281), .A2(new_n282), .A3(new_n288), .A4(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296));
  NOR3_X1   g095(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT26), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n275), .B1(new_n273), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT27), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G183gat), .ZN(new_n301));
  INV_X1    g100(.A(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT27), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT67), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT67), .ZN(new_n306));
  AOI21_X1  g105(.A(G190gat), .B1(new_n301), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT28), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT28), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n304), .A2(new_n309), .A3(G190gat), .ZN(new_n310));
  OAI221_X1 g109(.A(new_n296), .B1(new_n297), .B2(new_n299), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n267), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n266), .B1(new_n295), .B2(new_n311), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n264), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n312), .A2(new_n267), .ZN(new_n317));
  INV_X1    g116(.A(new_n264), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT29), .B1(new_n295), .B2(new_n311), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n267), .ZN(new_n320));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G64gat), .B(G92gat), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n321), .B(new_n322), .Z(new_n323));
  NAND4_X1  g122(.A1(new_n316), .A2(KEYINPUT30), .A3(new_n320), .A4(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n324), .A2(KEYINPUT75), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n316), .A2(new_n323), .A3(new_n320), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n323), .B(KEYINPUT74), .Z(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(new_n316), .B2(new_n320), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT30), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n324), .A2(KEYINPUT75), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT29), .B1(new_n263), .B2(new_n257), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n257), .B2(new_n263), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n335), .A2(KEYINPUT82), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(KEYINPUT82), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n340));
  INV_X1    g139(.A(G141gat), .ZN(new_n341));
  INV_X1    g140(.A(G148gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344));
  AND2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n343), .B(new_n344), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(G162gat), .ZN(new_n349));
  INV_X1    g148(.A(G162gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(KEYINPUT77), .ZN(new_n351));
  OAI21_X1  g150(.A(G155gat), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n347), .B1(new_n352), .B2(KEYINPUT2), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n345), .B2(new_n346), .ZN(new_n355));
  INV_X1    g154(.A(G155gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n350), .ZN(new_n357));
  NAND2_X1  g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(KEYINPUT76), .A3(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(G141gat), .A2(G148gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(KEYINPUT2), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n355), .A2(new_n359), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n340), .B1(new_n353), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n357), .A2(new_n358), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n350), .A2(KEYINPUT77), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n348), .A2(G162gat), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n356), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT2), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n362), .B(new_n366), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n363), .A2(new_n343), .A3(new_n344), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n345), .A2(new_n346), .A3(new_n354), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT76), .B1(new_n357), .B2(new_n358), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n375), .A3(KEYINPUT79), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n365), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n339), .A2(new_n377), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n353), .A2(new_n364), .A3(KEYINPUT3), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n264), .B1(new_n379), .B2(KEYINPUT29), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G228gat), .ZN(new_n382));
  INV_X1    g181(.A(G233gat), .ZN(new_n383));
  OAI22_X1  g182(.A1(new_n378), .A2(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n337), .B1(new_n371), .B2(new_n375), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n264), .A2(KEYINPUT29), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n353), .A2(new_n364), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n389), .A2(KEYINPUT83), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n382), .A2(new_n383), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(KEYINPUT83), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n390), .A2(new_n391), .A3(new_n380), .A4(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G22gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT31), .B(G50gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  MUX2_X1   g197(.A(G22gat), .B(new_n395), .S(new_n398), .Z(new_n399));
  AND3_X1   g198(.A1(new_n384), .A2(new_n393), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n384), .B2(new_n393), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT90), .B(KEYINPUT35), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n333), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT0), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT85), .ZN(new_n410));
  XOR2_X1   g209(.A(G127gat), .B(G134gat), .Z(new_n411));
  INV_X1    g210(.A(G113gat), .ZN(new_n412));
  INV_X1    g211(.A(G120gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G113gat), .A2(G120gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n411), .A2(new_n416), .A3(KEYINPUT1), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(G113gat), .A2(G120gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(G113gat), .A2(G120gat), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT68), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT68), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n414), .A2(new_n422), .A3(new_n415), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT1), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n425), .A2(KEYINPUT69), .A3(new_n411), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT69), .B1(new_n425), .B2(new_n411), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n418), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(new_n387), .ZN(new_n429));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT5), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n425), .A2(new_n411), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT69), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n425), .A2(KEYINPUT69), .A3(new_n411), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n417), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT3), .B1(new_n353), .B2(new_n364), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n371), .A2(new_n375), .A3(new_n337), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT78), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n436), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n379), .A2(new_n385), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT78), .B1(new_n442), .B2(new_n428), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n430), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT4), .B1(new_n428), .B2(new_n377), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT4), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n436), .A2(new_n446), .A3(new_n387), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT80), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n430), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n440), .B1(new_n436), .B2(new_n439), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n428), .A2(KEYINPUT78), .A3(new_n438), .A4(new_n437), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n445), .A2(new_n447), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n431), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT5), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n436), .A2(new_n446), .A3(new_n365), .A4(new_n376), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT4), .B1(new_n428), .B2(new_n388), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n453), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n410), .B1(new_n457), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n431), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n454), .B1(new_n453), .B2(new_n455), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n409), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT6), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n469), .B1(new_n468), .B2(new_n462), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n464), .A2(new_n472), .B1(new_n473), .B2(KEYINPUT6), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT34), .ZN(new_n476));
  NAND2_X1  g275(.A1(G227gat), .A2(G233gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n295), .A2(new_n311), .A3(new_n428), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n428), .B1(new_n295), .B2(new_n311), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n476), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n312), .A2(new_n436), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n478), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n476), .B1(new_n484), .B2(new_n477), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n483), .A2(G227gat), .A3(G233gat), .A4(new_n478), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT32), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT33), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g289(.A(G15gat), .B(G43gat), .Z(new_n491));
  XNOR2_X1  g290(.A(G71gat), .B(G99gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n488), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n493), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n487), .B(KEYINPUT32), .C1(new_n489), .C2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n486), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n486), .B1(new_n494), .B2(new_n496), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(KEYINPUT89), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n405), .A2(new_n475), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(KEYINPUT6), .B(new_n409), .C1(new_n457), .C2(new_n463), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n457), .B2(new_n470), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n504), .B1(new_n506), .B2(new_n473), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT81), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n331), .A2(new_n332), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n508), .B1(new_n507), .B2(new_n509), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n512));
  INV_X1    g311(.A(new_n486), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT70), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT70), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n515), .A2(new_n517), .A3(new_n402), .A4(new_n497), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n510), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT35), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n503), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n316), .A2(new_n522), .A3(new_n320), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT87), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n316), .A2(KEYINPUT87), .A3(new_n320), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n522), .B1(new_n316), .B2(new_n320), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(new_n323), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT38), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT88), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(KEYINPUT88), .A3(KEYINPUT38), .ZN(new_n534));
  INV_X1    g333(.A(new_n326), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n528), .A2(KEYINPUT38), .A3(new_n327), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n527), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n533), .A2(new_n474), .A3(new_n534), .A4(new_n537), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n331), .A2(new_n464), .A3(new_n332), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n459), .A2(new_n460), .B1(new_n451), .B2(new_n452), .ZN(new_n540));
  OR3_X1    g339(.A1(new_n540), .A2(KEYINPUT39), .A3(new_n430), .ZN(new_n541));
  INV_X1    g340(.A(new_n410), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n429), .A2(new_n430), .ZN(new_n543));
  OAI211_X1 g342(.A(KEYINPUT39), .B(new_n543), .C1(new_n540), .C2(new_n430), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT86), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT40), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT40), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n403), .B1(new_n539), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n538), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n403), .B1(new_n510), .B2(new_n511), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n497), .A2(KEYINPUT36), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n515), .A2(new_n555), .A3(new_n517), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT71), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n500), .A2(KEYINPUT36), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT71), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n515), .A2(new_n555), .A3(new_n559), .A4(new_n517), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n553), .A2(new_n554), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n256), .B1(new_n521), .B2(new_n562), .ZN(new_n563));
  AND3_X1   g362(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT7), .ZN(new_n566));
  INV_X1    g365(.A(G99gat), .ZN(new_n567));
  INV_X1    g366(.A(G106gat), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT8), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT104), .B(G85gat), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n566), .B(new_n569), .C1(G92gat), .C2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n564), .B1(new_n229), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n229), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT105), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n573), .B(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n574), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G190gat), .B(G218gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT103), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n574), .B(new_n580), .C1(new_n576), .C2(new_n578), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT106), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT102), .Z(new_n589));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n582), .A2(KEYINPUT106), .A3(new_n584), .ZN(new_n593));
  INV_X1    g392(.A(new_n591), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n592), .B1(new_n587), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G57gat), .B(G64gat), .ZN(new_n601));
  OAI22_X1  g400(.A1(new_n601), .A2(KEYINPUT97), .B1(KEYINPUT9), .B2(new_n598), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n601), .A2(KEYINPUT97), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT99), .ZN(new_n606));
  INV_X1    g405(.A(new_n600), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G57gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(KEYINPUT98), .A3(G64gat), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n606), .A2(new_n607), .A3(new_n609), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n236), .B1(new_n614), .B2(new_n613), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT100), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G183gat), .B(G211gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT101), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n623), .B(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n619), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n613), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n573), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n573), .A2(new_n633), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n573), .A2(new_n633), .A3(KEYINPUT10), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n632), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n634), .A2(new_n636), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n632), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n640), .A2(new_n642), .A3(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n597), .A2(new_n630), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n563), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n507), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  AND3_X1   g455(.A1(new_n652), .A2(new_n333), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(G8gat), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n652), .B2(new_n333), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT42), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(KEYINPUT42), .B2(new_n657), .ZN(G1325gat));
  INV_X1    g460(.A(G15gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n501), .A2(new_n502), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n652), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n561), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n652), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n667), .B2(new_n662), .ZN(G1326gat));
  NAND3_X1  g467(.A1(new_n563), .A2(new_n403), .A3(new_n651), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(new_n256), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n650), .A2(new_n629), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n521), .A2(new_n562), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n597), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT44), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n596), .B1(new_n521), .B2(new_n562), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n674), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n653), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n681), .A2(KEYINPUT109), .A3(new_n653), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(G29gat), .A3(new_n685), .ZN(new_n686));
  AOI211_X1 g485(.A(new_n596), .B(new_n674), .C1(new_n521), .C2(new_n562), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n215), .A3(new_n653), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(KEYINPUT107), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(KEYINPUT107), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(KEYINPUT45), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n686), .A2(new_n691), .A3(new_n694), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n687), .A2(new_n216), .A3(new_n333), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT46), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n216), .B1(new_n681), .B2(new_n333), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n697), .A2(new_n698), .ZN(G1329gat));
  INV_X1    g498(.A(new_n674), .ZN(new_n700));
  INV_X1    g499(.A(G43gat), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n561), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n675), .B2(new_n597), .ZN(new_n704));
  INV_X1    g503(.A(new_n679), .ZN(new_n705));
  AOI211_X1 g504(.A(new_n596), .B(new_n705), .C1(new_n521), .C2(new_n562), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n700), .B(new_n702), .C1(new_n704), .C2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n687), .A2(new_n664), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n701), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n710), .A2(KEYINPUT111), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n707), .A2(new_n709), .ZN(new_n714));
  INV_X1    g513(.A(new_n711), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n710), .A2(KEYINPUT47), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n712), .B1(new_n716), .B2(new_n717), .ZN(G1330gat));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n403), .B(new_n700), .C1(new_n704), .C2(new_n706), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(G50gat), .ZN(new_n721));
  NOR4_X1   g520(.A1(new_n596), .A2(G50gat), .A3(new_n629), .A4(new_n650), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n563), .A2(new_n403), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n720), .B2(G50gat), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT48), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n721), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI221_X4 g525(.A(new_n723), .B1(new_n719), .B2(KEYINPUT48), .C1(new_n720), .C2(G50gat), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(G1331gat));
  NAND4_X1  g527(.A1(new_n596), .A2(new_n256), .A3(new_n629), .A4(new_n650), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT113), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n562), .B2(new_n521), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n507), .B(KEYINPUT114), .Z(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n333), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT49), .B(G64gat), .Z(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n736), .B2(new_n738), .ZN(G1333gat));
  NAND2_X1  g538(.A1(new_n731), .A2(new_n666), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n663), .A2(G71gat), .ZN(new_n741));
  AOI22_X1  g540(.A1(new_n740), .A2(G71gat), .B1(new_n731), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n742), .B(new_n743), .Z(G1334gat));
  NAND2_X1  g543(.A1(new_n731), .A2(new_n403), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n672), .A2(new_n629), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT51), .B1(new_n676), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n678), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n749), .A2(new_n650), .A3(new_n751), .ZN(new_n752));
  OR3_X1    g551(.A1(new_n752), .A2(new_n507), .A3(new_n570), .ZN(new_n753));
  INV_X1    g552(.A(new_n650), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n677), .B2(new_n680), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n653), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT116), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n570), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n758), .A2(KEYINPUT116), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n753), .B1(new_n760), .B2(new_n761), .ZN(G1336gat));
  INV_X1    g561(.A(G92gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n333), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n752), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n757), .A2(new_n333), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G92gat), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n763), .B1(new_n757), .B2(new_n333), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT52), .B1(new_n765), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(G1337gat));
  NAND2_X1  g572(.A1(new_n664), .A2(new_n567), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n752), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n757), .A2(new_n666), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G99gat), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n567), .B1(new_n757), .B2(new_n666), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT117), .B1(new_n775), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1338gat));
  OAI211_X1 g582(.A(new_n403), .B(new_n755), .C1(new_n704), .C2(new_n706), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n784), .A2(G106gat), .B1(KEYINPUT118), .B2(KEYINPUT53), .ZN(new_n785));
  OR2_X1    g584(.A1(KEYINPUT118), .A2(KEYINPUT53), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n402), .A2(G106gat), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n749), .A2(new_n650), .A3(new_n751), .A4(new_n787), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n786), .B1(new_n785), .B2(new_n788), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(G1339gat));
  AOI21_X1  g590(.A(new_n239), .B1(new_n237), .B2(new_n238), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n246), .A2(new_n247), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n206), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n650), .A2(new_n253), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n637), .A2(new_n638), .A3(new_n632), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n640), .A2(KEYINPUT54), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n647), .B1(new_n640), .B2(KEYINPUT54), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  OR3_X1    g598(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n797), .B2(new_n798), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n649), .A3(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n596), .B(new_n795), .C1(new_n256), .C2(new_n802), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n587), .A2(new_n595), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n253), .A2(new_n794), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n592), .B(new_n804), .C1(new_n802), .C2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n630), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n596), .A2(new_n256), .A3(new_n629), .A4(new_n754), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT119), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n811), .A3(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n333), .A2(new_n507), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n813), .A2(new_n402), .A3(new_n664), .A4(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n815), .A2(new_n412), .A3(new_n256), .ZN(new_n816));
  INV_X1    g615(.A(new_n518), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n813), .A2(new_n817), .A3(new_n733), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n333), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n672), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n816), .B1(new_n820), .B2(new_n412), .ZN(G1340gat));
  NOR3_X1   g620(.A1(new_n815), .A2(new_n413), .A3(new_n754), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n650), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n413), .ZN(G1341gat));
  INV_X1    g623(.A(G127gat), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n819), .A2(new_n825), .A3(new_n629), .ZN(new_n826));
  OAI21_X1  g625(.A(G127gat), .B1(new_n815), .B2(new_n630), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1342gat));
  OR3_X1    g627(.A1(new_n596), .A2(G134gat), .A3(new_n333), .ZN(new_n829));
  OR3_X1    g628(.A1(new_n818), .A2(KEYINPUT56), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G134gat), .B1(new_n815), .B2(new_n596), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT56), .B1(new_n818), .B2(new_n829), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(G1343gat));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n807), .A2(new_n811), .A3(new_n808), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n811), .B1(new_n807), .B2(new_n808), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n733), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n666), .A2(new_n402), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n509), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n341), .A3(new_n672), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n834), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n561), .A2(new_n814), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n403), .B1(new_n835), .B2(new_n836), .ZN(new_n846));
  XNOR2_X1  g645(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n807), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n808), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n807), .A2(new_n849), .ZN(new_n852));
  OAI211_X1 g651(.A(KEYINPUT57), .B(new_n403), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n845), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n341), .B1(new_n854), .B2(new_n672), .ZN(new_n855));
  NOR4_X1   g654(.A1(new_n837), .A2(G141gat), .A3(new_n256), .A4(new_n839), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n843), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT58), .B1(new_n856), .B2(KEYINPUT122), .ZN(new_n858));
  AOI211_X1 g657(.A(new_n256), .B(new_n845), .C1(new_n848), .C2(new_n853), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n858), .B(new_n841), .C1(new_n859), .C2(new_n341), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n860), .ZN(G1344gat));
  NAND3_X1  g660(.A1(new_n840), .A2(new_n342), .A3(new_n650), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  INV_X1    g662(.A(new_n847), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n403), .B(new_n864), .C1(new_n835), .C2(new_n836), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n402), .B1(new_n807), .B2(new_n808), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(KEYINPUT57), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n844), .A2(new_n650), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT123), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n865), .B2(new_n867), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n342), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n863), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n863), .A2(G148gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n854), .B2(new_n650), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n862), .B1(new_n874), .B2(new_n876), .ZN(G1345gat));
  NAND3_X1  g676(.A1(new_n840), .A2(new_n356), .A3(new_n629), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n854), .A2(new_n629), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n356), .ZN(G1346gat));
  NOR2_X1   g679(.A1(new_n349), .A2(new_n351), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n840), .A2(new_n881), .A3(new_n597), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n854), .A2(new_n883), .A3(new_n597), .ZN(new_n884));
  INV_X1    g683(.A(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n883), .B1(new_n854), .B2(new_n597), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(G1347gat));
  NOR3_X1   g687(.A1(new_n733), .A2(new_n509), .A3(new_n663), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n813), .A2(new_n402), .A3(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(G169gat), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n890), .A2(new_n891), .A3(new_n256), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n653), .A2(new_n509), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n817), .B(new_n893), .C1(new_n835), .C2(new_n836), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(G169gat), .B1(new_n895), .B2(new_n672), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n892), .A2(new_n896), .ZN(G1348gat));
  OAI21_X1  g696(.A(G176gat), .B1(new_n890), .B2(new_n754), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n754), .A2(G176gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT125), .ZN(G1349gat));
  NAND4_X1  g700(.A1(new_n813), .A2(new_n402), .A3(new_n629), .A4(new_n889), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G183gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n630), .A2(new_n304), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT126), .B1(new_n894), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n893), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n907), .B1(new_n810), .B2(new_n812), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n817), .A4(new_n904), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n903), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n912));
  OR2_X1    g711(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n911), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(G1350gat));
  OR3_X1    g715(.A1(new_n894), .A2(G190gat), .A3(new_n596), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n890), .A2(new_n596), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n918), .A2(new_n919), .A3(G190gat), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n918), .B2(G190gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(G1351gat));
  AND2_X1   g721(.A1(new_n908), .A2(new_n838), .ZN(new_n923));
  AOI21_X1  g722(.A(G197gat), .B1(new_n923), .B2(new_n672), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n561), .A2(new_n732), .A3(new_n333), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n925), .B1(new_n865), .B2(new_n867), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n672), .A2(G197gat), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G1352gat));
  INV_X1    g727(.A(G204gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n923), .A2(new_n929), .A3(new_n650), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  INV_X1    g730(.A(new_n926), .ZN(new_n932));
  OAI21_X1  g731(.A(G204gat), .B1(new_n932), .B2(new_n754), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(G1353gat));
  NAND3_X1  g734(.A1(new_n923), .A2(new_n260), .A3(new_n629), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n260), .B1(new_n926), .B2(new_n629), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n937), .A2(KEYINPUT63), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(KEYINPUT63), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1354gat));
  OAI21_X1  g739(.A(G218gat), .B1(new_n932), .B2(new_n596), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n923), .A2(new_n261), .A3(new_n597), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1355gat));
endmodule


