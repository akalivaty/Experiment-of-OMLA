//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n215));
  XOR2_X1   g0015(.A(new_n214), .B(new_n215), .Z(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n205), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  INV_X1    g0029(.A(new_n201), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  AND2_X1   g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n216), .A2(new_n229), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  XOR2_X1   g0045(.A(G58), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G222), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(G223), .A3(G1698), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G77), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n258), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n264), .A2(KEYINPUT66), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G1), .A3(G13), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(new_n264), .B2(KEYINPUT66), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(new_n267), .A3(G274), .ZN(new_n273));
  INV_X1    g0073(.A(G226), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G179), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n277), .B1(new_n265), .B2(new_n268), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n210), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n282), .A2(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n287), .B1(G20), .B2(new_n203), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G1), .A2(G13), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(new_n290), .A3(new_n289), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n209), .A2(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G50), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n295), .A2(new_n297), .B1(G50), .B2(new_n294), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n281), .A2(G169), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n280), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n288), .A2(new_n292), .ZN(new_n301));
  INV_X1    g0101(.A(new_n298), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(KEYINPUT9), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n293), .B2(new_n298), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n303), .B(new_n305), .C1(new_n306), .C2(new_n281), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n281), .A2(G190), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT10), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n303), .A2(new_n305), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n279), .A2(G200), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n308), .A4(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n300), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n296), .A2(G77), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n295), .A2(new_n317), .B1(G77), .B2(new_n294), .ZN(new_n318));
  XOR2_X1   g0118(.A(KEYINPUT8), .B(G58), .Z(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT15), .B(G87), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n283), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n318), .B1(new_n322), .B2(new_n291), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n225), .A2(new_n257), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n219), .A2(G1698), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n262), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n290), .B1(G33), .B2(G41), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n256), .B2(G107), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G244), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n273), .B1(new_n331), .B2(new_n276), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n324), .B(KEYINPUT67), .C1(G169), .C2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT67), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n333), .A2(G169), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n323), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n333), .A2(G190), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n323), .C1(new_n306), .C2(new_n333), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT16), .ZN(new_n344));
  INV_X1    g0144(.A(G159), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n286), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT71), .ZN(new_n348));
  XNOR2_X1  g0148(.A(G58), .B(G68), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(G20), .ZN(new_n350));
  AND2_X1   g0150(.A1(G58), .A2(G68), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n348), .B(G20), .C1(new_n351), .C2(new_n201), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n347), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n254), .A2(new_n210), .A3(new_n255), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n255), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n218), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n344), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT7), .B1(new_n262), .B2(new_n210), .ZN(new_n361));
  INV_X1    g0161(.A(new_n358), .ZN(new_n362));
  OAI21_X1  g0162(.A(G68), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n351), .B2(new_n201), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT71), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n346), .B1(new_n365), .B2(new_n352), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n366), .A3(KEYINPUT16), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n360), .A2(new_n291), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n319), .A2(new_n296), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n369), .A2(new_n295), .B1(new_n319), .B2(new_n294), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT72), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n267), .A2(G232), .A3(new_n275), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n273), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(G223), .B(new_n257), .C1(new_n260), .C2(new_n261), .ZN(new_n376));
  OAI211_X1 g0176(.A(G226), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n375), .B1(new_n328), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G169), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(G179), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n372), .A2(new_n373), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n373), .B1(new_n372), .B2(new_n384), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n379), .A2(new_n328), .ZN(new_n389));
  INV_X1    g0189(.A(G190), .ZN(new_n390));
  INV_X1    g0190(.A(new_n375), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(G200), .B2(new_n380), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n368), .A2(new_n371), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT17), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n343), .A2(new_n388), .A3(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n285), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n397));
  INV_X1    g0197(.A(G77), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(new_n283), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n291), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT11), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n294), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n218), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT12), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n399), .A2(KEYINPUT11), .A3(new_n291), .ZN(new_n406));
  INV_X1    g0206(.A(new_n295), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(G68), .A3(new_n296), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n402), .A2(new_n405), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n274), .A2(new_n257), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n225), .A2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n260), .C2(new_n261), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n253), .A2(new_n205), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n328), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n267), .A2(G238), .A3(new_n275), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n273), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT13), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n267), .B1(new_n412), .B2(new_n414), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n273), .A2(new_n417), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT13), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n409), .B1(G200), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n416), .A2(new_n418), .A3(KEYINPUT68), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT68), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n421), .B2(new_n422), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(KEYINPUT13), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(G190), .A3(new_n420), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n424), .A2(G169), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT69), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT14), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(KEYINPUT14), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n424), .A2(G169), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n421), .A2(new_n422), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n338), .B1(new_n438), .B2(new_n419), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n429), .A2(KEYINPUT70), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT70), .B1(new_n429), .B2(new_n439), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n435), .B(new_n437), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n409), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NOR4_X1   g0244(.A1(new_n316), .A2(new_n396), .A3(new_n432), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G116), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G20), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT23), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n210), .B2(G107), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n210), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n452), .A2(KEYINPUT22), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(KEYINPUT22), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT24), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT24), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(new_n451), .C1(new_n453), .C2(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n291), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n271), .A2(G1), .ZN(new_n461));
  AND2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  NOR2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G264), .A3(new_n267), .ZN(new_n465));
  INV_X1    g0265(.A(G274), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n232), .B2(new_n266), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT5), .B(G41), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(new_n461), .ZN(new_n469));
  NOR2_X1   g0269(.A1(G250), .A2(G1698), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n226), .B2(G1698), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT75), .B(G294), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n471), .A2(new_n256), .B1(new_n472), .B2(G33), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n465), .B(new_n469), .C1(new_n473), .C2(new_n267), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n306), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(G190), .B2(new_n474), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n295), .B1(new_n209), .B2(G33), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT25), .B1(new_n403), .B2(new_n206), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n403), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n477), .A2(G107), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n460), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  XOR2_X1   g0282(.A(KEYINPUT75), .B(G294), .Z(new_n483));
  NAND2_X1  g0283(.A1(new_n226), .A2(G1698), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(G250), .B2(G1698), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n483), .A2(new_n253), .B1(new_n485), .B2(new_n262), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n468), .A2(new_n461), .B1(new_n232), .B2(new_n266), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n486), .A2(new_n328), .B1(new_n487), .B2(G264), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n338), .A3(new_n469), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n474), .A2(new_n381), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n292), .B1(new_n456), .B2(new_n458), .ZN(new_n491));
  INV_X1    g0291(.A(new_n481), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n489), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n482), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G244), .B(new_n257), .C1(new_n260), .C2(new_n261), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n257), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n328), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n464), .A2(new_n267), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n469), .B1(new_n503), .B2(new_n226), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(new_n390), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n504), .B1(new_n501), .B2(new_n328), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(G200), .B2(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n509));
  XNOR2_X1  g0309(.A(G97), .B(G107), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT6), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n512), .A2(new_n210), .B1(new_n398), .B2(new_n286), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n206), .B1(new_n357), .B2(new_n358), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n291), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n294), .A2(G97), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n477), .B2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n508), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n219), .A2(new_n257), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n331), .A2(G1698), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n260), .C2(new_n261), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n446), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n328), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n221), .B1(new_n209), .B2(G45), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n467), .A2(new_n461), .B1(new_n267), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(G190), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n267), .B1(new_n523), .B2(new_n446), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n267), .A2(G274), .A3(new_n461), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n526), .A2(new_n267), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(G200), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n207), .A2(G87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(KEYINPUT73), .A2(KEYINPUT19), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(KEYINPUT73), .A2(KEYINPUT19), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n413), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n536), .B1(new_n540), .B2(new_n210), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n210), .B(G68), .C1(new_n260), .C2(new_n261), .ZN(new_n542));
  INV_X1    g0342(.A(new_n539), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n537), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n283), .A2(new_n205), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n291), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n321), .A2(new_n403), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n477), .A2(G87), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n321), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n477), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n547), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n525), .A2(G179), .A3(new_n527), .ZN(new_n555));
  OAI21_X1  g0355(.A(G169), .B1(new_n529), .B2(new_n532), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n535), .A2(new_n551), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n502), .A2(new_n505), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n381), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n502), .A2(new_n338), .A3(new_n505), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n518), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n520), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G264), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n564));
  OAI211_X1 g0364(.A(G257), .B(new_n257), .C1(new_n260), .C2(new_n261), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n254), .A2(G303), .A3(new_n255), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n567), .A2(new_n328), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n464), .A2(G270), .A3(new_n267), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n469), .ZN(new_n570));
  OAI211_X1 g0370(.A(KEYINPUT21), .B(G169), .C1(new_n568), .C2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n569), .A2(new_n469), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n328), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(G179), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n499), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT74), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT20), .ZN(new_n578));
  INV_X1    g0378(.A(G116), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n577), .A2(new_n578), .B1(new_n579), .B2(G20), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n576), .A2(new_n580), .A3(new_n291), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(KEYINPUT74), .A3(KEYINPUT20), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n209), .A2(G33), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n407), .A2(G116), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n403), .A2(new_n579), .ZN(new_n585));
  NAND2_X1  g0385(.A1(KEYINPUT74), .A2(KEYINPUT20), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n576), .A2(new_n580), .A3(new_n291), .A4(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n582), .A2(new_n584), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n575), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n306), .B1(new_n572), .B2(new_n573), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n588), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n572), .A2(new_n573), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n591), .B(new_n592), .C1(new_n390), .C2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n381), .B1(new_n572), .B2(new_n573), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n588), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n589), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n563), .A2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n445), .A2(new_n494), .A3(new_n600), .ZN(G372));
  INV_X1    g0401(.A(new_n310), .ZN(new_n602));
  INV_X1    g0402(.A(new_n314), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n432), .A2(new_n340), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n395), .B1(new_n444), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n604), .B1(new_n606), .B2(new_n388), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT79), .B1(new_n607), .B2(new_n300), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT79), .ZN(new_n609));
  INV_X1    g0409(.A(new_n388), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n443), .B1(new_n432), .B2(new_n340), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n610), .B1(new_n611), .B2(new_n395), .ZN(new_n612));
  OAI221_X1 g0412(.A(new_n609), .B1(new_n280), .B2(new_n299), .C1(new_n612), .C2(new_n604), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n534), .A2(new_n550), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT76), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n381), .B1(new_n525), .B2(new_n527), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n529), .A2(new_n532), .A3(new_n338), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n555), .A2(KEYINPUT76), .A3(new_n556), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n615), .B1(new_n621), .B2(new_n554), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT78), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n518), .A2(new_n561), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n507), .A2(G169), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT26), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n338), .A2(new_n507), .B1(new_n515), .B2(new_n517), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(KEYINPUT78), .A3(new_n560), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n622), .A2(new_n626), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n535), .A2(new_n551), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n557), .A2(new_n554), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n631), .A2(new_n628), .A3(new_n632), .A4(new_n560), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n633), .A2(KEYINPUT26), .B1(new_n554), .B2(new_n621), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n489), .A2(new_n490), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n460), .B2(new_n481), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n570), .B1(new_n328), .B2(new_n567), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n595), .A2(KEYINPUT21), .B1(new_n637), .B2(G179), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n598), .B(KEYINPUT77), .C1(new_n638), .C2(new_n592), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT77), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n592), .B1(new_n571), .B2(new_n574), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT21), .B1(new_n595), .B2(new_n588), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n636), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n622), .A2(new_n482), .A3(new_n562), .A4(new_n520), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n630), .B(new_n634), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n445), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n614), .A2(new_n647), .ZN(G369));
  NOR3_X1   g0448(.A1(new_n568), .A2(new_n390), .A3(new_n570), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n649), .A2(new_n590), .A3(new_n588), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n650), .A2(new_n641), .A3(new_n642), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n588), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n639), .A2(new_n643), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n658), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n657), .B1(new_n491), .B2(new_n492), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n494), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n636), .A2(new_n657), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n657), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n636), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n482), .A2(new_n493), .A3(new_n669), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n589), .A2(new_n598), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n668), .A2(new_n670), .A3(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n213), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n536), .A2(new_n579), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n677), .A2(G1), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n231), .B2(new_n677), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n646), .A2(new_n669), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(KEYINPUT29), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n624), .A2(new_n625), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n686), .A2(new_n627), .A3(new_n558), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n621), .A2(new_n554), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n622), .A2(new_n626), .A3(new_n629), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT26), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n672), .A2(new_n636), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n689), .B(new_n691), .C1(new_n645), .C2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n685), .B1(new_n693), .B2(new_n669), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n684), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G330), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n465), .B1(new_n473), .B2(new_n267), .ZN(new_n697));
  NOR2_X1   g0497(.A1(G238), .A2(G1698), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n331), .B2(G1698), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n699), .A2(new_n256), .B1(G33), .B2(G116), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n527), .B1(new_n700), .B2(new_n267), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT80), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT80), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n529), .A2(new_n532), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n488), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n507), .A2(KEYINPUT30), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n572), .A2(G179), .A3(new_n573), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n706), .A2(new_n708), .A3(KEYINPUT81), .A4(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n702), .A2(new_n709), .A3(new_n705), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(new_n559), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT81), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n712), .B2(new_n707), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n704), .A2(G179), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n559), .A2(new_n474), .A3(new_n593), .A4(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n710), .A2(new_n713), .A3(new_n715), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n657), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT31), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n721), .A3(new_n657), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n519), .A2(new_n508), .B1(new_n628), .B2(new_n560), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n651), .A2(new_n724), .A3(new_n558), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n482), .A2(new_n493), .A3(new_n669), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT82), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n520), .A2(new_n558), .A3(new_n562), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT82), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n671), .A2(new_n728), .A3(new_n729), .A4(new_n651), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n696), .B1(new_n723), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n695), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n682), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(G13), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n735), .A2(new_n271), .A3(G20), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT83), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n676), .A2(new_n737), .A3(new_n209), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n663), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(G330), .B2(new_n661), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n213), .A2(new_n256), .ZN(new_n741));
  INV_X1    g0541(.A(G355), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n741), .A2(new_n742), .B1(G116), .B2(new_n213), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n247), .A2(G45), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n675), .A2(new_n256), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n231), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(new_n271), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n743), .B1(new_n744), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n735), .A2(new_n253), .A3(KEYINPUT84), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT84), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G13), .B2(G33), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n290), .B1(G20), .B2(new_n381), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n738), .B1(new_n749), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(G20), .A2(G179), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT85), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n390), .A2(G200), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G322), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n762), .A2(new_n390), .A3(G200), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT33), .B(G317), .Z(new_n767));
  OAI21_X1  g0567(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT89), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n210), .A2(G179), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n256), .B1(new_n773), .B2(G329), .ZN(new_n774));
  INV_X1    g0574(.A(G283), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n770), .A2(new_n390), .A3(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n763), .A2(new_n338), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n774), .B1(new_n775), .B2(new_n776), .C1(new_n483), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n762), .A2(new_n771), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n780), .B1(G311), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT88), .Z(new_n785));
  AND3_X1   g0585(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n785), .A2(G303), .B1(G326), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n769), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n776), .A2(new_n206), .ZN(new_n789));
  INV_X1    g0589(.A(new_n784), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n262), .B(new_n789), .C1(G87), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n772), .A2(new_n345), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT32), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n791), .B(new_n793), .C1(new_n398), .C2(new_n781), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G50), .B2(new_n786), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n764), .B(KEYINPUT86), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n224), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n778), .A2(G97), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n766), .B2(new_n218), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT87), .Z(new_n800));
  OAI21_X1  g0600(.A(new_n788), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n759), .B1(new_n801), .B2(new_n756), .ZN(new_n802));
  INV_X1    g0602(.A(new_n755), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n661), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n740), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  INV_X1    g0606(.A(new_n738), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n753), .A2(new_n756), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n398), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n324), .A2(new_n657), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n340), .A2(new_n342), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n340), .B2(new_n810), .ZN(new_n812));
  INV_X1    g0612(.A(new_n786), .ZN(new_n813));
  INV_X1    g0613(.A(G137), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n813), .A2(new_n814), .B1(new_n781), .B2(new_n345), .ZN(new_n815));
  INV_X1    g0615(.A(new_n766), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(G150), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G143), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n796), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT34), .Z(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n256), .B1(new_n772), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n776), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(G68), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n785), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n224), .B2(new_n779), .C1(new_n825), .C2(new_n202), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n256), .B1(new_n785), .B2(G107), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT90), .ZN(new_n829));
  INV_X1    g0629(.A(G303), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n813), .A2(new_n830), .B1(new_n775), .B2(new_n766), .ZN(new_n831));
  INV_X1    g0631(.A(new_n764), .ZN(new_n832));
  INV_X1    g0632(.A(G294), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n832), .A2(new_n833), .B1(new_n579), .B2(new_n781), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n776), .A2(new_n220), .ZN(new_n835));
  INV_X1    g0635(.A(G311), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n798), .B1(new_n836), .B2(new_n772), .ZN(new_n837));
  NOR4_X1   g0637(.A1(new_n831), .A2(new_n834), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n827), .B1(new_n829), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n756), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n809), .B1(new_n754), .B2(new_n812), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT91), .ZN(new_n842));
  INV_X1    g0642(.A(new_n732), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n340), .A2(new_n810), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n343), .B2(new_n810), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n683), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n646), .A2(new_n669), .A3(new_n812), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n738), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n732), .A2(new_n846), .A3(new_n847), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n842), .A2(new_n851), .ZN(G384));
  INV_X1    g0652(.A(new_n512), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n579), .B(new_n233), .C1(new_n853), .C2(KEYINPUT35), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(KEYINPUT35), .B2(new_n853), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT36), .ZN(new_n856));
  OAI21_X1  g0656(.A(G77), .B1(new_n224), .B2(new_n218), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n231), .A2(new_n857), .B1(G50), .B2(new_n218), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(G1), .A3(new_n735), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT92), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n409), .A2(new_n657), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n443), .A2(new_n431), .A3(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n409), .B(new_n657), .C1(new_n442), .C2(new_n432), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n340), .A2(new_n657), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n865), .B1(new_n847), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n363), .A2(new_n366), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n292), .B1(new_n869), .B2(new_n344), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n370), .B1(new_n870), .B2(new_n367), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n394), .B1(new_n871), .B2(new_n655), .ZN(new_n872));
  INV_X1    g0672(.A(new_n370), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n368), .A2(new_n873), .B1(new_n382), .B2(new_n383), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n372), .A2(new_n384), .ZN(new_n876));
  INV_X1    g0676(.A(new_n655), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n372), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n876), .A2(new_n878), .A3(new_n879), .A4(new_n394), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT93), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT93), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n875), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  INV_X1    g0684(.A(new_n387), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT17), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n394), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n394), .A2(new_n886), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n885), .A2(new_n887), .A3(new_n385), .A4(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n871), .A2(new_n655), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n884), .A4(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n881), .A2(KEYINPUT93), .B1(new_n889), .B2(new_n890), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n894), .B2(new_n884), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n868), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT94), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n388), .A2(new_n877), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n882), .A2(new_n884), .A3(new_n891), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n876), .A2(new_n878), .A3(new_n394), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(new_n879), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n878), .B1(new_n388), .B2(new_n395), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n892), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n443), .A2(new_n657), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n904), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n900), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n897), .B1(new_n896), .B2(new_n899), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n445), .B1(new_n684), .B2(new_n694), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n614), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n918), .B(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT40), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n893), .A2(new_n895), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n729), .B1(new_n600), .B2(new_n671), .ZN(new_n924));
  NOR4_X1   g0724(.A1(new_n726), .A2(new_n563), .A3(new_n599), .A4(KEYINPUT82), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n718), .A2(new_n721), .A3(new_n657), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n721), .B1(new_n718), .B2(new_n657), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n924), .A2(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n845), .B1(new_n863), .B2(new_n864), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n922), .B1(new_n923), .B2(new_n930), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n720), .A2(new_n722), .B1(new_n727), .B2(new_n730), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n863), .A2(new_n864), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n812), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT95), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n922), .B1(new_n892), .B2(new_n908), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT95), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n928), .A2(new_n929), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n931), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n445), .A2(new_n928), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(G330), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n921), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(G1), .B1(new_n735), .B2(G20), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n921), .A2(new_n944), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n861), .B1(new_n947), .B2(new_n948), .ZN(G367));
  NOR2_X1   g0749(.A1(new_n746), .A2(new_n242), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n757), .B1(new_n213), .B2(new_n321), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n813), .A2(new_n836), .B1(new_n483), .B2(new_n766), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT46), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n579), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n952), .B1(new_n785), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n953), .B1(new_n784), .B2(new_n579), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n781), .B2(new_n775), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n823), .A2(G97), .ZN(new_n958));
  INV_X1    g0758(.A(G317), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n958), .B(new_n262), .C1(new_n959), .C2(new_n772), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n957), .B(new_n960), .C1(G107), .C2(new_n778), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n955), .B(new_n961), .C1(new_n830), .C2(new_n796), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n256), .B1(new_n776), .B2(new_n398), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(G68), .B2(new_n778), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n202), .B2(new_n781), .C1(new_n284), .C2(new_n832), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n784), .A2(new_n224), .B1(new_n772), .B2(new_n814), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT103), .Z(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n818), .B2(new_n813), .C1(new_n345), .C2(new_n766), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n962), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT47), .Z(new_n970));
  OAI221_X1 g0770(.A(new_n738), .B1(new_n950), .B2(new_n951), .C1(new_n970), .C2(new_n840), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT104), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n550), .A2(new_n657), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n622), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT96), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n622), .A2(KEYINPUT96), .A3(new_n973), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(new_n688), .C2(new_n973), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT97), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n755), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n972), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n979), .B(KEYINPUT43), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n518), .A2(new_n657), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n724), .A2(new_n983), .B1(new_n686), .B2(new_n657), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT98), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n562), .B1(new_n986), .B2(new_n493), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n669), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n673), .A2(new_n984), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT42), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n982), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n978), .B(KEYINPUT97), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n988), .A2(new_n994), .A3(new_n990), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT99), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n995), .A2(new_n996), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n668), .A2(new_n986), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(KEYINPUT100), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n999), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1003), .A2(new_n997), .A3(new_n1001), .A4(new_n992), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT100), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n998), .A2(new_n999), .B1(new_n668), .B2(new_n986), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1002), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n737), .A2(new_n209), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n673), .A2(new_n670), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n1011), .A2(KEYINPUT101), .A3(new_n984), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT101), .B1(new_n1011), .B2(new_n984), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1011), .A2(new_n984), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT44), .Z(new_n1018));
  NAND3_X1  g0818(.A1(new_n1012), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1016), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1020), .A2(new_n663), .A3(new_n667), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n657), .B1(new_n589), .B2(new_n598), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n673), .B1(new_n667), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(KEYINPUT102), .B2(new_n662), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n662), .B(KEYINPUT102), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n1023), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1016), .A2(new_n1018), .A3(new_n668), .A4(new_n1019), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1021), .A2(new_n733), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n733), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n676), .B(KEYINPUT41), .Z(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1010), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n981), .B1(new_n1008), .B2(new_n1032), .ZN(G387));
  INV_X1    g0833(.A(KEYINPUT109), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT108), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1025), .A2(new_n1023), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1035), .B1(new_n695), .B2(new_n732), .C1(new_n1036), .C2(new_n1024), .ZN(new_n1037));
  OAI21_X1  g0837(.A(KEYINPUT108), .B1(new_n733), .B2(new_n1026), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n733), .A2(new_n1026), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n676), .A4(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n271), .B1(new_n218), .B2(new_n398), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n678), .B2(KEYINPUT105), .ZN(new_n1042));
  AND3_X1   g0842(.A1(new_n319), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT50), .B1(new_n319), .B2(new_n202), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1042), .B1(KEYINPUT105), .B2(new_n678), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n745), .B(new_n1045), .C1(new_n239), .C2(new_n271), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(G107), .B2(new_n213), .C1(new_n679), .C2(new_n741), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n807), .B1(new_n1047), .B2(new_n757), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n813), .A2(new_n345), .B1(new_n282), .B2(new_n766), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n832), .A2(new_n202), .B1(new_n218), .B2(new_n781), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n262), .B1(new_n773), .B2(G150), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n790), .A2(G77), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n778), .A2(new_n552), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1051), .A2(new_n958), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n1049), .A2(new_n1050), .A3(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n766), .A2(new_n836), .B1(new_n781), .B2(new_n830), .ZN(new_n1056));
  XOR2_X1   g0856(.A(KEYINPUT106), .B(G322), .Z(new_n1057));
  AOI21_X1  g0857(.A(new_n1056), .B1(new_n786), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n796), .B2(new_n959), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n472), .A2(new_n790), .B1(new_n778), .B2(G283), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT107), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT49), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n256), .B1(new_n773), .B2(G326), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n579), .B2(new_n776), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1055), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1048), .B1(new_n667), .B2(new_n803), .C1(new_n1071), .C2(new_n840), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1026), .A2(new_n1010), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1034), .B1(new_n1040), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1040), .A2(new_n1034), .A3(new_n1074), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(G393));
  INV_X1    g0878(.A(KEYINPUT110), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1021), .A2(new_n1079), .A3(new_n1027), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1027), .A2(new_n1079), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n985), .A2(new_n803), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT111), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n256), .B(new_n789), .C1(new_n773), .C2(new_n1057), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n775), .B2(new_n784), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G294), .B2(new_n782), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n813), .A2(new_n959), .B1(new_n832), .B2(new_n836), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n1090));
  OAI21_X1  g0890(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n766), .A2(new_n830), .B1(new_n779), .B2(new_n579), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT113), .Z(new_n1094));
  OAI22_X1  g0894(.A1(new_n813), .A2(new_n284), .B1(new_n832), .B2(new_n345), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT51), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n262), .B(new_n835), .C1(G143), .C2(new_n773), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G68), .A2(new_n790), .B1(new_n778), .B2(G77), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n282), .C2(new_n781), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G50), .B2(new_n816), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1092), .A2(new_n1094), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(new_n840), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n745), .A2(new_n250), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n758), .B1(G97), .B2(new_n675), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n807), .B(new_n1102), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1082), .A2(new_n1010), .B1(new_n1084), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1080), .A2(new_n1081), .A3(new_n1039), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1107), .A2(new_n676), .A3(new_n1028), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(G390));
  INV_X1    g0909(.A(new_n808), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n262), .B1(new_n772), .B2(new_n833), .C1(new_n218), .C2(new_n776), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n832), .A2(new_n579), .B1(new_n205), .B2(new_n781), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1111), .B(new_n1112), .C1(G77), .C2(new_n778), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n825), .A2(new_n220), .B1(new_n206), .B2(new_n766), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G283), .B2(new_n786), .ZN(new_n1115));
  INV_X1    g0915(.A(G125), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n256), .B1(new_n772), .B2(new_n1116), .C1(new_n779), .C2(new_n345), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n832), .A2(new_n821), .B1(new_n781), .B2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1117), .B(new_n1119), .C1(G50), .C2(new_n823), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n766), .A2(new_n814), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n790), .A2(G150), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT53), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1121), .B(new_n1123), .C1(G128), .C2(new_n786), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1113), .A2(new_n1115), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n738), .B1(new_n319), .B2(new_n1110), .C1(new_n1125), .C2(new_n840), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n904), .A2(new_n911), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n753), .ZN(new_n1128));
  NOR4_X1   g0928(.A1(new_n932), .A2(new_n696), .A3(new_n865), .A4(new_n845), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n868), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n912), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n904), .A2(new_n911), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n909), .A2(new_n1131), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n933), .B(KEYINPUT114), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n693), .A2(new_n669), .A3(new_n812), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n867), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1133), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1129), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1127), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n732), .A2(new_n812), .A3(new_n933), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1136), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n865), .B(KEYINPUT114), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1131), .B(new_n909), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1140), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1138), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT116), .B1(new_n1146), .B2(new_n1009), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT116), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1138), .A2(new_n1145), .A3(new_n1148), .A4(new_n1010), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1128), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n732), .A2(new_n445), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n614), .A2(new_n919), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n732), .A2(new_n812), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1143), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n847), .A2(new_n867), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n933), .B1(new_n732), .B2(new_n812), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n1129), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1152), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n1138), .A3(new_n1145), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT115), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n1161), .A3(new_n676), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1159), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1146), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1161), .B1(new_n1160), .B2(new_n676), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1150), .B1(new_n1165), .B2(new_n1166), .ZN(G378));
  AOI21_X1  g0967(.A(new_n930), .B1(new_n892), .B2(new_n903), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n939), .B(G330), .C1(new_n1168), .C2(KEYINPUT40), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n655), .B1(new_n301), .B2(new_n302), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n315), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT119), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n315), .A2(new_n1171), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n315), .A2(new_n1171), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT119), .B1(new_n1177), .B2(new_n1172), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g0979(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1176), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1169), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1186), .A2(new_n931), .A3(G330), .A4(new_n939), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n918), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n914), .A2(new_n916), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n1187), .A3(new_n1185), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1009), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n256), .A2(G41), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(G33), .A2(G41), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1193), .A2(G50), .A3(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n786), .A2(G116), .B1(G68), .B2(new_n778), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT117), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n766), .A2(new_n205), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n776), .A2(new_n224), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n773), .A2(G283), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1200), .A2(new_n1052), .A3(new_n1201), .A4(new_n1193), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n832), .A2(new_n206), .B1(new_n321), .B2(new_n781), .ZN(new_n1203));
  NOR4_X1   g1003(.A1(new_n1197), .A2(new_n1198), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1195), .B1(new_n1204), .B2(KEYINPUT58), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n764), .A2(G128), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n284), .B2(new_n779), .C1(new_n784), .C2(new_n1118), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n813), .A2(new_n1116), .B1(new_n821), .B2(new_n766), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(G137), .C2(new_n782), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  INV_X1    g1011(.A(G124), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1194), .B1(new_n772), .B2(new_n1212), .C1(new_n345), .C2(new_n776), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT118), .Z(new_n1214));
  INV_X1    g1014(.A(KEYINPUT59), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1214), .B1(new_n1209), .B2(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1205), .B1(KEYINPUT58), .B2(new_n1204), .C1(new_n1211), .C2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n756), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n807), .B1(new_n202), .B2(new_n808), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n1186), .C2(new_n754), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1192), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1152), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1160), .A2(new_n1223), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1190), .A2(new_n1187), .A3(new_n1185), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1185), .A2(new_n1187), .B1(new_n915), .B2(new_n917), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1224), .B(KEYINPUT57), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n676), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1189), .A2(new_n1191), .B1(new_n1160), .B2(new_n1223), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(KEYINPUT57), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1222), .B1(new_n1228), .B2(new_n1230), .ZN(G375));
  NAND3_X1  g1031(.A1(new_n1155), .A2(new_n1158), .A3(new_n1152), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1163), .A2(new_n1031), .A3(new_n1232), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n262), .B(new_n1199), .C1(G128), .C2(new_n773), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n202), .B2(new_n779), .C1(new_n284), .C2(new_n781), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n786), .A2(G132), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n766), .B2(new_n1118), .C1(new_n825), .C2(new_n345), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n796), .A2(new_n814), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1235), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G116), .A2(new_n816), .B1(new_n786), .B2(G294), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n825), .B2(new_n205), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n778), .A2(new_n552), .B1(new_n773), .B2(G303), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1242), .B1(new_n206), .B2(new_n781), .C1(new_n832), .C2(new_n775), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n262), .B1(new_n776), .B2(new_n398), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT120), .Z(new_n1245));
  NOR3_X1   g1045(.A1(new_n1241), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n756), .B1(new_n1239), .B2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1247), .B(new_n738), .C1(G68), .C2(new_n1110), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1143), .B2(new_n753), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1010), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1233), .A2(new_n1251), .ZN(G381));
  NOR2_X1   g1052(.A1(G375), .A2(G378), .ZN(new_n1253));
  INV_X1    g1053(.A(G387), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1076), .A2(new_n805), .A3(new_n1077), .ZN(new_n1255));
  NOR4_X1   g1055(.A1(new_n1255), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .ZN(G407));
  NAND2_X1  g1057(.A1(new_n656), .A2(G213), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1253), .A2(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(G407), .A2(G213), .A3(new_n1260), .ZN(G409));
  NAND4_X1  g1061(.A1(new_n1155), .A2(new_n1158), .A3(new_n1152), .A4(KEYINPUT60), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT123), .ZN(new_n1263));
  XOR2_X1   g1063(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n1264));
  NAND2_X1  g1064(.A1(new_n1232), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n1163), .A3(new_n676), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1251), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(G384), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G384), .B(new_n1251), .C1(new_n1263), .C2(new_n1266), .ZN(new_n1270));
  AND4_X1   g1070(.A1(G2897), .A2(new_n1269), .A3(new_n1259), .A4(new_n1270), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1269), .A2(new_n1270), .B1(G2897), .B2(new_n1259), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT121), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1192), .B2(new_n1221), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1010), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(KEYINPUT121), .A3(new_n1220), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1229), .A2(new_n1031), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(G378), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G378), .B(new_n1222), .C1(new_n1228), .C2(new_n1230), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1259), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1273), .B1(KEYINPUT124), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT124), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1285), .B1(new_n1286), .B2(new_n1259), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1077), .ZN(new_n1289));
  OAI21_X1  g1089(.A(G396), .B1(new_n1289), .B2(new_n1075), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n1255), .A3(G390), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(G390), .B1(new_n1290), .B2(new_n1255), .ZN(new_n1293));
  OAI21_X1  g1093(.A(G387), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1290), .A2(new_n1255), .ZN(new_n1295));
  INV_X1    g1095(.A(G390), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(new_n1254), .A3(new_n1291), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1294), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1259), .B(new_n1301), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1300), .B1(new_n1302), .B2(KEYINPUT63), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1301), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1283), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT63), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1288), .A2(new_n1303), .A3(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1299), .B1(new_n1283), .B2(new_n1273), .ZN(new_n1309));
  AND2_X1   g1109(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1310), .B1(new_n1302), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1305), .A2(new_n1311), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1309), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  AND2_X1   g1115(.A1(new_n1294), .A2(new_n1298), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1308), .B1(new_n1315), .B2(new_n1316), .ZN(G405));
  AND2_X1   g1117(.A1(G375), .A2(new_n1280), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1282), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT127), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1304), .A2(KEYINPUT126), .A3(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT126), .ZN(new_n1323));
  OAI21_X1  g1123(.A(KEYINPUT127), .B1(new_n1301), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1320), .A2(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1324), .B(new_n1322), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1316), .ZN(G402));
endmodule


