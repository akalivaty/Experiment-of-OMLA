

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588;

  XOR2_X1 U321 ( .A(n411), .B(n410), .Z(n289) );
  OR2_X1 U322 ( .A1(n536), .A2(n522), .ZN(n461) );
  XNOR2_X1 U323 ( .A(KEYINPUT25), .B(KEYINPUT99), .ZN(n463) );
  XNOR2_X1 U324 ( .A(n464), .B(n463), .ZN(n471) );
  XNOR2_X1 U325 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n396) );
  XNOR2_X1 U326 ( .A(n397), .B(n396), .ZN(n530) );
  XNOR2_X1 U327 ( .A(n418), .B(KEYINPUT54), .ZN(n419) );
  XNOR2_X1 U328 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U329 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U330 ( .A(n412), .B(n289), .ZN(n414) );
  XNOR2_X1 U331 ( .A(n384), .B(n383), .ZN(n387) );
  XNOR2_X1 U332 ( .A(n416), .B(n415), .ZN(n522) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U334 ( .A(n484), .B(KEYINPUT108), .ZN(n485) );
  XNOR2_X1 U335 ( .A(n487), .B(G29GAT), .ZN(n488) );
  XNOR2_X1 U336 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XNOR2_X1 U337 ( .A(n486), .B(n485), .ZN(G1331GAT) );
  XOR2_X1 U338 ( .A(G99GAT), .B(G85GAT), .Z(n366) );
  XOR2_X1 U339 ( .A(KEYINPUT65), .B(KEYINPUT77), .Z(n291) );
  XNOR2_X1 U340 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n290) );
  XNOR2_X1 U341 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U342 ( .A(n366), .B(n292), .Z(n298) );
  XOR2_X1 U343 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n294) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(G29GAT), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n296) );
  INV_X1 U346 ( .A(KEYINPUT71), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n341) );
  XOR2_X1 U348 ( .A(G36GAT), .B(G190GAT), .Z(n411) );
  XNOR2_X1 U349 ( .A(n341), .B(n411), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U351 ( .A(G106GAT), .B(G92GAT), .Z(n300) );
  NAND2_X1 U352 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XOR2_X1 U353 ( .A(n300), .B(n299), .Z(n301) );
  XNOR2_X1 U354 ( .A(n302), .B(n301), .ZN(n307) );
  XOR2_X1 U355 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n304) );
  XNOR2_X1 U356 ( .A(G134GAT), .B(KEYINPUT78), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U358 ( .A(G50GAT), .B(G162GAT), .Z(n431) );
  XNOR2_X1 U359 ( .A(n305), .B(n431), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n560) );
  XOR2_X1 U361 ( .A(KEYINPUT92), .B(KEYINPUT6), .Z(n309) );
  XNOR2_X1 U362 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U364 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n311) );
  XNOR2_X1 U365 ( .A(G120GAT), .B(KEYINPUT5), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U368 ( .A(KEYINPUT94), .B(G57GAT), .Z(n315) );
  XNOR2_X1 U369 ( .A(G29GAT), .B(G148GAT), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U372 ( .A(n318), .B(KEYINPUT91), .Z(n322) );
  XOR2_X1 U373 ( .A(KEYINPUT0), .B(KEYINPUT83), .Z(n320) );
  XNOR2_X1 U374 ( .A(G113GAT), .B(G134GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n443) );
  XNOR2_X1 U376 ( .A(n443), .B(G127GAT), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n329) );
  XOR2_X1 U378 ( .A(G155GAT), .B(KEYINPUT2), .Z(n324) );
  XNOR2_X1 U379 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n423) );
  XOR2_X1 U381 ( .A(G85GAT), .B(n423), .Z(n326) );
  NAND2_X1 U382 ( .A1(G225GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U384 ( .A(G162GAT), .B(n327), .Z(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n520) );
  XOR2_X1 U386 ( .A(G197GAT), .B(KEYINPUT29), .Z(n331) );
  XNOR2_X1 U387 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n345) );
  XOR2_X1 U389 ( .A(KEYINPUT70), .B(G15GAT), .Z(n333) );
  XNOR2_X1 U390 ( .A(G113GAT), .B(G141GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U392 ( .A(n334), .B(G36GAT), .Z(n336) );
  XOR2_X1 U393 ( .A(G169GAT), .B(G8GAT), .Z(n409) );
  XNOR2_X1 U394 ( .A(n409), .B(G50GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U396 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n338) );
  NAND2_X1 U397 ( .A1(G229GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U399 ( .A(n340), .B(n339), .Z(n343) );
  XOR2_X1 U400 ( .A(G1GAT), .B(G22GAT), .Z(n361) );
  XNOR2_X1 U401 ( .A(n341), .B(n361), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n573) );
  XNOR2_X1 U404 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n365) );
  XOR2_X1 U405 ( .A(KEYINPUT36), .B(n560), .Z(n584) );
  XOR2_X1 U406 ( .A(G57GAT), .B(KEYINPUT13), .Z(n367) );
  XOR2_X1 U407 ( .A(n367), .B(G78GAT), .Z(n347) );
  NAND2_X1 U408 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U410 ( .A(G211GAT), .B(KEYINPUT15), .Z(n349) );
  XNOR2_X1 U411 ( .A(KEYINPUT12), .B(KEYINPUT79), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U413 ( .A(n351), .B(n350), .Z(n356) );
  XOR2_X1 U414 ( .A(G64GAT), .B(KEYINPUT14), .Z(n353) );
  XNOR2_X1 U415 ( .A(G8GAT), .B(G183GAT), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U417 ( .A(G71GAT), .B(n354), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U419 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n358) );
  XNOR2_X1 U420 ( .A(G155GAT), .B(KEYINPUT82), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U422 ( .A(n360), .B(n359), .Z(n363) );
  XOR2_X1 U423 ( .A(G15GAT), .B(G127GAT), .Z(n449) );
  XNOR2_X1 U424 ( .A(n361), .B(n449), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n582) );
  NAND2_X1 U426 ( .A1(n584), .A2(n582), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n385) );
  XOR2_X1 U428 ( .A(n367), .B(n366), .Z(n369) );
  NAND2_X1 U429 ( .A1(G230GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U431 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n371) );
  XNOR2_X1 U432 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U434 ( .A(n373), .B(n372), .Z(n378) );
  XOR2_X1 U435 ( .A(G120GAT), .B(G71GAT), .Z(n448) );
  XOR2_X1 U436 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n375) );
  XNOR2_X1 U437 ( .A(G148GAT), .B(G106GAT), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U439 ( .A(G78GAT), .B(n376), .Z(n437) );
  XNOR2_X1 U440 ( .A(n448), .B(n437), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n384) );
  XOR2_X1 U442 ( .A(G204GAT), .B(G64GAT), .Z(n380) );
  XNOR2_X1 U443 ( .A(G176GAT), .B(G92GAT), .ZN(n379) );
  XNOR2_X1 U444 ( .A(n380), .B(n379), .ZN(n400) );
  XNOR2_X1 U445 ( .A(n400), .B(KEYINPUT76), .ZN(n382) );
  INV_X1 U446 ( .A(KEYINPUT33), .ZN(n381) );
  NOR2_X1 U447 ( .A1(n385), .A2(n387), .ZN(n386) );
  NAND2_X1 U448 ( .A1(n573), .A2(n386), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n387), .B(KEYINPUT41), .ZN(n563) );
  NOR2_X1 U450 ( .A1(n573), .A2(n563), .ZN(n389) );
  INV_X1 U451 ( .A(KEYINPUT46), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n389), .B(n388), .ZN(n391) );
  INV_X1 U453 ( .A(n560), .ZN(n545) );
  NOR2_X1 U454 ( .A1(n582), .A2(n545), .ZN(n390) );
  NAND2_X1 U455 ( .A1(n391), .A2(n390), .ZN(n393) );
  XOR2_X1 U456 ( .A(KEYINPUT47), .B(KEYINPUT112), .Z(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  NAND2_X1 U458 ( .A1(n395), .A2(n394), .ZN(n397) );
  XOR2_X1 U459 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n399) );
  XNOR2_X1 U460 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n450) );
  XNOR2_X1 U462 ( .A(n450), .B(n400), .ZN(n416) );
  XNOR2_X1 U463 ( .A(G218GAT), .B(G211GAT), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n401), .B(KEYINPUT89), .ZN(n403) );
  INV_X1 U465 ( .A(KEYINPUT88), .ZN(n402) );
  NAND2_X1 U466 ( .A1(n403), .A2(n402), .ZN(n406) );
  INV_X1 U467 ( .A(n403), .ZN(n404) );
  NAND2_X1 U468 ( .A1(n404), .A2(KEYINPUT88), .ZN(n405) );
  NAND2_X1 U469 ( .A1(n406), .A2(n405), .ZN(n408) );
  XNOR2_X1 U470 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n427) );
  XNOR2_X1 U472 ( .A(n409), .B(n427), .ZN(n412) );
  XOR2_X1 U473 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n410) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n522), .B(KEYINPUT120), .ZN(n417) );
  NOR2_X1 U477 ( .A1(n530), .A2(n417), .ZN(n420) );
  XOR2_X1 U478 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n418) );
  NAND2_X1 U479 ( .A1(n520), .A2(n421), .ZN(n422) );
  XOR2_X1 U480 ( .A(KEYINPUT64), .B(n422), .Z(n571) );
  XOR2_X1 U481 ( .A(n423), .B(KEYINPUT24), .Z(n425) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n435) );
  XOR2_X1 U485 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n429) );
  XNOR2_X1 U486 ( .A(KEYINPUT90), .B(KEYINPUT87), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U488 ( .A(n430), .B(G204GAT), .Z(n433) );
  XNOR2_X1 U489 ( .A(G22GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n465) );
  NAND2_X1 U493 ( .A1(n571), .A2(n465), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n438), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U495 ( .A(G176GAT), .B(G99GAT), .Z(n440) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G190GAT), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n455) );
  XOR2_X1 U498 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n442) );
  XNOR2_X1 U499 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n441) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n447) );
  XOR2_X1 U501 ( .A(n443), .B(KEYINPUT85), .Z(n445) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n447), .B(n446), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n455), .B(n454), .ZN(n466) );
  NAND2_X1 U509 ( .A1(n456), .A2(n466), .ZN(n568) );
  NOR2_X1 U510 ( .A1(n560), .A2(n568), .ZN(n460) );
  XNOR2_X1 U511 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n458) );
  INV_X1 U512 ( .A(G190GAT), .ZN(n457) );
  XNOR2_X1 U513 ( .A(KEYINPUT28), .B(n465), .ZN(n534) );
  INV_X1 U514 ( .A(KEYINPUT101), .ZN(n473) );
  INV_X1 U515 ( .A(n466), .ZN(n536) );
  NAND2_X1 U516 ( .A1(n461), .A2(n465), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n462), .B(KEYINPUT100), .ZN(n464) );
  XOR2_X1 U518 ( .A(n522), .B(KEYINPUT27), .Z(n475) );
  NOR2_X1 U519 ( .A1(n466), .A2(n465), .ZN(n468) );
  XNOR2_X1 U520 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n467) );
  XNOR2_X1 U521 ( .A(n468), .B(n467), .ZN(n469) );
  XOR2_X1 U522 ( .A(KEYINPUT97), .B(n469), .Z(n572) );
  NAND2_X1 U523 ( .A1(n475), .A2(n572), .ZN(n470) );
  NAND2_X1 U524 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U525 ( .A(n473), .B(n472), .ZN(n474) );
  NAND2_X1 U526 ( .A1(n474), .A2(n520), .ZN(n479) );
  INV_X1 U527 ( .A(n475), .ZN(n476) );
  NOR2_X1 U528 ( .A1(n520), .A2(n476), .ZN(n531) );
  AND2_X1 U529 ( .A1(n534), .A2(n536), .ZN(n477) );
  NAND2_X1 U530 ( .A1(n531), .A2(n477), .ZN(n478) );
  NAND2_X1 U531 ( .A1(n479), .A2(n478), .ZN(n480) );
  XOR2_X1 U532 ( .A(KEYINPUT102), .B(n480), .Z(n492) );
  NOR2_X1 U533 ( .A1(n582), .A2(n492), .ZN(n481) );
  NAND2_X1 U534 ( .A1(n481), .A2(n584), .ZN(n482) );
  XNOR2_X1 U535 ( .A(n482), .B(KEYINPUT37), .ZN(n519) );
  NOR2_X1 U536 ( .A1(n387), .A2(n573), .ZN(n493) );
  NAND2_X1 U537 ( .A1(n519), .A2(n493), .ZN(n483) );
  XNOR2_X1 U538 ( .A(KEYINPUT38), .B(n483), .ZN(n505) );
  NOR2_X1 U539 ( .A1(n534), .A2(n505), .ZN(n486) );
  INV_X1 U540 ( .A(G50GAT), .ZN(n484) );
  NOR2_X1 U541 ( .A1(n505), .A2(n520), .ZN(n489) );
  XNOR2_X1 U542 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n487) );
  XNOR2_X1 U543 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  NAND2_X1 U544 ( .A1(n560), .A2(n582), .ZN(n490) );
  XNOR2_X1 U545 ( .A(KEYINPUT16), .B(n490), .ZN(n491) );
  NOR2_X1 U546 ( .A1(n492), .A2(n491), .ZN(n509) );
  NAND2_X1 U547 ( .A1(n509), .A2(n493), .ZN(n494) );
  XOR2_X1 U548 ( .A(KEYINPUT103), .B(n494), .Z(n502) );
  NOR2_X1 U549 ( .A1(n520), .A2(n502), .ZN(n495) );
  XOR2_X1 U550 ( .A(KEYINPUT34), .B(n495), .Z(n496) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(n496), .ZN(G1324GAT) );
  NOR2_X1 U552 ( .A1(n522), .A2(n502), .ZN(n497) );
  XOR2_X1 U553 ( .A(G8GAT), .B(n497), .Z(G1325GAT) );
  NOR2_X1 U554 ( .A1(n502), .A2(n536), .ZN(n501) );
  XOR2_X1 U555 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n499) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U558 ( .A(n501), .B(n500), .ZN(G1326GAT) );
  NOR2_X1 U559 ( .A1(n534), .A2(n502), .ZN(n503) );
  XOR2_X1 U560 ( .A(G22GAT), .B(n503), .Z(G1327GAT) );
  NOR2_X1 U561 ( .A1(n522), .A2(n505), .ZN(n504) );
  XOR2_X1 U562 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  NOR2_X1 U563 ( .A1(n536), .A2(n505), .ZN(n507) );
  XNOR2_X1 U564 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n506) );
  XNOR2_X1 U565 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U566 ( .A(n508), .B(G43GAT), .ZN(G1330GAT) );
  INV_X1 U567 ( .A(n573), .ZN(n537) );
  NOR2_X1 U568 ( .A1(n537), .A2(n563), .ZN(n518) );
  NAND2_X1 U569 ( .A1(n509), .A2(n518), .ZN(n515) );
  NOR2_X1 U570 ( .A1(n520), .A2(n515), .ZN(n511) );
  XNOR2_X1 U571 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n522), .A2(n515), .ZN(n513) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n513), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n536), .A2(n515), .ZN(n514) );
  XOR2_X1 U577 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U578 ( .A1(n534), .A2(n515), .ZN(n517) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U581 ( .A1(n519), .A2(n518), .ZN(n527) );
  NOR2_X1 U582 ( .A1(n520), .A2(n527), .ZN(n521) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n521), .Z(G1336GAT) );
  NOR2_X1 U584 ( .A1(n522), .A2(n527), .ZN(n523) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n536), .A2(n527), .ZN(n525) );
  XNOR2_X1 U587 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(n526), .ZN(G1338GAT) );
  NOR2_X1 U590 ( .A1(n534), .A2(n527), .ZN(n528) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  INV_X1 U593 ( .A(n531), .ZN(n532) );
  NOR2_X1 U594 ( .A1(n530), .A2(n532), .ZN(n533) );
  XNOR2_X1 U595 ( .A(KEYINPUT114), .B(n533), .ZN(n549) );
  NAND2_X1 U596 ( .A1(n534), .A2(n549), .ZN(n535) );
  NOR2_X1 U597 ( .A1(n536), .A2(n535), .ZN(n546) );
  NAND2_X1 U598 ( .A1(n546), .A2(n537), .ZN(n538) );
  XNOR2_X1 U599 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  INV_X1 U601 ( .A(n563), .ZN(n539) );
  NAND2_X1 U602 ( .A1(n546), .A2(n539), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n543) );
  NAND2_X1 U605 ( .A1(n546), .A2(n582), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n572), .A2(n549), .ZN(n550) );
  XNOR2_X1 U612 ( .A(KEYINPUT116), .B(n550), .ZN(n559) );
  NOR2_X1 U613 ( .A1(n559), .A2(n573), .ZN(n552) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n551) );
  XNOR2_X1 U615 ( .A(n552), .B(n551), .ZN(G1344GAT) );
  NOR2_X1 U616 ( .A1(n559), .A2(n563), .ZN(n557) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n554) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(KEYINPUT118), .B(n555), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  INV_X1 U622 ( .A(n582), .ZN(n569) );
  NOR2_X1 U623 ( .A1(n559), .A2(n569), .ZN(n558) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n558), .Z(G1346GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  NOR2_X1 U627 ( .A1(n573), .A2(n568), .ZN(n562) );
  XOR2_X1 U628 ( .A(G169GAT), .B(n562), .Z(G1348GAT) );
  NOR2_X1 U629 ( .A1(n568), .A2(n563), .ZN(n567) );
  XOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n565) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U635 ( .A(G183GAT), .B(n570), .Z(G1350GAT) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n579) );
  NOR2_X1 U637 ( .A1(n573), .A2(n579), .ZN(n578) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n575) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT125), .B(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  INV_X1 U644 ( .A(n579), .ZN(n585) );
  NAND2_X1 U645 ( .A1(n585), .A2(n387), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

