//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  AOI21_X1  g000(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n202));
  OAI21_X1  g001(.A(new_n202), .B1(G169gat), .B2(G176gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT26), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n204), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT27), .B(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(KEYINPUT28), .A3(new_n210), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n208), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n218), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n204), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT25), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n226), .A2(new_n223), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n221), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n216), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT29), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G226gat), .A2(G233gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G197gat), .B(G204gat), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT72), .B(G218gat), .Z(new_n239));
  INV_X1    g038(.A(G211gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n238), .B1(new_n241), .B2(KEYINPUT22), .ZN(new_n242));
  XNOR2_X1  g041(.A(G211gat), .B(G218gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n242), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n236), .B(KEYINPUT73), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n233), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n237), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n242), .B(new_n243), .ZN(new_n249));
  INV_X1    g048(.A(new_n236), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n233), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n246), .B1(new_n233), .B2(new_n234), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n249), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G8gat), .B(G36gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT74), .ZN(new_n255));
  XNOR2_X1  g054(.A(G64gat), .B(G92gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n248), .A2(new_n253), .A3(KEYINPUT30), .A4(new_n257), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n258), .A2(KEYINPUT76), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n248), .A2(new_n253), .A3(new_n257), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n257), .B(KEYINPUT75), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n261), .B1(new_n248), .B2(new_n253), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n258), .A2(KEYINPUT76), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n259), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G148gat), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT78), .B1(new_n268), .B2(G141gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT78), .ZN(new_n270));
  INV_X1    g069(.A(G141gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(G148gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(G141gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT79), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(KEYINPUT80), .B(G155gat), .Z(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G162gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n278), .A2(KEYINPUT2), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n276), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n271), .A2(G148gat), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT2), .B1(new_n284), .B2(new_n273), .ZN(new_n285));
  AND2_X1   g084(.A1(new_n279), .A2(KEYINPUT77), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n281), .B1(new_n279), .B2(KEYINPUT77), .ZN(new_n287));
  NOR3_X1   g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n245), .A2(new_n290), .A3(new_n234), .ZN(new_n291));
  NAND2_X1  g090(.A1(G228gat), .A2(G233gat), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n292), .B1(new_n290), .B2(KEYINPUT3), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n288), .B1(new_n276), .B2(new_n282), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT29), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT86), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n245), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(KEYINPUT86), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n294), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G22gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n249), .A2(KEYINPUT29), .ZN(new_n305));
  INV_X1    g104(.A(new_n296), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n290), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n297), .A2(new_n245), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n292), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n303), .A2(new_n304), .A3(new_n311), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n307), .A2(new_n309), .B1(G228gat), .B2(G233gat), .ZN(new_n313));
  OAI21_X1  g112(.A(G22gat), .B1(new_n313), .B2(new_n302), .ZN(new_n314));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT31), .B(G50gat), .ZN(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  NAND4_X1  g116(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT87), .A4(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n312), .A2(KEYINPUT87), .A3(new_n314), .ZN(new_n319));
  INV_X1    g118(.A(new_n317), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT87), .B1(new_n312), .B2(new_n314), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n318), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G227gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G113gat), .ZN(new_n326));
  INV_X1    g125(.A(G120gat), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT1), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(new_n326), .B2(new_n327), .ZN(new_n329));
  INV_X1    g128(.A(G127gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(KEYINPUT66), .A3(G134gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G127gat), .B(G134gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n329), .B(new_n331), .C1(new_n333), .C2(KEYINPUT66), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT67), .B(G113gat), .Z(new_n335));
  OAI211_X1 g134(.A(new_n328), .B(new_n332), .C1(new_n335), .C2(new_n327), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n233), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n216), .B(new_n337), .C1(new_n229), .C2(new_n232), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n325), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT71), .B1(new_n342), .B2(KEYINPUT34), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT71), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT34), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n341), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n342), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT70), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(new_n341), .B2(new_n345), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT32), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n339), .A2(new_n340), .A3(new_n325), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT68), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT68), .A4(new_n325), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n353), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT33), .B1(new_n356), .B2(new_n357), .ZN(new_n359));
  XNOR2_X1  g158(.A(G15gat), .B(G43gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n358), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n356), .A2(new_n357), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT32), .ZN(new_n365));
  INV_X1    g164(.A(new_n362), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n366), .A2(KEYINPUT69), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT33), .B1(new_n366), .B2(KEYINPUT69), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n352), .B1(new_n363), .B2(new_n370), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n343), .A2(new_n346), .B1(new_n348), .B2(new_n350), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n358), .B1(new_n367), .B2(new_n368), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(new_n366), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n372), .B(new_n373), .C1(new_n374), .C2(new_n359), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n323), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n290), .A2(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n295), .A2(new_n296), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n337), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n295), .A2(new_n338), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n295), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n380), .A2(new_n381), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n290), .A2(new_n337), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n382), .ZN(new_n389));
  INV_X1    g188(.A(new_n381), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT83), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n384), .A2(new_n385), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n395), .A2(new_n381), .A3(new_n380), .A4(new_n387), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n386), .A2(KEYINPUT83), .A3(new_n391), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(G57gat), .B(G85gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n398), .A2(KEYINPUT6), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n398), .B2(new_n403), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n397), .A2(new_n396), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT83), .B1(new_n386), .B2(new_n391), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n398), .A2(KEYINPUT84), .A3(new_n403), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n404), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI211_X1 g214(.A(KEYINPUT85), .B(new_n406), .C1(new_n411), .C2(new_n412), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n267), .B(new_n377), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT35), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n267), .A2(new_n371), .A3(new_n375), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n323), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n407), .A2(new_n408), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT6), .B1(new_n421), .B2(new_n402), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT88), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n409), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n398), .A2(KEYINPUT88), .A3(new_n403), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n422), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT35), .B1(new_n426), .B2(new_n404), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n267), .B1(new_n415), .B2(new_n416), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n323), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n376), .B(KEYINPUT36), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n395), .A2(new_n380), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n390), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n388), .A2(new_n381), .A3(new_n382), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(KEYINPUT39), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT39), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n432), .A2(new_n436), .A3(new_n390), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n402), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT40), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n435), .A2(KEYINPUT40), .A3(new_n402), .A4(new_n437), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n266), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n425), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(new_n323), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n248), .A2(new_n253), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n446), .A2(KEYINPUT37), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n237), .A2(new_n249), .A3(new_n247), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n245), .B1(new_n251), .B2(new_n252), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT37), .ZN(new_n450));
  XOR2_X1   g249(.A(KEYINPUT89), .B(KEYINPUT38), .Z(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n261), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n447), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n260), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n257), .B1(new_n446), .B2(KEYINPUT37), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n451), .B1(new_n447), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(new_n426), .A3(new_n404), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n431), .B1(new_n445), .B2(new_n459), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n418), .A2(new_n428), .B1(new_n430), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT94), .ZN(new_n462));
  NAND2_X1  g261(.A1(G229gat), .A2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT16), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(G1gat), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n467), .B(KEYINPUT93), .C1(G1gat), .C2(new_n465), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(G8gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G43gat), .B(G50gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT15), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NOR3_X1   g274(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n476));
  OAI22_X1  g275(.A1(new_n471), .A2(KEYINPUT15), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G29gat), .A2(G36gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n473), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NOR4_X1   g279(.A1(KEYINPUT90), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n482));
  NOR2_X1   g281(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n483));
  INV_X1    g282(.A(G36gat), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n474), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT91), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(new_n474), .C1(new_n481), .C2(new_n485), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n489), .A3(new_n478), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n480), .B1(new_n490), .B2(new_n473), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n470), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT92), .B1(new_n491), .B2(KEYINPUT17), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT92), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n479), .B1(new_n486), .B2(KEYINPUT91), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n472), .B1(new_n496), .B2(new_n489), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n494), .B(new_n495), .C1(new_n497), .C2(new_n480), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n469), .B1(KEYINPUT17), .B2(new_n491), .ZN(new_n500));
  AOI211_X1 g299(.A(new_n464), .B(new_n492), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n462), .B1(new_n501), .B2(KEYINPUT18), .ZN(new_n502));
  XNOR2_X1  g301(.A(G113gat), .B(G141gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(G197gat), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT11), .B(G169gat), .Z(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT12), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n491), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(new_n469), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n463), .B(KEYINPUT13), .Z(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n501), .B2(KEYINPUT18), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n499), .A2(new_n500), .ZN(new_n514));
  INV_X1    g313(.A(new_n492), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n514), .A2(KEYINPUT18), .A3(new_n463), .A4(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n502), .B(new_n508), .C1(new_n513), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n463), .A3(new_n515), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT18), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n519), .A2(new_n520), .B1(new_n510), .B2(new_n511), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT94), .B1(new_n519), .B2(new_n520), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n521), .B(new_n516), .C1(new_n522), .C2(new_n507), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n461), .A2(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(G134gat), .B(G162gat), .Z(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(KEYINPUT41), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n490), .A2(new_n473), .ZN(new_n532));
  INV_X1    g331(.A(new_n480), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(KEYINPUT17), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(KEYINPUT100), .A3(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g335(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(G85gat), .A3(G92gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT101), .ZN(new_n541));
  NAND2_X1  g340(.A1(G99gat), .A2(G106gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G85gat), .ZN(new_n544));
  INV_X1    g343(.A(G92gat), .ZN(new_n545));
  AOI22_X1  g344(.A1(KEYINPUT8), .A2(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n539), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n541), .B1(new_n540), .B2(new_n542), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n548), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n550), .A2(new_n539), .A3(new_n543), .A4(new_n546), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(new_n493), .B2(new_n498), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n529), .A2(KEYINPUT41), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n491), .B2(new_n553), .ZN(new_n557));
  OAI21_X1  g356(.A(G190gat), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n552), .B1(new_n491), .B2(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n499), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n557), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n210), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G218gat), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT99), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n562), .A3(G218gat), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n531), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n210), .B1(new_n560), .B2(new_n561), .ZN(new_n568));
  AOI211_X1 g367(.A(G190gat), .B(new_n557), .C1(new_n499), .C2(new_n559), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n564), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT99), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n570), .A2(new_n571), .A3(new_n566), .A4(new_n531), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n528), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(G57gat), .A2(G64gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT95), .ZN(new_n576));
  NAND2_X1  g375(.A1(G57gat), .A2(G64gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(G57gat), .A2(G64gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(G57gat), .A2(G64gat), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT95), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT97), .ZN(new_n584));
  NAND2_X1  g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT96), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OR2_X1    g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT96), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n589), .A2(new_n590), .A3(new_n585), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n582), .A2(new_n584), .A3(new_n588), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n575), .A2(KEYINPUT9), .A3(new_n577), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n585), .A3(new_n589), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT21), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(new_n330), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n588), .A2(new_n591), .A3(new_n578), .A4(new_n581), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT97), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n583), .B(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n594), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g403(.A(KEYINPUT98), .B(new_n594), .C1(new_n599), .C2(new_n601), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(KEYINPUT21), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n470), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n598), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G155gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n570), .A2(new_n571), .A3(new_n566), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n530), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(new_n527), .A3(new_n572), .ZN(new_n618));
  INV_X1    g417(.A(G230gat), .ZN(new_n619));
  INV_X1    g418(.A(G233gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n592), .A2(new_n594), .A3(new_n549), .A4(new_n551), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n552), .A2(new_n602), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT10), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(new_n549), .B2(new_n551), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n604), .A2(new_n605), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n622), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n623), .A2(new_n624), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n621), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n629), .A2(new_n631), .A3(new_n635), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n574), .A2(new_n615), .A3(new_n618), .A4(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n526), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n415), .A2(new_n416), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g446(.A(KEYINPUT16), .B(G8gat), .Z(new_n648));
  NAND3_X1  g447(.A1(new_n644), .A2(new_n266), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(G8gat), .B1(new_n643), .B2(new_n267), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  MUX2_X1   g450(.A(new_n649), .B(new_n651), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g451(.A(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n376), .B(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(G15gat), .B1(new_n643), .B2(new_n654), .ZN(new_n655));
  OR2_X1    g454(.A1(new_n376), .A2(G15gat), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n655), .B1(new_n643), .B2(new_n656), .ZN(G1326gat));
  NAND3_X1  g456(.A1(new_n644), .A2(KEYINPUT102), .A3(new_n323), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  INV_X1    g458(.A(new_n323), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n643), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT43), .B(G22gat), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n658), .B2(new_n661), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(G1327gat));
  AND3_X1   g464(.A1(new_n617), .A2(new_n527), .A3(new_n572), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n527), .B1(new_n617), .B2(new_n572), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n668), .A2(new_n615), .A3(new_n639), .ZN(new_n669));
  INV_X1    g468(.A(new_n459), .ZN(new_n670));
  INV_X1    g469(.A(new_n322), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n319), .A3(new_n320), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n672), .B(new_n318), .C1(new_n443), .C2(new_n442), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n654), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n674), .B1(new_n323), .B2(new_n429), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n417), .A2(KEYINPUT35), .B1(new_n420), .B2(new_n427), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n524), .B(new_n669), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n415), .A2(new_n416), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(G29gat), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT45), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT45), .ZN(new_n682));
  NOR4_X1   g481(.A1(new_n677), .A2(new_n682), .A3(G29gat), .A4(new_n679), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n461), .B2(new_n668), .ZN(new_n686));
  INV_X1    g485(.A(new_n668), .ZN(new_n687));
  OAI211_X1 g486(.A(KEYINPUT44), .B(new_n687), .C1(new_n675), .C2(new_n676), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n615), .A2(new_n639), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n524), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n518), .A2(new_n523), .A3(KEYINPUT103), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n686), .A2(new_n645), .A3(new_n688), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G29gat), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n684), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n684), .A2(KEYINPUT104), .A3(new_n696), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1328gat));
  NOR3_X1   g500(.A1(new_n677), .A2(G36gat), .A3(new_n267), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT46), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n704), .A2(new_n266), .A3(new_n694), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n705), .B2(new_n484), .ZN(G1329gat));
  NAND4_X1  g505(.A1(new_n686), .A2(new_n431), .A3(new_n688), .A4(new_n694), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G43gat), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n677), .A2(G43gat), .A3(new_n376), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT47), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n710), .B(new_n712), .ZN(G1330gat));
  OR3_X1    g512(.A1(new_n677), .A2(G50gat), .A3(new_n660), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n714), .A2(KEYINPUT48), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n686), .A2(new_n323), .A3(new_n688), .A4(new_n694), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G50gat), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n716), .A2(new_n717), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n715), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n716), .A2(G50gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n714), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n721), .A2(new_n725), .ZN(G1331gat));
  NAND2_X1  g525(.A1(new_n418), .A2(new_n428), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n430), .A2(new_n460), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n615), .ZN(new_n730));
  NOR4_X1   g529(.A1(new_n687), .A2(new_n693), .A3(new_n730), .A4(new_n640), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n679), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n645), .A2(KEYINPUT107), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  INV_X1    g537(.A(KEYINPUT49), .ZN(new_n739));
  INV_X1    g538(.A(G64gat), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n732), .B(new_n266), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1333gat));
  INV_X1    g542(.A(G71gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n731), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n376), .B(KEYINPUT109), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR4_X1   g546(.A1(new_n745), .A2(KEYINPUT108), .A3(new_n744), .A4(new_n654), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n654), .A2(new_n744), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n732), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n747), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g552(.A1(new_n732), .A2(new_n323), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g554(.A1(new_n693), .A2(new_n615), .A3(new_n640), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n704), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757), .B2(new_n679), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n693), .A2(new_n615), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n687), .B(new_n759), .C1(new_n675), .C2(new_n676), .ZN(new_n760));
  NAND2_X1  g559(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT110), .B(KEYINPUT51), .Z(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n729), .A2(new_n687), .A3(new_n759), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n645), .A2(new_n544), .A3(new_n639), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n758), .B1(new_n767), .B2(new_n768), .ZN(G1336gat));
  NAND4_X1  g568(.A1(new_n686), .A2(new_n266), .A3(new_n688), .A4(new_n756), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G92gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n266), .A2(new_n545), .A3(new_n639), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n767), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT52), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n771), .B(new_n775), .C1(new_n767), .C2(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1337gat));
  OAI21_X1  g576(.A(G99gat), .B1(new_n757), .B2(new_n654), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n376), .A2(G99gat), .A3(new_n640), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT111), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n767), .B2(new_n780), .ZN(G1338gat));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n660), .A2(new_n640), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n766), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(G106gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n660), .A2(new_n788), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n686), .A2(new_n688), .A3(new_n756), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n782), .A2(new_n783), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n785), .B1(new_n789), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(G106gat), .B1(new_n766), .B2(new_n786), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n796), .A2(new_n793), .A3(new_n784), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n795), .A2(new_n797), .ZN(G1339gat));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n604), .A2(new_n627), .A3(new_n605), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n621), .B(new_n800), .C1(new_n630), .C2(KEYINPUT10), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n801), .A2(new_n629), .A3(KEYINPUT54), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n803), .B(new_n622), .C1(new_n625), .C2(new_n628), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n636), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n804), .A2(KEYINPUT113), .A3(new_n636), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n802), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n799), .B1(new_n809), .B2(KEYINPUT55), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n801), .A2(new_n629), .A3(KEYINPUT54), .ZN(new_n811));
  INV_X1    g610(.A(new_n808), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT113), .B1(new_n804), .B2(new_n636), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(KEYINPUT114), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT55), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n638), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n691), .B2(new_n692), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n519), .A2(new_n520), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n822), .A2(new_n507), .A3(new_n516), .A4(new_n512), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n463), .B1(new_n514), .B2(new_n515), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n510), .A2(new_n511), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n506), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n823), .A2(new_n639), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n668), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n823), .A2(new_n826), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n817), .A2(new_n829), .A3(new_n819), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n666), .B2(new_n667), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n615), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n641), .A2(new_n693), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n660), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n679), .A2(new_n419), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n525), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n834), .A2(new_n420), .A3(new_n736), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n335), .A3(new_n693), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(G1340gat));
  OAI21_X1  g640(.A(G120gat), .B1(new_n837), .B2(new_n640), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n839), .A2(new_n327), .A3(new_n639), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n843), .B1(new_n842), .B2(new_n844), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(G1341gat));
  NOR3_X1   g646(.A1(new_n837), .A2(new_n330), .A3(new_n730), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n839), .A2(new_n615), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n849), .A2(KEYINPUT116), .ZN(new_n850));
  AOI21_X1  g649(.A(G127gat), .B1(new_n849), .B2(KEYINPUT116), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(G1342gat));
  AOI21_X1  g651(.A(G134gat), .B1(KEYINPUT117), .B2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n839), .A2(new_n687), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n835), .A2(new_n687), .A3(new_n836), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n858), .A2(new_n859), .A3(G134gat), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n858), .B2(G134gat), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n856), .B(new_n857), .C1(new_n860), .C2(new_n861), .ZN(G1343gat));
  NAND3_X1  g661(.A1(new_n645), .A2(new_n267), .A3(new_n654), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT119), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n814), .A2(new_n815), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n638), .A3(new_n818), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n523), .B2(new_n518), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n574), .B(new_n618), .C1(new_n867), .C2(new_n827), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n615), .B1(new_n868), .B2(new_n831), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT57), .B(new_n323), .C1(new_n869), .C2(new_n833), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g671(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n834), .B2(new_n323), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n864), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G141gat), .B1(new_n875), .B2(new_n525), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n834), .A2(new_n736), .ZN(new_n877));
  NOR4_X1   g676(.A1(new_n877), .A2(new_n660), .A3(new_n266), .A4(new_n431), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n525), .A2(G141gat), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT58), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n693), .B(new_n864), .C1(new_n872), .C2(new_n874), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n882), .A2(G141gat), .B1(new_n878), .B2(new_n879), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(G1344gat));
  NOR2_X1   g684(.A1(new_n268), .A2(KEYINPUT59), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n875), .B2(new_n640), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n323), .B(new_n873), .C1(new_n832), .C2(new_n833), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n641), .A2(new_n524), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n323), .B1(new_n869), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n893), .A2(new_n639), .A3(new_n864), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT59), .B1(new_n894), .B2(new_n268), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n878), .A2(new_n268), .A3(new_n639), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1345gat));
  OAI21_X1  g697(.A(new_n277), .B1(new_n875), .B2(new_n730), .ZN(new_n899));
  INV_X1    g698(.A(new_n277), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n878), .A2(new_n900), .A3(new_n615), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1346gat));
  INV_X1    g701(.A(G162gat), .ZN(new_n903));
  OR3_X1    g702(.A1(new_n875), .A2(new_n903), .A3(new_n668), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n878), .A2(new_n687), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n903), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n904), .A2(new_n906), .ZN(G1347gat));
  NOR3_X1   g706(.A1(new_n736), .A2(new_n267), .A3(new_n746), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n835), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n205), .A3(new_n525), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n834), .A2(new_n679), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n323), .A2(new_n267), .A3(new_n376), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n693), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n910), .B1(new_n205), .B2(new_n915), .ZN(G1348gat));
  OAI21_X1  g715(.A(G176gat), .B1(new_n909), .B2(new_n640), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n639), .A2(new_n206), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n913), .B2(new_n918), .ZN(G1349gat));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(KEYINPUT122), .B2(KEYINPUT60), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n908), .A2(new_n834), .A3(new_n660), .A4(new_n615), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G183gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n615), .A2(new_n209), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n913), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n920), .A2(KEYINPUT60), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n928), .B1(new_n922), .B2(new_n926), .ZN(G1350gat));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n210), .A3(new_n687), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n835), .A2(new_n687), .A3(new_n908), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n931), .A2(new_n932), .A3(G190gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n931), .B2(G190gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G1351gat));
  NOR3_X1   g734(.A1(new_n431), .A2(new_n660), .A3(new_n267), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n911), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n693), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n734), .A2(new_n266), .A3(new_n654), .A4(new_n735), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n888), .B2(new_n892), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n524), .A2(G197gat), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  INV_X1    g742(.A(G204gat), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n639), .A2(new_n944), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n937), .A2(KEYINPUT62), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT62), .B1(new_n937), .B2(new_n945), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n941), .A2(new_n639), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n946), .B(new_n947), .C1(new_n944), .C2(new_n948), .ZN(G1353gat));
  NOR2_X1   g748(.A1(new_n730), .A2(G211gat), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  OR3_X1    g750(.A1(new_n937), .A2(KEYINPUT124), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT124), .B1(new_n937), .B2(new_n951), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n940), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n893), .A2(new_n615), .A3(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g757(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n941), .A2(KEYINPUT125), .A3(new_n615), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n958), .A2(G211gat), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI211_X1 g762(.A(new_n730), .B(new_n940), .C1(new_n888), .C2(new_n892), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n240), .B1(new_n964), .B2(KEYINPUT125), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n959), .B1(new_n965), .B2(new_n958), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n954), .B1(new_n963), .B2(new_n966), .ZN(G1354gat));
  AOI21_X1  g766(.A(G218gat), .B1(new_n938), .B2(new_n687), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n668), .A2(new_n239), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n941), .B2(new_n969), .ZN(G1355gat));
endmodule


