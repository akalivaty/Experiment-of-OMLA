//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n468), .A2(KEYINPUT69), .A3(new_n472), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n471), .A2(G137), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n478), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n462), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n465), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n464), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n477), .A2(new_n482), .B1(G101), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n475), .A2(new_n476), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G112), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n472), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n481), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT71), .Z(new_n492));
  NAND2_X1  g067(.A1(new_n482), .A2(new_n472), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI211_X1 g069(.A(new_n489), .B(new_n492), .C1(G124), .C2(new_n494), .ZN(G162));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OR2_X1    g071(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(G138), .A3(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n481), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n500), .B2(KEYINPUT73), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n481), .B2(new_n499), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n496), .A2(KEYINPUT74), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT3), .B(G2104), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n510), .B2(new_n499), .ZN(new_n511));
  INV_X1    g086(.A(G138), .ZN(new_n512));
  NOR3_X1   g087(.A1(new_n469), .A2(new_n470), .A3(new_n512), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n513), .A2(KEYINPUT75), .A3(new_n509), .A4(new_n508), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n501), .A2(new_n503), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(G126), .A2(G2105), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n479), .A2(new_n480), .A3(new_n465), .A4(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(G102), .A2(G2105), .ZN(new_n518));
  INV_X1    g093(.A(G2105), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n518), .B(G2104), .C1(G114), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT72), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT76), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n480), .A2(new_n465), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n524), .A2(new_n513), .A3(KEYINPUT73), .A4(new_n479), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(new_n503), .A3(KEYINPUT4), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n511), .A2(new_n514), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n521), .B(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n523), .A2(new_n532), .ZN(G164));
  NAND2_X1  g108(.A1(KEYINPUT77), .A2(G651), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT6), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G50), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT78), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT5), .B(G543), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G75), .A2(G543), .ZN(new_n543));
  XOR2_X1   g118(.A(KEYINPUT5), .B(G543), .Z(new_n544));
  INV_X1    g119(.A(G62), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n542), .A2(G88), .B1(new_n546), .B2(G651), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n540), .A2(new_n547), .ZN(G303));
  INV_X1    g123(.A(G303), .ZN(G166));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT79), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT7), .ZN(new_n552));
  INV_X1    g127(.A(G51), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n537), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n536), .A2(G89), .ZN(new_n555));
  NAND2_X1  g130(.A1(G63), .A2(G651), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n544), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(G168));
  NAND2_X1  g133(.A1(new_n538), .A2(G52), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n542), .A2(G90), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n541), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G651), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(G301));
  INV_X1    g139(.A(G301), .ZN(G171));
  NAND2_X1  g140(.A1(G68), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G56), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n544), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n538), .A2(G43), .B1(new_n568), .B2(G651), .ZN(new_n569));
  XOR2_X1   g144(.A(KEYINPUT80), .B(G81), .Z(new_n570));
  NAND2_X1  g145(.A1(new_n542), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  NAND4_X1  g149(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND4_X1  g152(.A1(G319), .A2(G483), .A3(G661), .A4(new_n577), .ZN(G188));
  AOI22_X1  g153(.A1(new_n541), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n562), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT82), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G53), .ZN(new_n583));
  OR3_X1    g158(.A1(new_n537), .A2(KEYINPUT9), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT9), .B1(new_n537), .B2(new_n583), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n542), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n536), .A2(new_n541), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT81), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(G91), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n582), .A2(new_n586), .A3(new_n591), .ZN(G299));
  INV_X1    g167(.A(G168), .ZN(G286));
  AND2_X1   g168(.A1(new_n588), .A2(new_n590), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G87), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n541), .A2(G74), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n538), .A2(G49), .B1(G651), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(G288));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G61), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n544), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n538), .A2(G48), .B1(new_n601), .B2(G651), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n588), .A2(new_n590), .ZN(new_n603));
  INV_X1    g178(.A(G86), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(G305));
  NAND2_X1  g180(.A1(new_n538), .A2(G47), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n542), .A2(G85), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n541), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n606), .B(new_n607), .C1(new_n562), .C2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n594), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n603), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n541), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n538), .A2(G54), .B1(new_n617), .B2(G651), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n610), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n610), .B1(new_n619), .B2(G868), .ZN(G321));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(G299), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(G168), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(new_n622), .B2(G168), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n572), .A2(new_n622), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n615), .A2(new_n618), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n630), .B2(new_n622), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n509), .A2(new_n483), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT12), .Z(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  INV_X1    g211(.A(G111), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  AOI22_X1  g214(.A1(new_n472), .A2(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n638), .B2(new_n639), .ZN(new_n641));
  INV_X1    g216(.A(G123), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n641), .B1(new_n493), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(G135), .B2(new_n490), .ZN(new_n644));
  INV_X1    g219(.A(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n644), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(G2096), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n636), .A2(new_n646), .A3(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n650));
  XOR2_X1   g225(.A(KEYINPUT15), .B(G2435), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2438), .ZN(new_n652));
  XOR2_X1   g227(.A(G2427), .B(G2430), .Z(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n652), .B2(new_n653), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G14), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(G2100), .Z(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n645), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n680), .A2(new_n681), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n679), .A2(new_n684), .A3(new_n682), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n679), .A2(new_n684), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n687));
  AOI211_X1 g262(.A(new_n683), .B(new_n685), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n686), .B2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT86), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n693), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n692), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n695), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n696), .A2(new_n700), .ZN(G229));
  XNOR2_X1  g276(.A(KEYINPUT92), .B(KEYINPUT36), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G22), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT90), .Z(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G303), .B2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G1971), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n707), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT91), .ZN(new_n713));
  MUX2_X1   g288(.A(G6), .B(G305), .S(G16), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n704), .A2(G23), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n595), .A2(new_n597), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(new_n704), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT33), .B(G1976), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n710), .A2(new_n713), .A3(new_n716), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT34), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G25), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT87), .ZN(new_n726));
  OAI221_X1 g301(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n471), .C2(G107), .ZN(new_n727));
  INV_X1    g302(.A(G119), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n493), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G131), .B2(new_n490), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT88), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n726), .B1(new_n731), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT89), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  MUX2_X1   g311(.A(G24), .B(G290), .S(G16), .Z(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(G1986), .Z(new_n738));
  NAND3_X1  g313(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n703), .B1(new_n723), .B2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n739), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n722), .A2(KEYINPUT34), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n722), .A2(KEYINPUT34), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n741), .A2(new_n742), .A3(new_n743), .A4(new_n702), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n704), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n573), .B2(new_n704), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT93), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1341), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n724), .A2(G26), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT28), .ZN(new_n751));
  OAI221_X1 g326(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n471), .C2(G116), .ZN(new_n752));
  INV_X1    g327(.A(G128), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n493), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G140), .B2(new_n490), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n751), .B1(new_n755), .B2(new_n724), .ZN(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G4), .A2(G16), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n629), .B2(new_n704), .ZN(new_n761));
  INV_X1    g336(.A(G1348), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n749), .A2(new_n758), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(KEYINPUT94), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(KEYINPUT94), .ZN(new_n767));
  NOR2_X1   g342(.A1(G27), .A2(G29), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G164), .B2(G29), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n766), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G162), .A2(G29), .ZN(new_n773));
  OR2_X1    g348(.A1(G29), .A2(G35), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n775), .A2(KEYINPUT29), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(KEYINPUT29), .ZN(new_n777));
  INV_X1    g352(.A(G2090), .ZN(new_n778));
  OR3_X1    g353(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G16), .A2(G21), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G168), .B2(G16), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT97), .B(G1966), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT24), .ZN(new_n784));
  INV_X1    g359(.A(G34), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n784), .B2(new_n785), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G160), .B2(new_n724), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT26), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n791), .A2(new_n792), .B1(G105), .B2(new_n483), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n494), .B2(G129), .ZN(new_n795));
  INV_X1    g370(.A(G141), .ZN(new_n796));
  INV_X1    g371(.A(new_n490), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n724), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n724), .B2(G32), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT27), .B(G1996), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n783), .B1(G2084), .B2(new_n788), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n704), .A2(G20), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT23), .Z(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G299), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G1956), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G5), .A2(G16), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT98), .Z(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G301), .B2(new_n704), .ZN(new_n811));
  INV_X1    g386(.A(G1961), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT30), .B(G28), .ZN(new_n814));
  OR2_X1    g389(.A1(KEYINPUT31), .A2(G11), .ZN(new_n815));
  NAND2_X1  g390(.A1(KEYINPUT31), .A2(G11), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n814), .A2(new_n724), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n647), .B2(new_n724), .ZN(new_n818));
  NOR4_X1   g393(.A1(new_n803), .A2(new_n808), .A3(new_n813), .A4(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n778), .B1(new_n776), .B2(new_n777), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n779), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n724), .A2(G33), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT25), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n490), .A2(G139), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n509), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(new_n471), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT95), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n823), .B1(new_n830), .B2(G29), .ZN(new_n831));
  INV_X1    g406(.A(G2072), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n801), .A2(new_n802), .B1(G2084), .B2(new_n788), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n832), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT96), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n772), .A2(new_n821), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n745), .A2(KEYINPUT99), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT99), .B1(new_n745), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(G311));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n745), .A2(new_n842), .A3(new_n838), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n745), .B2(new_n838), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(G150));
  NOR2_X1   g420(.A1(new_n629), .A2(new_n626), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  INV_X1    g423(.A(G67), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n544), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n562), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  AOI22_X1  g428(.A1(G55), .A2(new_n538), .B1(new_n542), .B2(G93), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n572), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n847), .B(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n858), .A2(new_n859), .A3(G860), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n855), .A2(G860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT37), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n860), .A2(new_n862), .ZN(G145));
  XNOR2_X1  g438(.A(new_n730), .B(KEYINPUT105), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n634), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n494), .A2(G130), .B1(G142), .B2(new_n490), .ZN(new_n866));
  OR3_X1    g441(.A1(new_n471), .A2(KEYINPUT104), .A3(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT104), .B1(new_n471), .B2(G118), .ZN(new_n868));
  OR2_X1    g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n867), .A2(G2104), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n865), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n829), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n755), .B(KEYINPUT103), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n521), .B1(new_n526), .B2(new_n527), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n798), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n877), .A2(new_n798), .A3(new_n878), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n873), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n830), .A3(new_n879), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n872), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n644), .B(KEYINPUT102), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n485), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(G162), .Z(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n882), .A2(new_n884), .A3(new_n872), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n889), .B1(new_n893), .B2(new_n885), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(KEYINPUT106), .B(G37), .Z(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g473(.A(G303), .B(G290), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n718), .B(G305), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(G303), .B(G290), .ZN(new_n902));
  XNOR2_X1  g477(.A(G288), .B(G305), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n901), .A2(KEYINPUT109), .A3(new_n904), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT109), .B1(new_n901), .B2(new_n904), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  MUX2_X1   g484(.A(new_n905), .B(new_n909), .S(KEYINPUT42), .Z(new_n910));
  XNOR2_X1  g485(.A(new_n630), .B(new_n856), .ZN(new_n911));
  NAND2_X1  g486(.A1(G299), .A2(KEYINPUT107), .ZN(new_n912));
  OR2_X1    g487(.A1(G299), .A2(KEYINPUT107), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n619), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n629), .A2(KEYINPUT107), .A3(G299), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(KEYINPUT41), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n914), .A2(new_n921), .A3(new_n915), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT108), .B1(new_n917), .B2(new_n921), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n918), .B1(new_n925), .B2(new_n911), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n910), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n910), .A2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n855), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n929), .B1(G868), .B2(new_n930), .ZN(G295));
  OAI21_X1  g506(.A(new_n929), .B1(G868), .B2(new_n930), .ZN(G331));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n856), .A2(G171), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n856), .A2(G171), .ZN(new_n935));
  OR3_X1    g510(.A1(new_n934), .A2(new_n935), .A3(G286), .ZN(new_n936));
  OAI21_X1  g511(.A(G286), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n923), .B2(new_n924), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n916), .B1(new_n936), .B2(new_n937), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n908), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n920), .A2(new_n922), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n940), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n896), .B1(new_n945), .B2(new_n908), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n939), .A2(new_n941), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n909), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n949), .A2(new_n942), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n933), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(G37), .B1(new_n948), .B2(new_n909), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n950), .B1(new_n954), .B2(new_n942), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n943), .A2(new_n946), .A3(KEYINPUT43), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n953), .B1(new_n957), .B2(new_n933), .ZN(G397));
  NOR2_X1   g533(.A1(new_n875), .A2(G1384), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n475), .A2(G40), .A3(new_n484), .A4(new_n476), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G1996), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(new_n798), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n963), .B(KEYINPUT110), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n755), .B(new_n757), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n799), .A2(new_n965), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n967), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n730), .B(new_n734), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(G290), .B(G1986), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n964), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n959), .A2(new_n962), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(G2067), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n875), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n529), .B1(new_n528), .B2(new_n531), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n982), .A2(new_n983), .A3(G1384), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n962), .B(new_n981), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n979), .B1(new_n986), .B2(new_n762), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(new_n629), .ZN(new_n988));
  INV_X1    g563(.A(new_n521), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n528), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n961), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n523), .A2(new_n991), .A3(new_n532), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n993), .B1(KEYINPUT50), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n807), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(G1384), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n962), .B1(new_n875), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n994), .B2(new_n997), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT56), .B(G2072), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n996), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n582), .A2(new_n591), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n582), .A2(KEYINPUT114), .A3(new_n591), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n586), .A3(new_n1008), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT113), .B(KEYINPUT57), .Z(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT115), .B1(G299), .B2(new_n1012), .ZN(new_n1013));
  OR3_X1    g588(.A1(G299), .A2(KEYINPUT115), .A3(new_n1012), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n988), .B1(new_n1004), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1004), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n996), .A2(KEYINPUT116), .A3(new_n1003), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1020), .A3(new_n1016), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n987), .A2(KEYINPUT60), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT60), .ZN(new_n1024));
  AOI211_X1 g599(.A(new_n1024), .B(new_n979), .C1(new_n986), .C2(new_n762), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n619), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n986), .A2(new_n762), .ZN(new_n1028));
  INV_X1    g603(.A(new_n979), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(KEYINPUT60), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(KEYINPUT118), .A3(new_n629), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1023), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT61), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n996), .A2(new_n1003), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n1015), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1021), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1016), .A2(new_n1004), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1015), .B1(new_n996), .B2(new_n1003), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1035), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n572), .A2(KEYINPUT117), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1001), .A2(new_n965), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT58), .B(G1341), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n959), .B2(new_n962), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1042), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT59), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(new_n1042), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1038), .A2(new_n1041), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1022), .B1(new_n1034), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n1053));
  AOI211_X1 g628(.A(new_n1053), .B(KEYINPUT53), .C1(new_n1001), .C2(new_n770), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1000), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n770), .B(new_n1055), .C1(new_n984), .C2(KEYINPUT45), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT122), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n986), .A2(new_n812), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n961), .B1(new_n992), .B2(new_n997), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n523), .A2(new_n532), .A3(new_n998), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n770), .A3(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1063), .A2(KEYINPUT121), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1061), .A2(new_n1062), .A3(new_n1065), .A4(new_n770), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT53), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1060), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G171), .B1(new_n1059), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT123), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1071), .B(G171), .C1(new_n1059), .C2(new_n1068), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1053), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1056), .A2(KEYINPUT122), .A3(new_n1057), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n473), .A2(KEYINPUT53), .A3(G40), .A4(new_n770), .ZN(new_n1077));
  INV_X1    g652(.A(new_n484), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(KEYINPUT124), .B2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g654(.A(new_n1079), .B1(KEYINPUT124), .B2(new_n1078), .C1(new_n875), .C2(new_n999), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(new_n960), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n986), .B2(new_n812), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1076), .A2(G301), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1070), .A2(new_n1072), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G8), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n980), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n961), .A2(G2084), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1966), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1062), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n962), .B1(new_n959), .B2(KEYINPUT45), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1087), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(G286), .A2(G8), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT119), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT120), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(new_n1096), .B(KEYINPUT119), .Z(new_n1099));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1088), .A2(new_n1089), .B1(new_n1101), .B2(new_n1091), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1099), .B(new_n1100), .C1(new_n1102), .C2(new_n1087), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1098), .A2(new_n1103), .A3(KEYINPUT51), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT120), .B(new_n1106), .C1(new_n1095), .C2(new_n1097), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1066), .A2(KEYINPUT53), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1063), .A2(KEYINPUT121), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1109), .A2(new_n1110), .B1(new_n812), .B2(new_n986), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1076), .A2(new_n1111), .A3(G301), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1082), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1112), .A2(new_n1114), .A3(KEYINPUT54), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n978), .A2(G8), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(G1976), .B2(new_n718), .ZN(new_n1117));
  INV_X1    g692(.A(G1976), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT52), .B1(G288), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(G305), .A2(G1981), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n602), .B1(new_n604), .B2(new_n589), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G1981), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT49), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1121), .A2(KEYINPUT49), .A3(new_n1123), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1120), .B1(new_n1116), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1117), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT111), .B(G2090), .Z(new_n1133));
  NOR2_X1   g708(.A1(new_n995), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1001), .A2(G1971), .ZN(new_n1135));
  OAI21_X1  g710(.A(G8), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(G303), .A2(G8), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT55), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1138), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n986), .A2(new_n1133), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1140), .B(G8), .C1(new_n1141), .C2(new_n1135), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1132), .A2(new_n1139), .A3(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1108), .A2(new_n1115), .A3(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1052), .A2(new_n1086), .A3(new_n1144), .ZN(new_n1145));
  OAI221_X1 g720(.A(new_n1120), .B1(new_n1130), .B2(new_n1117), .C1(new_n1116), .C2(new_n1128), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1121), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n718), .A2(new_n1118), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT112), .Z(new_n1149));
  AOI21_X1  g724(.A(new_n1147), .B1(new_n1149), .B2(new_n1128), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1146), .A2(new_n1142), .B1(new_n1150), .B2(new_n1116), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1102), .A2(new_n1087), .A3(G286), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1132), .A2(new_n1139), .A3(new_n1142), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1152), .A2(KEYINPUT63), .ZN(new_n1156));
  OAI21_X1  g731(.A(G8), .B1(new_n1141), .B2(new_n1135), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1138), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1156), .A2(new_n1142), .A3(new_n1132), .A4(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1151), .B1(new_n1155), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1104), .A2(new_n1162), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1143), .A3(new_n1163), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1108), .A2(KEYINPUT62), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1160), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n977), .B1(new_n1145), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT46), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n966), .A2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT125), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n968), .B1(new_n798), .B2(new_n969), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1168), .B2(new_n966), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1173), .A2(KEYINPUT47), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(KEYINPUT47), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1174), .A2(KEYINPUT126), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT126), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1177));
  INV_X1    g752(.A(new_n731), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n972), .A2(new_n1178), .A3(new_n734), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n755), .A2(new_n757), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n968), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n963), .A2(G1986), .A3(G290), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT127), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT48), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1181), .B1(new_n975), .B2(new_n1184), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1176), .A2(new_n1177), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1167), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g762(.A(G227), .ZN(new_n1189));
  OAI211_X1 g763(.A(G319), .B(new_n1189), .C1(new_n663), .C2(new_n664), .ZN(new_n1190));
  AOI21_X1  g764(.A(new_n1190), .B1(new_n696), .B2(new_n700), .ZN(new_n1191));
  OAI211_X1 g765(.A(new_n897), .B(new_n1191), .C1(new_n955), .C2(new_n956), .ZN(G225));
  INV_X1    g766(.A(G225), .ZN(G308));
endmodule


