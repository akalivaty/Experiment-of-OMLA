//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n463), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT69), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(G126), .B2(new_n480), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n464), .B2(new_n465), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(KEYINPUT70), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(new_n492), .C1(new_n465), .C2(new_n464), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n489), .A2(new_n495), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G50), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n502), .A2(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n511), .A2(new_n514), .ZN(G166));
  NAND3_X1  g090(.A1(new_n506), .A2(G89), .A3(new_n508), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT7), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n517), .B(KEYINPUT72), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  OAI211_X1 g098(.A(KEYINPUT73), .B(new_n516), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n507), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n525), .A2(G51), .B1(new_n508), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(new_n520), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT73), .B1(new_n531), .B2(new_n516), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT74), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n516), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n536), .A2(new_n537), .A3(new_n524), .A4(new_n527), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n533), .A2(new_n538), .ZN(G168));
  AOI22_X1  g114(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n513), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n543), .A2(new_n507), .B1(new_n509), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(G171));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n547), .A2(new_n507), .B1(new_n509), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n513), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(new_n509), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n559), .A2(KEYINPUT76), .A3(G91), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n509), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  XOR2_X1   g139(.A(KEYINPUT5), .B(G543), .Z(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n560), .A2(new_n563), .B1(G651), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OR3_X1    g144(.A1(new_n507), .A2(KEYINPUT9), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT9), .B1(new_n507), .B2(new_n569), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  OAI21_X1  g151(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n577));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  INV_X1    g153(.A(G49), .ZN(new_n579));
  OAI221_X1 g154(.A(new_n577), .B1(new_n509), .B2(new_n578), .C1(new_n579), .C2(new_n507), .ZN(G288));
  INV_X1    g155(.A(G48), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n581), .A2(new_n507), .B1(new_n509), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n508), .A2(G61), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT77), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n513), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n588), .A2(KEYINPUT78), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(KEYINPUT78), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n584), .B1(new_n589), .B2(new_n590), .ZN(G305));
  XNOR2_X1  g166(.A(KEYINPUT79), .B(G85), .ZN(new_n592));
  AOI22_X1  g167(.A1(G47), .A2(new_n525), .B1(new_n559), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n513), .B2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n509), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G54), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n507), .A2(new_n600), .B1(new_n601), .B2(new_n513), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI221_X1 g179(.A(KEYINPUT80), .B1(new_n601), .B2(new_n513), .C1(new_n600), .C2(new_n507), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n596), .B1(new_n608), .B2(G868), .ZN(G321));
  XNOR2_X1  g184(.A(G321), .B(KEYINPUT81), .ZN(G284));
  NOR2_X1   g185(.A1(G299), .A2(G868), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g187(.A(new_n611), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n608), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n608), .A2(new_n614), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT82), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(new_n552), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(G282));
  INV_X1    g198(.A(new_n621), .ZN(G323));
  NAND2_X1  g199(.A1(new_n476), .A2(new_n477), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n470), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n478), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n480), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n463), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n631), .A3(new_n637), .ZN(G156));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT84), .Z(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n643), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT85), .Z(new_n658));
  NOR2_X1   g233(.A1(G2072), .A2(G2078), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n442), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n656), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(KEYINPUT17), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n656), .B(new_n657), .C1(new_n442), .C2(new_n659), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n658), .A2(new_n656), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n666), .B1(new_n662), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT87), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n673), .A2(new_n674), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n681), .A2(new_n677), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT88), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n675), .A2(new_n681), .A3(new_n677), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G229));
  NOR2_X1   g266(.A1(G16), .A2(G21), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G168), .B2(G16), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT92), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT93), .B(G1966), .Z(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NOR2_X1   g275(.A1(G171), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G5), .B2(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(G1961), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n705), .A2(G32), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT26), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n478), .A2(G141), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n480), .A2(G129), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n470), .A2(G105), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n708), .A2(new_n709), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(G29), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT27), .B(G1996), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n702), .B2(new_n703), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n705), .A2(G33), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n625), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(new_n463), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT25), .ZN(new_n720));
  NAND2_X1  g295(.A1(G103), .A2(G2104), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G2105), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n463), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n478), .A2(G139), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n717), .B1(new_n725), .B2(new_n705), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(G2072), .Z(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT30), .B(G28), .ZN(new_n728));
  OR2_X1    g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  NAND2_X1  g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n728), .A2(new_n705), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n636), .B2(new_n705), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n713), .B2(new_n714), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n704), .A2(new_n716), .A3(new_n727), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n705), .A2(G27), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G164), .B2(new_n705), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2078), .ZN(new_n737));
  INV_X1    g312(.A(G34), .ZN(new_n738));
  AOI21_X1  g313(.A(G29), .B1(new_n738), .B2(KEYINPUT24), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(KEYINPUT24), .B2(new_n738), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n474), .B2(new_n705), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  OR3_X1    g319(.A1(new_n737), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n699), .A2(new_n734), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n697), .A2(new_n698), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n746), .A2(KEYINPUT94), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n705), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n705), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2090), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n608), .A2(G16), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G4), .B2(G16), .ZN(new_n754));
  INV_X1    g329(.A(G1348), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  AOI21_X1  g332(.A(KEYINPUT23), .B1(new_n700), .B2(G20), .ZN(new_n758));
  AND3_X1   g333(.A1(new_n700), .A2(KEYINPUT23), .A3(G20), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n758), .B(new_n759), .C1(G299), .C2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT95), .B(G1956), .Z(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n700), .A2(G19), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n552), .B2(new_n700), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1341), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n705), .A2(G26), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT28), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n478), .A2(G140), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n480), .A2(G128), .ZN(new_n770));
  OR2_X1    g345(.A1(G104), .A2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n771), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n772));
  AND3_X1   g347(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(new_n705), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n766), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n756), .A2(new_n757), .A3(new_n763), .A4(new_n776), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n752), .B(new_n777), .C1(new_n762), .C2(new_n760), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n748), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT96), .ZN(new_n781));
  AOI21_X1  g356(.A(KEYINPUT94), .B1(new_n746), .B2(new_n747), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(KEYINPUT96), .B1(new_n779), .B2(new_n782), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n700), .A2(G6), .ZN(new_n786));
  INV_X1    g361(.A(G305), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n700), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT90), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT32), .B(G1981), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n789), .A2(new_n791), .ZN(new_n793));
  MUX2_X1   g368(.A(G23), .B(G288), .S(G16), .Z(new_n794));
  XOR2_X1   g369(.A(KEYINPUT33), .B(G1976), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n700), .A2(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G166), .B2(new_n700), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1971), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n792), .A2(new_n793), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(KEYINPUT34), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT34), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n792), .A2(new_n793), .A3(new_n803), .A4(new_n800), .ZN(new_n804));
  MUX2_X1   g379(.A(G24), .B(G290), .S(G16), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1986), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n705), .A2(G25), .ZN(new_n807));
  NOR2_X1   g382(.A1(G95), .A2(G2105), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT89), .Z(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(new_n463), .B2(G107), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n478), .A2(G131), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n480), .A2(G119), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n807), .B1(new_n816), .B2(new_n705), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n806), .A2(new_n820), .ZN(new_n821));
  AND3_X1   g396(.A1(new_n804), .A2(KEYINPUT91), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(KEYINPUT91), .B1(new_n804), .B2(new_n821), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n802), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(new_n802), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n784), .A2(new_n785), .B1(new_n825), .B2(new_n827), .ZN(G311));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n827), .ZN(new_n829));
  INV_X1    g404(.A(new_n785), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n779), .A2(KEYINPUT96), .A3(new_n782), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(G150));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n614), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n506), .A2(G55), .A3(G543), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT98), .B(G93), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n835), .B(KEYINPUT99), .C1(new_n509), .C2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  OR3_X1    g413(.A1(new_n565), .A2(new_n505), .A3(new_n836), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT99), .B1(new_n839), .B2(new_n835), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n513), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(KEYINPUT97), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n841), .A2(new_n844), .A3(new_n513), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n838), .A2(new_n840), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n619), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n842), .B(KEYINPUT97), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(new_n552), .C1(new_n840), .C2(new_n838), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n834), .B(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n852), .A2(new_n853), .A3(G860), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n846), .A2(G860), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  NAND2_X1  g432(.A1(new_n478), .A2(G142), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT101), .Z(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  INV_X1    g435(.A(G118), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(G2105), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(G130), .B2(new_n480), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n627), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n725), .A2(KEYINPUT100), .ZN(new_n868));
  INV_X1    g443(.A(new_n712), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n867), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n500), .B(new_n773), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n816), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n871), .B(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n474), .B(new_n636), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G162), .ZN(new_n877));
  AOI21_X1  g452(.A(G37), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n871), .B(new_n873), .ZN(new_n879));
  INV_X1    g454(.A(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g458(.A(new_n617), .B(new_n850), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n599), .A2(new_n606), .A3(new_n568), .A4(new_n572), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI22_X1  g461(.A1(new_n606), .A2(new_n599), .B1(new_n568), .B2(new_n572), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT41), .B1(new_n886), .B2(new_n887), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n607), .A2(G299), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n892), .A3(new_n885), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n889), .B1(new_n884), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n787), .A2(G290), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G166), .B(G288), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n787), .A2(G290), .ZN(new_n900));
  OR3_X1    g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n898), .B2(new_n900), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(KEYINPUT103), .B2(KEYINPUT42), .ZN(new_n904));
  NAND2_X1  g479(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n904), .B(new_n905), .Z(new_n906));
  AND2_X1   g481(.A1(new_n896), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n896), .A2(new_n906), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n846), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(G868), .B2(new_n910), .ZN(G295));
  OAI21_X1  g486(.A(new_n909), .B1(G868), .B2(new_n910), .ZN(G331));
  NAND3_X1  g487(.A1(new_n888), .A2(KEYINPUT104), .A3(new_n892), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n890), .A2(new_n914), .A3(new_n893), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n533), .A2(new_n538), .A3(G301), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(G301), .B1(new_n533), .B2(new_n538), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n917), .A2(new_n918), .A3(new_n850), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n847), .A2(new_n849), .ZN(new_n920));
  NAND2_X1  g495(.A1(G168), .A2(G171), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n916), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n913), .B(new_n915), .C1(new_n919), .C2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n850), .B1(new_n917), .B2(new_n918), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n921), .A2(new_n920), .A3(new_n916), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n888), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n903), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT105), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n924), .A2(new_n925), .A3(new_n888), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n924), .A2(new_n925), .B1(new_n893), .B2(new_n890), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(G37), .B1(new_n938), .B2(new_n903), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n933), .A2(new_n934), .A3(new_n935), .A4(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n931), .B1(new_n927), .B2(new_n928), .ZN(new_n941));
  AOI211_X1 g516(.A(KEYINPUT105), .B(new_n903), .C1(new_n923), .C2(new_n926), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n935), .B(new_n939), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT106), .ZN(new_n944));
  INV_X1    g519(.A(new_n939), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n938), .A2(new_n903), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n940), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n933), .A2(KEYINPUT43), .A3(new_n939), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n935), .B1(new_n945), .B2(new_n946), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT44), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(new_n954), .ZN(G397));
  INV_X1    g530(.A(G2067), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n773), .B(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT108), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(new_n712), .ZN(new_n959));
  INV_X1    g534(.A(G40), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n468), .A2(new_n472), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  OAI211_X1 g538(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n964));
  INV_X1    g539(.A(new_n486), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(G114), .B2(new_n463), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n499), .A2(new_n964), .A3(new_n966), .A4(new_n497), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n463), .A2(G138), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n476), .B2(new_n477), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT4), .B1(new_n969), .B2(KEYINPUT71), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n963), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n959), .A2(new_n962), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n974), .B1(G1996), .B2(new_n958), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n973), .A2(new_n962), .ZN(new_n976));
  INV_X1    g551(.A(G1996), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n975), .B1(new_n712), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n815), .B(new_n819), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  NOR2_X1   g557(.A1(G290), .A2(G1986), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n976), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n962), .A2(G2090), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n987), .B(new_n963), .C1(new_n967), .C2(new_n970), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n987), .B1(new_n500), .B2(new_n963), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n971), .A2(KEYINPUT109), .A3(KEYINPUT50), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT110), .B(new_n986), .C1(new_n992), .C2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1971), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n960), .B1(new_n971), .B2(new_n972), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n473), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n996), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n971), .A2(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1003), .A2(new_n989), .A3(new_n988), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n993), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT110), .B1(new_n1005), .B2(new_n986), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT111), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n986), .B1(new_n992), .B2(new_n994), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n1001), .A4(new_n995), .ZN(new_n1012));
  INV_X1    g587(.A(G8), .ZN(new_n1013));
  NOR2_X1   g588(.A1(G166), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n1015));
  OR2_X1    g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(KEYINPUT112), .B2(KEYINPUT55), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1007), .A2(new_n1012), .A3(G8), .A4(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n971), .A2(new_n962), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(new_n1013), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1021), .B(new_n1023), .C1(new_n1022), .C2(G288), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n500), .A2(new_n963), .A3(new_n961), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1025), .B(G8), .C1(new_n1022), .C2(G288), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  INV_X1    g602(.A(G1981), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n584), .B(new_n1028), .C1(new_n589), .C2(new_n590), .ZN(new_n1029));
  OAI21_X1  g604(.A(G1981), .B1(new_n583), .B2(new_n588), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT113), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1021), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1024), .B(new_n1027), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n988), .B1(new_n991), .B2(KEYINPUT114), .ZN(new_n1037));
  OR3_X1    g612(.A1(new_n971), .A2(KEYINPUT114), .A3(KEYINPUT50), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n961), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1001), .B1(new_n1039), .B2(G2090), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G8), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1018), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1036), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1019), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT123), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT123), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1019), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n999), .A2(new_n473), .ZN(new_n1048));
  INV_X1    g623(.A(G2078), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n997), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT45), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n971), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n972), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n500), .A2(new_n963), .A3(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1051), .A2(G2078), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1054), .A2(new_n961), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n962), .B1(new_n1004), .B2(new_n993), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1052), .B(new_n1058), .C1(G1961), .C2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g635(.A(G171), .B(KEYINPUT54), .Z(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1005), .A2(new_n961), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n703), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT121), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT121), .B1(new_n469), .B2(new_n471), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1065), .A2(new_n1066), .A3(new_n468), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n997), .A2(new_n1067), .A3(KEYINPUT122), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT122), .B1(new_n997), .B2(new_n1067), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n999), .B(new_n1057), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1061), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1064), .A2(new_n1070), .A3(new_n1052), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1062), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1005), .A2(new_n742), .A3(new_n961), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n961), .B1(new_n971), .B2(new_n972), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT45), .B1(new_n500), .B2(new_n963), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n698), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT115), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(new_n698), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1074), .A2(G168), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1080), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1054), .A2(new_n961), .A3(new_n1056), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1079), .B1(new_n1084), .B2(new_n698), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(G168), .B1(new_n1086), .B2(new_n1074), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT51), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1081), .A2(new_n1089), .A3(G8), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1073), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1045), .A2(new_n1047), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1045), .A2(new_n1091), .A3(KEYINPUT124), .A4(new_n1047), .ZN(new_n1095));
  INV_X1    g670(.A(G1956), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1039), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1048), .A2(new_n997), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(G299), .B(KEYINPUT57), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(new_n607), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1063), .A2(new_n755), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1025), .A2(KEYINPUT116), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1025), .A2(KEYINPUT116), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n956), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT117), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1108), .B(KEYINPUT117), .C1(new_n1059), .C2(G1348), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1103), .A2(new_n1112), .B1(new_n1101), .B2(new_n1100), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1109), .A2(new_n1111), .A3(KEYINPUT60), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT60), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n608), .ZN(new_n1116));
  OAI211_X1 g691(.A(KEYINPUT60), .B(new_n607), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n997), .A2(new_n977), .A3(new_n473), .A4(new_n999), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT118), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1107), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT58), .B(G1341), .Z(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(new_n1105), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1048), .A2(new_n1125), .A3(new_n977), .A4(new_n997), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1121), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1119), .B1(new_n1127), .B2(new_n552), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1127), .A2(new_n1119), .A3(new_n552), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(KEYINPUT59), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1127), .A2(new_n1119), .A3(new_n552), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(new_n1128), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1100), .A2(KEYINPUT120), .A3(new_n1101), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1101), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1136), .A2(new_n1097), .A3(KEYINPUT120), .A4(new_n1099), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1135), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1131), .B(new_n1134), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1113), .B1(new_n1118), .B2(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1094), .A2(new_n1095), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1144), .A2(G1976), .A3(G288), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1029), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1021), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1019), .B2(new_n1036), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1150));
  AOI211_X1 g725(.A(G2084), .B(new_n962), .C1(new_n1004), .C2(new_n993), .ZN(new_n1151));
  OAI211_X1 g726(.A(G8), .B(G168), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1149), .B1(new_n1044), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1007), .A2(G8), .A3(new_n1012), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1042), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1152), .A2(new_n1149), .A3(new_n1036), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(new_n1019), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1148), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1081), .A2(new_n1089), .A3(G8), .ZN(new_n1159));
  OAI21_X1  g734(.A(G286), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1160), .A2(G8), .A3(new_n1081), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1159), .B1(KEYINPUT51), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT125), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1060), .A2(G171), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(KEYINPUT62), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1164), .A2(new_n1166), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1158), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n985), .B1(new_n1143), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n983), .A2(new_n976), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT48), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n981), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT46), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n978), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT126), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n978), .A2(new_n1177), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n974), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT47), .Z(new_n1182));
  NAND2_X1  g757(.A1(new_n1176), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n773), .A2(new_n956), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n816), .A2(new_n818), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1184), .B1(new_n979), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1183), .B1(new_n976), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1173), .A2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g763(.A(G319), .B1(new_n653), .B2(new_n654), .ZN(new_n1190));
  OR2_X1    g764(.A1(new_n1190), .A2(G227), .ZN(new_n1191));
  NOR2_X1   g765(.A1(G229), .A2(new_n1191), .ZN(new_n1192));
  AND3_X1   g766(.A1(new_n948), .A2(new_n882), .A3(new_n1192), .ZN(G308));
  NAND3_X1  g767(.A1(new_n948), .A2(new_n882), .A3(new_n1192), .ZN(G225));
endmodule


