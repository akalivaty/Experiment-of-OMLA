

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n528), .A2(n527), .ZN(G164) );
  NAND2_X2 U553 ( .A1(n796), .A2(n696), .ZN(n738) );
  NOR2_X1 U554 ( .A1(G164), .A2(G1384), .ZN(n796) );
  NOR2_X2 U555 ( .A1(n553), .A2(n552), .ZN(G160) );
  INV_X1 U556 ( .A(KEYINPUT31), .ZN(n708) );
  INV_X1 U557 ( .A(n950), .ZN(n763) );
  AND2_X1 U558 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X2 U559 ( .A(KEYINPUT66), .B(G2104), .Z(n523) );
  NAND2_X1 U560 ( .A1(n523), .A2(G2105), .ZN(n518) );
  XNOR2_X2 U561 ( .A(n518), .B(KEYINPUT67), .ZN(n892) );
  NAND2_X1 U562 ( .A1(n892), .A2(G126), .ZN(n521) );
  AND2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U564 ( .A1(n891), .A2(G114), .ZN(n519) );
  XOR2_X1 U565 ( .A(KEYINPUT95), .B(n519), .Z(n520) );
  NAND2_X1 U566 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U567 ( .A(n522), .B(KEYINPUT96), .ZN(n528) );
  NOR2_X4 U568 ( .A1(G2105), .A2(n523), .ZN(n896) );
  NAND2_X1 U569 ( .A1(n896), .A2(G102), .ZN(n526) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  XOR2_X1 U571 ( .A(KEYINPUT17), .B(n524), .Z(n895) );
  NAND2_X1 U572 ( .A1(n895), .A2(G138), .ZN(n525) );
  NAND2_X1 U573 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U574 ( .A(G651), .B(KEYINPUT70), .Z(n537) );
  NOR2_X1 U575 ( .A1(G543), .A2(n537), .ZN(n529) );
  XOR2_X1 U576 ( .A(KEYINPUT1), .B(n529), .Z(n654) );
  NAND2_X1 U577 ( .A1(G63), .A2(n654), .ZN(n533) );
  XNOR2_X1 U578 ( .A(G543), .B(KEYINPUT0), .ZN(n530) );
  XNOR2_X1 U579 ( .A(n530), .B(KEYINPUT69), .ZN(n646) );
  NOR2_X1 U580 ( .A1(G651), .A2(n646), .ZN(n531) );
  XOR2_X1 U581 ( .A(KEYINPUT65), .B(n531), .Z(n655) );
  NAND2_X1 U582 ( .A1(G51), .A2(n655), .ZN(n532) );
  NAND2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U584 ( .A(KEYINPUT6), .B(n534), .ZN(n543) );
  NOR2_X1 U585 ( .A1(G651), .A2(G543), .ZN(n663) );
  NAND2_X1 U586 ( .A1(G89), .A2(n663), .ZN(n535) );
  XNOR2_X1 U587 ( .A(n535), .B(KEYINPUT4), .ZN(n536) );
  XNOR2_X1 U588 ( .A(n536), .B(KEYINPUT78), .ZN(n539) );
  NOR2_X1 U589 ( .A1(n646), .A2(n537), .ZN(n658) );
  NAND2_X1 U590 ( .A1(G76), .A2(n658), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U592 ( .A(KEYINPUT79), .B(n540), .ZN(n541) );
  XNOR2_X1 U593 ( .A(KEYINPUT5), .B(n541), .ZN(n542) );
  NOR2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U595 ( .A(KEYINPUT7), .B(n544), .Z(G168) );
  NAND2_X1 U596 ( .A1(G101), .A2(n896), .ZN(n546) );
  INV_X1 U597 ( .A(KEYINPUT68), .ZN(n545) );
  XNOR2_X1 U598 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U599 ( .A(n547), .B(KEYINPUT23), .ZN(n549) );
  NAND2_X1 U600 ( .A1(G113), .A2(n891), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U602 ( .A1(G125), .A2(n892), .ZN(n551) );
  NAND2_X1 U603 ( .A1(G137), .A2(n895), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U605 ( .A(G2438), .B(G2454), .Z(n555) );
  XNOR2_X1 U606 ( .A(G2435), .B(G2430), .ZN(n554) );
  XNOR2_X1 U607 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U608 ( .A(n556), .B(G2427), .Z(n558) );
  XNOR2_X1 U609 ( .A(G1341), .B(G1348), .ZN(n557) );
  XNOR2_X1 U610 ( .A(n558), .B(n557), .ZN(n562) );
  XOR2_X1 U611 ( .A(G2443), .B(G2446), .Z(n560) );
  XNOR2_X1 U612 ( .A(KEYINPUT110), .B(G2451), .ZN(n559) );
  XNOR2_X1 U613 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U614 ( .A(n562), .B(n561), .Z(n563) );
  AND2_X1 U615 ( .A1(G14), .A2(n563), .ZN(G401) );
  NAND2_X1 U616 ( .A1(G64), .A2(n654), .ZN(n565) );
  NAND2_X1 U617 ( .A1(G52), .A2(n655), .ZN(n564) );
  NAND2_X1 U618 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U619 ( .A1(G77), .A2(n658), .ZN(n567) );
  NAND2_X1 U620 ( .A1(G90), .A2(n663), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U622 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U623 ( .A1(n570), .A2(n569), .ZN(G171) );
  AND2_X1 U624 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U625 ( .A(G57), .ZN(G237) );
  INV_X1 U626 ( .A(G132), .ZN(G219) );
  INV_X1 U627 ( .A(G82), .ZN(G220) );
  NAND2_X1 U628 ( .A1(G62), .A2(n654), .ZN(n572) );
  NAND2_X1 U629 ( .A1(G50), .A2(n655), .ZN(n571) );
  NAND2_X1 U630 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U631 ( .A(KEYINPUT86), .B(n573), .Z(n579) );
  NAND2_X1 U632 ( .A1(n663), .A2(G88), .ZN(n574) );
  XOR2_X1 U633 ( .A(KEYINPUT87), .B(n574), .Z(n576) );
  NAND2_X1 U634 ( .A1(n658), .A2(G75), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U636 ( .A(KEYINPUT88), .B(n577), .Z(n578) );
  NAND2_X1 U637 ( .A1(n579), .A2(n578), .ZN(G303) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U640 ( .A(n580), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U641 ( .A(G223), .ZN(n837) );
  NAND2_X1 U642 ( .A1(n837), .A2(G567), .ZN(n581) );
  XNOR2_X1 U643 ( .A(n581), .B(KEYINPUT11), .ZN(n582) );
  XNOR2_X1 U644 ( .A(KEYINPUT73), .B(n582), .ZN(G234) );
  NAND2_X1 U645 ( .A1(G56), .A2(n654), .ZN(n583) );
  XOR2_X1 U646 ( .A(KEYINPUT14), .B(n583), .Z(n589) );
  NAND2_X1 U647 ( .A1(n663), .A2(G81), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G68), .A2(n658), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT13), .B(n587), .Z(n588) );
  NOR2_X1 U652 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U653 ( .A1(n655), .A2(G43), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n591), .A2(n590), .ZN(n946) );
  INV_X1 U655 ( .A(G860), .ZN(n614) );
  OR2_X1 U656 ( .A1(n946), .A2(n614), .ZN(G153) );
  XOR2_X1 U657 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U659 ( .A1(G79), .A2(n658), .ZN(n592) );
  XNOR2_X1 U660 ( .A(n592), .B(KEYINPUT76), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G66), .A2(n654), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G54), .A2(n655), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G92), .A2(n663), .ZN(n595) );
  XNOR2_X1 U665 ( .A(KEYINPUT75), .B(n595), .ZN(n596) );
  NOR2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n601) );
  XOR2_X1 U668 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n600) );
  XNOR2_X1 U669 ( .A(n601), .B(n600), .ZN(n909) );
  INV_X1 U670 ( .A(n909), .ZN(n963) );
  INV_X1 U671 ( .A(G868), .ZN(n677) );
  NAND2_X1 U672 ( .A1(n963), .A2(n677), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U674 ( .A1(G78), .A2(n658), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G91), .A2(n663), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U677 ( .A1(n655), .A2(G53), .ZN(n606) );
  XOR2_X1 U678 ( .A(KEYINPUT72), .B(n606), .Z(n607) );
  NOR2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n654), .A2(G65), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n610), .A2(n609), .ZN(G299) );
  NOR2_X1 U682 ( .A1(G286), .A2(n677), .ZN(n612) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U685 ( .A(KEYINPUT80), .B(n613), .ZN(G297) );
  NAND2_X1 U686 ( .A1(n614), .A2(G559), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n615), .A2(n909), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U689 ( .A1(G868), .A2(n946), .ZN(n619) );
  NAND2_X1 U690 ( .A1(G868), .A2(n909), .ZN(n617) );
  NOR2_X1 U691 ( .A1(G559), .A2(n617), .ZN(n618) );
  NOR2_X1 U692 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U693 ( .A1(G111), .A2(n891), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G135), .A2(n895), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n627) );
  NAND2_X1 U696 ( .A1(G123), .A2(n892), .ZN(n622) );
  XOR2_X1 U697 ( .A(KEYINPUT18), .B(n622), .Z(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(KEYINPUT81), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G99), .A2(n896), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n977) );
  XNOR2_X1 U702 ( .A(n977), .B(G2096), .ZN(n629) );
  INV_X1 U703 ( .A(G2100), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(G156) );
  NAND2_X1 U705 ( .A1(G80), .A2(n658), .ZN(n631) );
  NAND2_X1 U706 ( .A1(G67), .A2(n654), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n663), .A2(G93), .ZN(n632) );
  XOR2_X1 U709 ( .A(KEYINPUT82), .B(n632), .Z(n633) );
  NOR2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n655), .A2(G55), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n676) );
  NAND2_X1 U713 ( .A1(n909), .A2(G559), .ZN(n674) );
  XNOR2_X1 U714 ( .A(n946), .B(n674), .ZN(n637) );
  NOR2_X1 U715 ( .A1(G860), .A2(n637), .ZN(n638) );
  XOR2_X1 U716 ( .A(n676), .B(n638), .Z(G145) );
  NAND2_X1 U717 ( .A1(G72), .A2(n658), .ZN(n640) );
  NAND2_X1 U718 ( .A1(G47), .A2(n655), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G60), .A2(n654), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G85), .A2(n663), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n645), .B(KEYINPUT71), .ZN(G290) );
  INV_X1 U725 ( .A(G303), .ZN(G166) );
  NAND2_X1 U726 ( .A1(n646), .A2(G87), .ZN(n647) );
  XNOR2_X1 U727 ( .A(KEYINPUT84), .B(n647), .ZN(n653) );
  NAND2_X1 U728 ( .A1(G49), .A2(n655), .ZN(n649) );
  NAND2_X1 U729 ( .A1(G74), .A2(G651), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U731 ( .A1(n654), .A2(n650), .ZN(n651) );
  XOR2_X1 U732 ( .A(KEYINPUT83), .B(n651), .Z(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(G288) );
  NAND2_X1 U734 ( .A1(G61), .A2(n654), .ZN(n657) );
  NAND2_X1 U735 ( .A1(G48), .A2(n655), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n662) );
  XOR2_X1 U737 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n660) );
  NAND2_X1 U738 ( .A1(n658), .A2(G73), .ZN(n659) );
  XOR2_X1 U739 ( .A(n660), .B(n659), .Z(n661) );
  NOR2_X1 U740 ( .A1(n662), .A2(n661), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n663), .A2(G86), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(G305) );
  INV_X1 U743 ( .A(G299), .ZN(n955) );
  XNOR2_X1 U744 ( .A(n955), .B(G290), .ZN(n671) );
  XNOR2_X1 U745 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n667) );
  XNOR2_X1 U746 ( .A(G288), .B(KEYINPUT19), .ZN(n666) );
  XNOR2_X1 U747 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U748 ( .A(G166), .B(n668), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n669), .B(n676), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n672), .B(G305), .ZN(n673) );
  XNOR2_X1 U752 ( .A(n673), .B(n946), .ZN(n908) );
  XNOR2_X1 U753 ( .A(n674), .B(n908), .ZN(n675) );
  NAND2_X1 U754 ( .A1(n675), .A2(G868), .ZN(n679) );
  NAND2_X1 U755 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U756 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n680) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n680), .Z(n681) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n681), .ZN(n682) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n682), .ZN(n683) );
  NAND2_X1 U761 ( .A1(n683), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U763 ( .A1(G661), .A2(G483), .ZN(n694) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n684) );
  XNOR2_X1 U765 ( .A(KEYINPUT22), .B(n684), .ZN(n685) );
  NAND2_X1 U766 ( .A1(n685), .A2(G96), .ZN(n686) );
  NOR2_X1 U767 ( .A1(n686), .A2(G218), .ZN(n687) );
  XNOR2_X1 U768 ( .A(n687), .B(KEYINPUT91), .ZN(n843) );
  NAND2_X1 U769 ( .A1(G2106), .A2(n843), .ZN(n688) );
  XNOR2_X1 U770 ( .A(n688), .B(KEYINPUT92), .ZN(n692) );
  NAND2_X1 U771 ( .A1(G69), .A2(G120), .ZN(n689) );
  NOR2_X1 U772 ( .A1(G237), .A2(n689), .ZN(n690) );
  NAND2_X1 U773 ( .A1(G108), .A2(n690), .ZN(n842) );
  NAND2_X1 U774 ( .A1(G567), .A2(n842), .ZN(n691) );
  NAND2_X1 U775 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U776 ( .A(KEYINPUT93), .B(n693), .Z(n845) );
  NOR2_X1 U777 ( .A1(n694), .A2(n845), .ZN(n695) );
  XNOR2_X1 U778 ( .A(n695), .B(KEYINPUT94), .ZN(n840) );
  NAND2_X1 U779 ( .A1(G36), .A2(n840), .ZN(G176) );
  NOR2_X1 U780 ( .A1(G1976), .A2(G288), .ZN(n949) );
  AND2_X1 U781 ( .A1(KEYINPUT33), .A2(n949), .ZN(n698) );
  NAND2_X1 U782 ( .A1(G160), .A2(G40), .ZN(n795) );
  INV_X1 U783 ( .A(n795), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n738), .A2(G8), .ZN(n697) );
  XOR2_X2 U785 ( .A(KEYINPUT100), .B(n697), .Z(n780) );
  NAND2_X1 U786 ( .A1(n698), .A2(n780), .ZN(n771) );
  OR2_X1 U787 ( .A1(G1981), .A2(G305), .ZN(n772) );
  NAND2_X1 U788 ( .A1(G1981), .A2(G305), .ZN(n699) );
  NAND2_X1 U789 ( .A1(n772), .A2(n699), .ZN(n943) );
  INV_X1 U790 ( .A(n780), .ZN(n764) );
  NOR2_X1 U791 ( .A1(n764), .A2(G1966), .ZN(n756) );
  NOR2_X1 U792 ( .A1(G2084), .A2(n738), .ZN(n752) );
  NOR2_X1 U793 ( .A1(n756), .A2(n752), .ZN(n700) );
  NAND2_X1 U794 ( .A1(G8), .A2(n700), .ZN(n701) );
  XNOR2_X1 U795 ( .A(n701), .B(KEYINPUT30), .ZN(n702) );
  NOR2_X1 U796 ( .A1(n702), .A2(G168), .ZN(n707) );
  XOR2_X1 U797 ( .A(G2078), .B(KEYINPUT25), .Z(n927) );
  NOR2_X1 U798 ( .A1(n927), .A2(n738), .ZN(n704) );
  INV_X1 U799 ( .A(n738), .ZN(n712) );
  NOR2_X1 U800 ( .A1(n712), .A2(G1961), .ZN(n703) );
  NOR2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U802 ( .A(KEYINPUT101), .B(n705), .ZN(n710) );
  NOR2_X1 U803 ( .A1(G171), .A2(n710), .ZN(n706) );
  NOR2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n709) );
  XNOR2_X1 U805 ( .A(n709), .B(n708), .ZN(n754) );
  NAND2_X1 U806 ( .A1(n710), .A2(G171), .ZN(n737) );
  NAND2_X1 U807 ( .A1(n712), .A2(G2072), .ZN(n711) );
  XNOR2_X1 U808 ( .A(n711), .B(KEYINPUT27), .ZN(n714) );
  INV_X1 U809 ( .A(G1956), .ZN(n1009) );
  NOR2_X1 U810 ( .A1(n1009), .A2(n712), .ZN(n713) );
  NOR2_X1 U811 ( .A1(n714), .A2(n713), .ZN(n717) );
  NOR2_X1 U812 ( .A1(n717), .A2(n955), .ZN(n716) );
  XOR2_X1 U813 ( .A(KEYINPUT28), .B(KEYINPUT102), .Z(n715) );
  XNOR2_X1 U814 ( .A(n716), .B(n715), .ZN(n734) );
  NAND2_X1 U815 ( .A1(n717), .A2(n955), .ZN(n732) );
  INV_X1 U816 ( .A(G1996), .ZN(n918) );
  NOR2_X1 U817 ( .A1(n738), .A2(n918), .ZN(n719) );
  XOR2_X1 U818 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n718) );
  XNOR2_X1 U819 ( .A(n719), .B(n718), .ZN(n721) );
  NAND2_X1 U820 ( .A1(n738), .A2(G1341), .ZN(n720) );
  NAND2_X1 U821 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U822 ( .A1(n946), .A2(n722), .ZN(n728) );
  NAND2_X1 U823 ( .A1(n909), .A2(n728), .ZN(n727) );
  INV_X1 U824 ( .A(G2067), .ZN(n924) );
  NOR2_X1 U825 ( .A1(n738), .A2(n924), .ZN(n723) );
  XNOR2_X1 U826 ( .A(n723), .B(KEYINPUT103), .ZN(n725) );
  NAND2_X1 U827 ( .A1(n738), .A2(G1348), .ZN(n724) );
  NAND2_X1 U828 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U829 ( .A1(n727), .A2(n726), .ZN(n730) );
  OR2_X1 U830 ( .A1(n909), .A2(n728), .ZN(n729) );
  NAND2_X1 U831 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U832 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U833 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U834 ( .A(KEYINPUT29), .B(n735), .Z(n736) );
  NAND2_X1 U835 ( .A1(n737), .A2(n736), .ZN(n753) );
  INV_X1 U836 ( .A(G8), .ZN(n744) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n738), .ZN(n739) );
  XNOR2_X1 U838 ( .A(n739), .B(KEYINPUT104), .ZN(n741) );
  NOR2_X1 U839 ( .A1(n764), .A2(G1971), .ZN(n740) );
  NOR2_X1 U840 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U841 ( .A1(n742), .A2(G303), .ZN(n743) );
  OR2_X1 U842 ( .A1(n744), .A2(n743), .ZN(n746) );
  AND2_X1 U843 ( .A1(n753), .A2(n746), .ZN(n745) );
  NAND2_X1 U844 ( .A1(n754), .A2(n745), .ZN(n750) );
  INV_X1 U845 ( .A(n746), .ZN(n748) );
  AND2_X1 U846 ( .A1(G286), .A2(G8), .ZN(n747) );
  OR2_X1 U847 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U848 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U849 ( .A(n751), .B(KEYINPUT32), .ZN(n760) );
  NAND2_X1 U850 ( .A1(G8), .A2(n752), .ZN(n758) );
  AND2_X1 U851 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U852 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U853 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U854 ( .A1(n760), .A2(n759), .ZN(n776) );
  NOR2_X1 U855 ( .A1(G1971), .A2(G303), .ZN(n761) );
  NOR2_X1 U856 ( .A1(n949), .A2(n761), .ZN(n762) );
  NAND2_X1 U857 ( .A1(n776), .A2(n762), .ZN(n766) );
  NAND2_X1 U858 ( .A1(G1976), .A2(G288), .ZN(n950) );
  NOR2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U860 ( .A1(KEYINPUT33), .A2(n767), .ZN(n768) );
  XOR2_X1 U861 ( .A(KEYINPUT105), .B(n768), .Z(n769) );
  NOR2_X1 U862 ( .A1(n943), .A2(n769), .ZN(n770) );
  NAND2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n784) );
  XOR2_X1 U864 ( .A(n772), .B(KEYINPUT24), .Z(n773) );
  AND2_X1 U865 ( .A1(n773), .A2(n780), .ZN(n782) );
  NOR2_X1 U866 ( .A1(G2090), .A2(G303), .ZN(n774) );
  XOR2_X1 U867 ( .A(KEYINPUT106), .B(n774), .Z(n775) );
  NOR2_X1 U868 ( .A1(n744), .A2(n775), .ZN(n778) );
  INV_X1 U869 ( .A(n776), .ZN(n777) );
  NOR2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n819) );
  XOR2_X1 U874 ( .A(G2067), .B(KEYINPUT37), .Z(n785) );
  XNOR2_X1 U875 ( .A(KEYINPUT97), .B(n785), .ZN(n829) );
  NAND2_X1 U876 ( .A1(n896), .A2(G104), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n895), .A2(G140), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U879 ( .A(KEYINPUT34), .B(n788), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n892), .A2(G128), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n891), .A2(G116), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U883 ( .A(KEYINPUT35), .B(n791), .Z(n792) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U885 ( .A(KEYINPUT36), .B(n794), .ZN(n875) );
  NOR2_X1 U886 ( .A1(n829), .A2(n875), .ZN(n975) );
  NOR2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n831) );
  NAND2_X1 U888 ( .A1(n975), .A2(n831), .ZN(n828) );
  NAND2_X1 U889 ( .A1(G107), .A2(n891), .ZN(n798) );
  NAND2_X1 U890 ( .A1(G131), .A2(n895), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n892), .A2(G119), .ZN(n799) );
  XNOR2_X1 U893 ( .A(n799), .B(KEYINPUT98), .ZN(n801) );
  NAND2_X1 U894 ( .A1(G95), .A2(n896), .ZN(n800) );
  NAND2_X1 U895 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n874) );
  INV_X1 U897 ( .A(G1991), .ZN(n923) );
  NOR2_X1 U898 ( .A1(n874), .A2(n923), .ZN(n813) );
  NAND2_X1 U899 ( .A1(G105), .A2(n896), .ZN(n804) );
  XNOR2_X1 U900 ( .A(n804), .B(KEYINPUT38), .ZN(n811) );
  NAND2_X1 U901 ( .A1(G129), .A2(n892), .ZN(n806) );
  NAND2_X1 U902 ( .A1(G141), .A2(n895), .ZN(n805) );
  NAND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n809) );
  NAND2_X1 U904 ( .A1(G117), .A2(n891), .ZN(n807) );
  XNOR2_X1 U905 ( .A(KEYINPUT99), .B(n807), .ZN(n808) );
  NOR2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(n902) );
  AND2_X1 U908 ( .A1(n902), .A2(G1996), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n979) );
  INV_X1 U910 ( .A(n831), .ZN(n814) );
  NOR2_X1 U911 ( .A1(n979), .A2(n814), .ZN(n822) );
  INV_X1 U912 ( .A(n822), .ZN(n815) );
  NAND2_X1 U913 ( .A1(n828), .A2(n815), .ZN(n817) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n959) );
  AND2_X1 U915 ( .A1(n959), .A2(n831), .ZN(n816) );
  NOR2_X1 U916 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U917 ( .A1(n819), .A2(n818), .ZN(n835) );
  NOR2_X1 U918 ( .A1(G1996), .A2(n902), .ZN(n989) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n820) );
  AND2_X1 U920 ( .A1(n923), .A2(n874), .ZN(n981) );
  NOR2_X1 U921 ( .A1(n820), .A2(n981), .ZN(n821) );
  NOR2_X1 U922 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U923 ( .A(KEYINPUT107), .B(n823), .Z(n824) );
  NOR2_X1 U924 ( .A1(n989), .A2(n824), .ZN(n825) );
  XNOR2_X1 U925 ( .A(n825), .B(KEYINPUT108), .ZN(n826) );
  XNOR2_X1 U926 ( .A(n826), .B(KEYINPUT39), .ZN(n827) );
  NAND2_X1 U927 ( .A1(n828), .A2(n827), .ZN(n830) );
  NAND2_X1 U928 ( .A1(n829), .A2(n875), .ZN(n973) );
  NAND2_X1 U929 ( .A1(n830), .A2(n973), .ZN(n832) );
  NAND2_X1 U930 ( .A1(n832), .A2(n831), .ZN(n833) );
  XOR2_X1 U931 ( .A(KEYINPUT109), .B(n833), .Z(n834) );
  NAND2_X1 U932 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U933 ( .A(KEYINPUT40), .B(n836), .ZN(G329) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U936 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n839) );
  XOR2_X1 U938 ( .A(KEYINPUT111), .B(n839), .Z(n841) );
  NAND2_X1 U939 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G69), .ZN(G235) );
  NOR2_X1 U944 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n844), .B(KEYINPUT112), .ZN(G325) );
  INV_X1 U946 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U947 ( .A(KEYINPUT113), .B(n845), .ZN(G319) );
  XOR2_X1 U948 ( .A(G2100), .B(G2096), .Z(n847) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(G2678), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U951 ( .A(KEYINPUT43), .B(G2090), .Z(n849) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U953 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U954 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U955 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n853), .B(n852), .ZN(G227) );
  XOR2_X1 U957 ( .A(G2474), .B(G1976), .Z(n855) );
  XNOR2_X1 U958 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U959 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U960 ( .A(n856), .B(KEYINPUT114), .Z(n858) );
  XNOR2_X1 U961 ( .A(G1981), .B(G1956), .ZN(n857) );
  XNOR2_X1 U962 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U963 ( .A(G1986), .B(G1971), .Z(n860) );
  XNOR2_X1 U964 ( .A(G1966), .B(G1961), .ZN(n859) );
  XNOR2_X1 U965 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U966 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U967 ( .A(KEYINPUT115), .B(KEYINPUT41), .ZN(n863) );
  XNOR2_X1 U968 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U969 ( .A1(G112), .A2(n891), .ZN(n866) );
  NAND2_X1 U970 ( .A1(G136), .A2(n895), .ZN(n865) );
  NAND2_X1 U971 ( .A1(n866), .A2(n865), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G124), .A2(n892), .ZN(n867) );
  XNOR2_X1 U973 ( .A(n867), .B(KEYINPUT44), .ZN(n868) );
  XNOR2_X1 U974 ( .A(n868), .B(KEYINPUT116), .ZN(n870) );
  NAND2_X1 U975 ( .A1(G100), .A2(n896), .ZN(n869) );
  NAND2_X1 U976 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U977 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U978 ( .A(KEYINPUT117), .B(n873), .Z(G162) );
  XNOR2_X1 U979 ( .A(G162), .B(n977), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U981 ( .A(n877), .B(n876), .ZN(n881) );
  XOR2_X1 U982 ( .A(KEYINPUT46), .B(KEYINPUT118), .Z(n879) );
  XNOR2_X1 U983 ( .A(KEYINPUT119), .B(KEYINPUT48), .ZN(n878) );
  XNOR2_X1 U984 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U985 ( .A(n881), .B(n880), .Z(n890) );
  NAND2_X1 U986 ( .A1(G139), .A2(n895), .ZN(n883) );
  NAND2_X1 U987 ( .A1(G103), .A2(n896), .ZN(n882) );
  NAND2_X1 U988 ( .A1(n883), .A2(n882), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G115), .A2(n891), .ZN(n885) );
  NAND2_X1 U990 ( .A1(G127), .A2(n892), .ZN(n884) );
  NAND2_X1 U991 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n886), .Z(n887) );
  NOR2_X1 U993 ( .A1(n888), .A2(n887), .ZN(n984) );
  XNOR2_X1 U994 ( .A(G160), .B(n984), .ZN(n889) );
  XNOR2_X1 U995 ( .A(n890), .B(n889), .ZN(n906) );
  NAND2_X1 U996 ( .A1(G118), .A2(n891), .ZN(n894) );
  NAND2_X1 U997 ( .A1(G130), .A2(n892), .ZN(n893) );
  NAND2_X1 U998 ( .A1(n894), .A2(n893), .ZN(n901) );
  NAND2_X1 U999 ( .A1(G142), .A2(n895), .ZN(n898) );
  NAND2_X1 U1000 ( .A1(G106), .A2(n896), .ZN(n897) );
  NAND2_X1 U1001 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U1002 ( .A(n899), .B(KEYINPUT45), .Z(n900) );
  NOR2_X1 U1003 ( .A1(n901), .A2(n900), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1005 ( .A(G164), .B(n904), .ZN(n905) );
  XNOR2_X1 U1006 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n907), .ZN(G395) );
  XOR2_X1 U1008 ( .A(n908), .B(G286), .Z(n911) );
  XNOR2_X1 U1009 ( .A(G171), .B(n909), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n912), .ZN(G397) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n914), .ZN(n916) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n915) );
  AND2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n917), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1020 ( .A(G32), .B(n918), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n919), .A2(G28), .ZN(n922) );
  XOR2_X1 U1022 ( .A(KEYINPUT121), .B(G2072), .Z(n920) );
  XNOR2_X1 U1023 ( .A(G33), .B(n920), .ZN(n921) );
  NOR2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n931) );
  XNOR2_X1 U1025 ( .A(n923), .B(G25), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n924), .B(G26), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(G27), .B(n927), .ZN(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n932), .B(KEYINPUT53), .ZN(n935) );
  XOR2_X1 U1032 ( .A(G2084), .B(G34), .Z(n933) );
  XNOR2_X1 U1033 ( .A(KEYINPUT54), .B(n933), .ZN(n934) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(G35), .B(G2090), .ZN(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(KEYINPUT55), .B(n938), .ZN(n940) );
  INV_X1 U1038 ( .A(G29), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n941), .A2(G11), .ZN(n972) );
  XNOR2_X1 U1041 ( .A(KEYINPUT56), .B(G16), .ZN(n969) );
  XOR2_X1 U1042 ( .A(G168), .B(G1966), .Z(n942) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1044 ( .A(KEYINPUT57), .B(n944), .Z(n945) );
  XNOR2_X1 U1045 ( .A(KEYINPUT122), .B(n945), .ZN(n967) );
  XOR2_X1 U1046 ( .A(G171), .B(G1961), .Z(n948) );
  XNOR2_X1 U1047 ( .A(n946), .B(G1341), .ZN(n947) );
  NOR2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n962) );
  XNOR2_X1 U1049 ( .A(KEYINPUT123), .B(n949), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(G1971), .B(G303), .ZN(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(KEYINPUT124), .B(n954), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(n955), .B(G1956), .ZN(n956) );
  NAND2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1057 ( .A(KEYINPUT125), .B(n960), .Z(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(G1348), .B(n963), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1063 ( .A(KEYINPUT126), .B(n970), .Z(n971) );
  NOR2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n1000) );
  INV_X1 U1065 ( .A(n973), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n983) );
  XOR2_X1 U1067 ( .A(G2084), .B(G160), .Z(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n994) );
  XOR2_X1 U1072 ( .A(G2072), .B(n984), .Z(n986) );
  XOR2_X1 U1073 ( .A(G164), .B(G2078), .Z(n985) );
  NOR2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(KEYINPUT50), .B(n987), .ZN(n992) );
  XOR2_X1 U1076 ( .A(G2090), .B(G162), .Z(n988) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1078 ( .A(KEYINPUT51), .B(n990), .Z(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1081 ( .A(KEYINPUT52), .B(n995), .Z(n996) );
  NOR2_X1 U1082 ( .A1(KEYINPUT55), .A2(n996), .ZN(n997) );
  XOR2_X1 U1083 ( .A(KEYINPUT120), .B(n997), .Z(n998) );
  NAND2_X1 U1084 ( .A1(G29), .A2(n998), .ZN(n999) );
  NAND2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1025) );
  XOR2_X1 U1086 ( .A(G1966), .B(G21), .Z(n1008) );
  XNOR2_X1 U1087 ( .A(G1986), .B(G24), .ZN(n1005) );
  XNOR2_X1 U1088 ( .A(G1971), .B(G22), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G1976), .B(G23), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(KEYINPUT127), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(KEYINPUT58), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1021) );
  XOR2_X1 U1095 ( .A(G1961), .B(G5), .Z(n1019) );
  XNOR2_X1 U1096 ( .A(G20), .B(n1009), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G1981), .B(G6), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(KEYINPUT59), .B(G1348), .Z(n1014) );
  XNOR2_X1 U1102 ( .A(G4), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(n1017), .B(KEYINPUT60), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1022), .Z(n1023) );
  NOR2_X1 U1108 ( .A1(G16), .A2(n1023), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1110 ( .A(n1026), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

