//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G227), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G953), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT80), .A3(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT3), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n198), .A2(new_n194), .A3(KEYINPUT80), .A4(G104), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G107), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n196), .A2(new_n197), .A3(new_n199), .A4(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n204), .B(new_n206), .C1(KEYINPUT1), .C2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n205), .A2(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n203), .A2(G143), .ZN(new_n211));
  OAI211_X1 g025(.A(G128), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT82), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n194), .A3(G104), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT82), .B1(new_n194), .B2(G104), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n200), .A2(G107), .ZN(new_n216));
  OAI211_X1 g030(.A(G101), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n202), .A2(new_n208), .A3(new_n212), .A4(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n218), .B(KEYINPUT10), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT0), .A4(G128), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n210), .A2(new_n211), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT0), .B(G128), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n196), .A2(new_n199), .A3(new_n201), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G101), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(KEYINPUT81), .A3(G101), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT81), .B1(new_n225), .B2(G101), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n224), .B(new_n227), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G134), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G137), .ZN(new_n233));
  INV_X1    g047(.A(G137), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT64), .B1(new_n234), .B2(G134), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT11), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AOI211_X1 g051(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n234), .C2(G134), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n234), .A2(G134), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n232), .B2(G137), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n240), .B1(new_n242), .B2(KEYINPUT11), .ZN(new_n243));
  INV_X1    g057(.A(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n235), .A2(new_n236), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n239), .A2(KEYINPUT67), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT67), .B1(new_n239), .B2(new_n246), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n219), .A2(new_n231), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT83), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n219), .A2(new_n231), .A3(KEYINPUT83), .A4(new_n249), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n219), .A2(new_n231), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n237), .A2(G131), .A3(new_n238), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n244), .B1(new_n243), .B2(new_n245), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n239), .A2(KEYINPUT67), .A3(new_n246), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n193), .B1(new_n254), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT12), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT84), .ZN(new_n265));
  AND4_X1   g079(.A1(new_n202), .A2(new_n208), .A3(new_n212), .A4(new_n217), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n202), .A2(new_n217), .B1(new_n212), .B2(new_n208), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n202), .A2(new_n217), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n212), .A2(new_n208), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT84), .A3(new_n218), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n268), .A2(new_n261), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n239), .A2(new_n246), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n266), .B2(new_n267), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT12), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  AOI211_X1 g091(.A(new_n192), .B(new_n277), .C1(new_n252), .C2(new_n253), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n187), .B(new_n188), .C1(new_n263), .C2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n187), .A2(new_n188), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n254), .A2(new_n262), .A3(new_n193), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n277), .B1(new_n252), .B2(new_n253), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n282), .B(G469), .C1(new_n193), .C2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT9), .B(G234), .ZN(new_n286));
  OAI21_X1  g100(.A(G221), .B1(new_n286), .B2(G902), .ZN(new_n287));
  OAI21_X1  g101(.A(G214), .B1(G237), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G210), .B1(G237), .B2(G902), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G125), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n270), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n293), .B1(new_n224), .B2(new_n292), .ZN(new_n294));
  INV_X1    g108(.A(G224), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(G953), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n294), .B(new_n296), .Z(new_n297));
  XOR2_X1   g111(.A(G116), .B(G119), .Z(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT2), .B(G113), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n298), .A2(KEYINPUT66), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT2), .B(G113), .Z(new_n302));
  XNOR2_X1  g116(.A(G116), .B(G119), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI22_X1  g118(.A1(new_n300), .A2(new_n304), .B1(new_n303), .B2(new_n302), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n227), .B(new_n305), .C1(new_n229), .C2(new_n230), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT5), .ZN(new_n307));
  INV_X1    g121(.A(G119), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(G116), .ZN(new_n309));
  OAI211_X1 g123(.A(G113), .B(new_n309), .C1(new_n298), .C2(new_n307), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n300), .B2(new_n304), .ZN(new_n311));
  OR2_X1    g125(.A1(new_n311), .A2(new_n269), .ZN(new_n312));
  XNOR2_X1  g126(.A(G110), .B(G122), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n306), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT6), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n306), .A2(new_n312), .ZN(new_n316));
  INV_X1    g130(.A(new_n313), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT85), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n322));
  AOI211_X1 g136(.A(new_n322), .B(new_n318), .C1(new_n306), .C2(new_n312), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n297), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT7), .B1(new_n295), .B2(G953), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n294), .B(new_n326), .ZN(new_n327));
  XOR2_X1   g141(.A(new_n313), .B(KEYINPUT8), .Z(new_n328));
  NAND2_X1  g142(.A1(new_n311), .A2(new_n269), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n312), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n314), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n188), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n291), .B1(new_n325), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n297), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n314), .A2(KEYINPUT6), .B1(new_n316), .B2(new_n319), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(new_n323), .ZN(new_n337));
  AOI21_X1  g151(.A(G902), .B1(new_n331), .B2(new_n314), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n290), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n289), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n285), .A2(new_n287), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT91), .ZN(new_n342));
  INV_X1    g156(.A(G475), .ZN(new_n343));
  INV_X1    g157(.A(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G125), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n292), .A2(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G146), .ZN(new_n348));
  XNOR2_X1  g162(.A(G125), .B(G140), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n203), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n349), .B2(new_n203), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(G237), .A2(G953), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(G143), .A3(G214), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(G143), .B1(new_n355), .B2(G214), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT18), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n359), .A2(new_n244), .A3(KEYINPUT86), .ZN(new_n360));
  OR3_X1    g174(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n360), .B1(new_n357), .B2(new_n358), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n354), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT17), .B(G131), .C1(new_n357), .C2(new_n358), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT88), .ZN(new_n365));
  OAI21_X1  g179(.A(G131), .B1(new_n357), .B2(new_n358), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n355), .A2(G214), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n205), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n244), .A3(new_n356), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT17), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT16), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n344), .A3(G125), .ZN(new_n373));
  OAI211_X1 g187(.A(G146), .B(new_n373), .C1(new_n347), .C2(new_n372), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n349), .A2(KEYINPUT16), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n373), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n203), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n363), .B1(new_n365), .B2(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(G113), .B(G122), .Z(new_n380));
  XOR2_X1   g194(.A(KEYINPUT87), .B(G104), .Z(new_n381));
  XOR2_X1   g195(.A(new_n380), .B(new_n381), .Z(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n382), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n363), .B(new_n384), .C1(new_n365), .C2(new_n378), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n343), .B1(new_n386), .B2(new_n188), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT20), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n366), .A2(new_n369), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n349), .A2(KEYINPUT19), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n349), .A2(KEYINPUT19), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n203), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n374), .A2(KEYINPUT75), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT75), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n375), .A2(new_n395), .A3(G146), .A4(new_n373), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n390), .A2(new_n393), .A3(new_n394), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n363), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n382), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n385), .ZN(new_n400));
  NOR2_X1   g214(.A1(G475), .A2(G902), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n389), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n400), .A2(new_n389), .A3(new_n401), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n388), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G217), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n286), .A2(new_n405), .A3(G953), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT89), .B1(new_n207), .B2(G143), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT89), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n205), .A3(G128), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n205), .A2(G128), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n232), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G116), .B(G122), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n194), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(G107), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT13), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n409), .B1(G128), .B2(new_n205), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n207), .A2(KEYINPUT89), .A3(G143), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT90), .A3(new_n413), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT90), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT13), .B1(new_n408), .B2(new_n410), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n425), .B1(new_n426), .B2(new_n412), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n411), .A2(new_n420), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n424), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n419), .B1(new_n430), .B2(G134), .ZN(new_n431));
  INV_X1    g245(.A(G122), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G116), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n194), .B1(new_n433), .B2(KEYINPUT14), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n416), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n416), .A2(new_n434), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n411), .A2(new_n413), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G134), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n414), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n407), .B1(new_n431), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n414), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n435), .A3(new_n436), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n412), .B1(new_n411), .B2(new_n420), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n428), .B1(new_n444), .B2(KEYINPUT90), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n232), .B1(new_n445), .B2(new_n427), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n443), .B(new_n406), .C1(new_n446), .C2(new_n419), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n188), .ZN(new_n449));
  INV_X1    g263(.A(G478), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(KEYINPUT15), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(G902), .B1(new_n441), .B2(new_n447), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(KEYINPUT15), .B2(new_n450), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G952), .ZN(new_n456));
  AOI211_X1 g270(.A(G953), .B(new_n456), .C1(G234), .C2(G237), .ZN(new_n457));
  INV_X1    g271(.A(G953), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n188), .B(new_n458), .C1(G234), .C2(G237), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(G898), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n404), .A2(new_n455), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n341), .A2(new_n342), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n285), .A2(new_n462), .A3(new_n340), .A4(new_n287), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT91), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT69), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n355), .A2(G210), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n466), .B(KEYINPUT69), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n469), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT26), .B(G101), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n471), .A2(new_n473), .A3(new_n475), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n224), .B1(new_n247), .B2(new_n248), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n232), .A2(G137), .ZN(new_n481));
  OAI21_X1  g295(.A(G131), .B1(new_n481), .B2(new_n240), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n212), .A2(new_n208), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n246), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(KEYINPUT30), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n224), .B1(new_n257), .B2(new_n258), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n484), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT65), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n223), .B1(new_n239), .B2(new_n246), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n212), .A2(new_n208), .A3(new_n482), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n257), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(KEYINPUT65), .B(new_n488), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n485), .B(new_n305), .C1(new_n489), .C2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n492), .A2(new_n305), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n480), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n479), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT28), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n223), .B1(new_n259), .B2(new_n260), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n298), .A2(new_n299), .ZN(new_n501));
  OAI221_X1 g315(.A(new_n501), .B1(new_n300), .B2(new_n304), .C1(new_n257), .C2(new_n491), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n499), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n480), .A2(new_n496), .B1(new_n487), .B2(new_n305), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n479), .B(new_n503), .C1(new_n504), .C2(new_n499), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT29), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n188), .B1(new_n498), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT28), .B1(new_n480), .B2(new_n496), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n479), .A2(KEYINPUT29), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n305), .B1(new_n500), .B2(new_n492), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT72), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT72), .B(new_n305), .C1(new_n500), .C2(new_n492), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n497), .A3(new_n514), .ZN(new_n515));
  AOI211_X1 g329(.A(new_n509), .B(new_n510), .C1(new_n515), .C2(KEYINPUT28), .ZN(new_n516));
  OAI21_X1  g330(.A(G472), .B1(new_n508), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(G472), .A2(G902), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n518), .B(KEYINPUT71), .Z(new_n519));
  INV_X1    g333(.A(KEYINPUT32), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n477), .A2(new_n478), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n305), .B1(new_n490), .B2(new_n492), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n499), .B1(new_n497), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n522), .B(new_n523), .C1(new_n525), .C2(new_n509), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n479), .A2(new_n497), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n492), .B1(new_n261), .B2(new_n224), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT65), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n274), .A2(new_n224), .B1(new_n483), .B2(new_n246), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n529), .B1(new_n530), .B2(KEYINPUT30), .ZN(new_n531));
  AOI22_X1  g345(.A1(KEYINPUT30), .A2(new_n528), .B1(new_n531), .B2(new_n493), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n527), .B1(new_n532), .B2(new_n305), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT31), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n526), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n500), .A2(new_n502), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(new_n523), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n495), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n524), .B1(new_n500), .B2(new_n502), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT28), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n479), .B1(new_n540), .B2(new_n503), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n538), .B1(new_n541), .B2(new_n522), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n521), .B1(new_n535), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n523), .B1(new_n525), .B2(new_n509), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n533), .A2(new_n534), .B1(new_n544), .B2(KEYINPUT70), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n495), .A2(new_n537), .ZN(new_n546));
  AOI22_X1  g360(.A1(KEYINPUT31), .A2(new_n546), .B1(new_n541), .B2(new_n522), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n519), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n517), .B(new_n543), .C1(new_n548), .C2(KEYINPUT32), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT79), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n405), .B1(G234), .B2(new_n188), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT24), .B(G110), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n308), .A2(G128), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n207), .A2(G119), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT73), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n554), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT74), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n308), .A2(G128), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n555), .B(new_n564), .C1(new_n565), .C2(KEYINPUT23), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G110), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n562), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT74), .B1(new_n561), .B2(new_n567), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n353), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n351), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n394), .A2(new_n396), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n458), .A2(G221), .A3(G234), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT77), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT78), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(KEYINPUT77), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT78), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n576), .A2(KEYINPUT77), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT22), .B(G137), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n578), .A2(new_n582), .A3(new_n584), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n377), .A2(new_n374), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n566), .A2(G110), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n558), .A2(new_n560), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(new_n553), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n575), .A2(new_n589), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n573), .A2(new_n394), .A3(new_n396), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n569), .B2(new_n570), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n588), .B1(new_n598), .B2(new_n594), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n188), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT25), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n552), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n551), .A2(G902), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n549), .A2(new_n550), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n550), .B1(new_n549), .B2(new_n608), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n463), .B(new_n465), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  INV_X1    g426(.A(G472), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n546), .A2(KEYINPUT31), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n509), .B1(KEYINPUT28), .B2(new_n539), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT70), .B1(new_n615), .B2(new_n479), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n614), .A2(new_n616), .A3(new_n526), .A4(new_n538), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n613), .B1(new_n617), .B2(new_n188), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(KEYINPUT92), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT92), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n620), .B(new_n613), .C1(new_n617), .C2(new_n188), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n619), .A2(new_n621), .A3(new_n548), .ZN(new_n622));
  INV_X1    g436(.A(new_n461), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n340), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n441), .A2(new_n447), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n441), .B2(new_n447), .ZN(new_n627));
  OAI211_X1 g441(.A(G478), .B(new_n188), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT94), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT93), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n449), .B2(new_n450), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n453), .A2(KEYINPUT93), .A3(G478), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n628), .B(new_n629), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n449), .A2(new_n630), .A3(new_n450), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT93), .B1(new_n453), .B2(G478), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n629), .B1(new_n637), .B2(new_n628), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n404), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n624), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n285), .A2(new_n287), .ZN(new_n641));
  INV_X1    g455(.A(new_n608), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n622), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n400), .A2(new_n401), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT20), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n400), .A2(new_n389), .A3(new_n401), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(KEYINPUT95), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT95), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n402), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n651), .A2(new_n455), .A3(new_n388), .A4(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n647), .B1(new_n654), .B2(new_n461), .ZN(new_n655));
  AOI211_X1 g469(.A(KEYINPUT95), .B(new_n389), .C1(new_n400), .C2(new_n401), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n403), .A2(new_n402), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n656), .B1(new_n657), .B2(KEYINPUT95), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n387), .B1(new_n452), .B2(new_n454), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n658), .A2(KEYINPUT96), .A3(new_n623), .A4(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n655), .A2(new_n340), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT97), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n655), .A2(new_n660), .A3(KEYINPUT97), .A4(new_n340), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n622), .A3(new_n643), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  INV_X1    g482(.A(KEYINPUT98), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n575), .A2(new_n595), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n589), .A2(KEYINPUT36), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n606), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n669), .B1(new_n605), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(KEYINPUT25), .B1(new_n600), .B2(new_n188), .ZN(new_n676));
  AOI211_X1 g490(.A(new_n602), .B(G902), .C1(new_n596), .C2(new_n599), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n551), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(KEYINPUT98), .A3(new_n673), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n463), .A2(new_n622), .A3(new_n465), .A4(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n459), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n457), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n654), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n341), .A2(new_n549), .A3(new_n680), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XNOR2_X1  g505(.A(new_n687), .B(KEYINPUT39), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n641), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT40), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n536), .B1(new_n511), .B2(new_n512), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n523), .A3(new_n514), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n536), .B1(new_n532), .B2(new_n305), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n188), .B(new_n697), .C1(new_n698), .C2(new_n523), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G472), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n543), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n519), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT32), .B1(new_n617), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT99), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n702), .B1(new_n535), .B2(new_n542), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n520), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n617), .A2(new_n521), .B1(new_n699), .B2(G472), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT99), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n337), .A2(new_n290), .A3(new_n338), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n290), .B1(new_n337), .B2(new_n338), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n713), .A2(KEYINPUT38), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(KEYINPUT38), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n404), .A2(new_n455), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n288), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n716), .A2(new_n680), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n695), .A2(new_n710), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  NOR2_X1   g535(.A1(new_n657), .A2(new_n387), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT94), .ZN(new_n724));
  AOI211_X1 g538(.A(new_n722), .B(new_n688), .C1(new_n724), .C2(new_n633), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n341), .A2(new_n725), .A3(new_n549), .A4(new_n680), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  OAI21_X1  g541(.A(new_n188), .B1(new_n263), .B2(new_n278), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n729), .A2(new_n287), .A3(new_n279), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n549), .A2(new_n730), .A3(new_n608), .ZN(new_n731));
  INV_X1    g545(.A(new_n624), .ZN(new_n732));
  INV_X1    g546(.A(new_n639), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT41), .B(G113), .Z(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  AND3_X1   g551(.A1(new_n549), .A2(new_n730), .A3(new_n608), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n665), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  NAND3_X1  g554(.A1(new_n549), .A2(new_n680), .A3(new_n462), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n340), .A2(new_n287), .A3(new_n729), .A4(new_n279), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n308), .ZN(G21));
  INV_X1    g558(.A(KEYINPUT101), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n509), .B1(new_n515), .B2(KEYINPUT28), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT100), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n523), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n499), .B1(new_n696), .B2(new_n514), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n749), .A2(KEYINPUT100), .A3(new_n509), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n745), .B(new_n614), .C1(new_n748), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n538), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n746), .A2(new_n747), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT100), .B1(new_n749), .B2(new_n509), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n523), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n745), .B1(new_n755), .B2(new_n614), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n702), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n618), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n729), .A2(new_n287), .A3(new_n279), .A4(new_n623), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n717), .A2(new_n340), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n757), .A2(new_n608), .A3(new_n758), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  NAND2_X1  g577(.A1(new_n724), .A2(new_n633), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n404), .A3(new_n687), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n742), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n757), .A2(new_n766), .A3(new_n758), .A4(new_n680), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G125), .ZN(G27));
  NOR3_X1   g582(.A1(new_n711), .A2(new_n712), .A3(new_n289), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n285), .A2(new_n769), .A3(new_n287), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(KEYINPUT42), .A3(new_n725), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT102), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n543), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n617), .A2(KEYINPUT102), .A3(new_n521), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n517), .B1(new_n548), .B2(KEYINPUT32), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n608), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT103), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n706), .A2(new_n773), .A3(new_n517), .A4(new_n774), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(KEYINPUT103), .A3(new_n608), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n771), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n770), .A2(new_n549), .A3(new_n608), .A4(new_n725), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT42), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n782), .A2(new_n785), .A3(KEYINPUT104), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT104), .ZN(new_n787));
  INV_X1    g601(.A(new_n771), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n780), .A2(KEYINPUT103), .A3(new_n608), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT103), .B1(new_n780), .B2(new_n608), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n783), .A2(new_n784), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G131), .ZN(G33));
  AND3_X1   g609(.A1(new_n770), .A2(new_n549), .A3(new_n608), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n689), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  INV_X1    g612(.A(new_n769), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n764), .A2(new_n722), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT43), .B1(new_n722), .B2(KEYINPUT105), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n764), .B(new_n722), .C1(KEYINPUT105), .C2(KEYINPUT43), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT106), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT106), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(new_n806), .A3(new_n803), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n622), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n680), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT44), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n799), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n813));
  INV_X1    g627(.A(new_n282), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n283), .A2(new_n193), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n282), .B(KEYINPUT45), .C1(new_n193), .C2(new_n283), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(G469), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(KEYINPUT46), .A3(new_n281), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT46), .B1(new_n818), .B2(new_n281), .ZN(new_n821));
  INV_X1    g635(.A(new_n279), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n287), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n823), .A2(new_n824), .A3(new_n693), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n812), .B(new_n825), .C1(new_n811), .C2(new_n810), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G137), .ZN(G39));
  OR4_X1    g641(.A1(new_n549), .A2(new_n765), .A3(new_n608), .A4(new_n799), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT47), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n829), .B1(new_n823), .B2(new_n824), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n821), .A2(new_n822), .ZN(new_n831));
  OAI211_X1 g645(.A(KEYINPUT47), .B(new_n287), .C1(new_n831), .C2(new_n820), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n828), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(new_n344), .ZN(G42));
  INV_X1    g648(.A(new_n800), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n716), .A2(new_n835), .A3(new_n287), .A4(new_n288), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n729), .A2(new_n279), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT49), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n836), .A2(new_n838), .A3(new_n710), .A4(new_n642), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT107), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n639), .A2(KEYINPUT108), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n722), .A2(new_n455), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT108), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n764), .A2(new_n843), .A3(new_n404), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n622), .A3(new_n732), .A4(new_n643), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n611), .A2(new_n681), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n738), .A2(new_n640), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n549), .A2(new_n680), .ZN(new_n849));
  INV_X1    g663(.A(new_n742), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n462), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n739), .A2(new_n762), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n791), .A2(new_n792), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT104), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n791), .A2(new_n787), .A3(new_n792), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n285), .A2(new_n769), .A3(new_n287), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n765), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n757), .A2(new_n858), .A3(new_n758), .A4(new_n680), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n455), .A2(new_n387), .A3(new_n688), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n849), .A2(new_n658), .A3(new_n770), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n797), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n853), .A2(new_n855), .A3(new_n856), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  INV_X1    g679(.A(new_n767), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n701), .A2(new_n703), .A3(KEYINPUT99), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n708), .B1(new_n706), .B2(new_n707), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n760), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n285), .A2(new_n287), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n605), .A2(new_n674), .A3(new_n688), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n690), .B(new_n726), .C1(new_n869), .C2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n865), .B1(new_n866), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n690), .A2(new_n726), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n710), .A2(new_n871), .A3(new_n870), .A4(new_n872), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(KEYINPUT52), .A3(new_n767), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT53), .B1(new_n864), .B2(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n786), .A2(new_n793), .A3(new_n862), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n882), .A2(new_n883), .A3(new_n879), .A4(new_n853), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n881), .A2(new_n884), .A3(KEYINPUT54), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n864), .B2(new_n880), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n779), .A2(new_n781), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n888), .A2(new_n788), .B1(new_n784), .B2(new_n783), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT109), .B1(new_n889), .B2(new_n852), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n731), .B1(new_n663), .B2(new_n664), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n891), .A2(new_n735), .A3(new_n743), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT109), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n854), .A2(new_n892), .A3(new_n893), .A4(new_n762), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n611), .A2(KEYINPUT53), .A3(new_n681), .A4(new_n846), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n862), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n890), .A2(new_n894), .A3(new_n879), .A4(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n886), .A2(new_n887), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT111), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n730), .A2(new_n899), .A3(new_n769), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n729), .A2(new_n287), .A3(new_n279), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT111), .B1(new_n799), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n704), .A2(new_n709), .A3(new_n457), .A4(new_n608), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n456), .B(G953), .C1(new_n905), .C2(new_n733), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n686), .B1(new_n802), .B2(new_n803), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(new_n608), .A3(new_n758), .A4(new_n757), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n907), .A2(new_n902), .A3(new_n900), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT48), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n888), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n909), .B2(new_n888), .ZN(new_n912));
  OAI221_X1 g726(.A(new_n906), .B1(new_n742), .B2(new_n908), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n908), .A2(new_n799), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n830), .A2(new_n832), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n837), .A2(new_n287), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT110), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(KEYINPUT50), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n716), .A2(new_n289), .A3(new_n730), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n908), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n757), .A2(new_n758), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n642), .ZN(new_n923));
  INV_X1    g737(.A(new_n919), .ZN(new_n924));
  INV_X1    g738(.A(new_n920), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n907), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n922), .B1(new_n675), .B2(new_n679), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n764), .A2(new_n404), .ZN(new_n929));
  AOI22_X1  g743(.A1(new_n928), .A2(new_n909), .B1(new_n905), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n917), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT51), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT51), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n917), .A2(new_n927), .A3(new_n933), .A4(new_n930), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n913), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n885), .A2(new_n898), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT112), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n885), .A2(new_n898), .A3(new_n935), .A4(KEYINPUT112), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n456), .A2(new_n458), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n840), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT113), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(KEYINPUT113), .B(new_n840), .C1(new_n938), .C2(new_n941), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(G75));
  INV_X1    g760(.A(KEYINPUT56), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n886), .A2(new_n897), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(G902), .ZN(new_n949));
  INV_X1    g763(.A(G210), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n336), .A2(new_n323), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT114), .Z(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT55), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT115), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(new_n297), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n951), .B(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n458), .A2(G952), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT116), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n957), .A2(new_n960), .ZN(G51));
  NAND2_X1  g775(.A1(new_n948), .A2(KEYINPUT54), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n898), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n280), .B(KEYINPUT57), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n263), .A2(new_n278), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT117), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n949), .A2(new_n818), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n958), .B1(new_n968), .B2(new_n969), .ZN(G54));
  INV_X1    g784(.A(KEYINPUT58), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n949), .A2(new_n971), .A3(new_n343), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n972), .A2(new_n400), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n400), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n974), .A3(new_n958), .ZN(G60));
  OR2_X1    g789(.A1(new_n626), .A2(new_n627), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n885), .A2(new_n898), .ZN(new_n977));
  NAND2_X1  g791(.A1(G478), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT59), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n976), .A2(new_n979), .ZN(new_n981));
  AOI211_X1 g795(.A(new_n960), .B(new_n980), .C1(new_n963), .C2(new_n981), .ZN(G63));
  NAND4_X1  g796(.A1(new_n794), .A2(new_n879), .A3(new_n853), .A4(new_n863), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n890), .A2(new_n894), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n879), .A2(new_n896), .ZN(new_n985));
  AOI22_X1  g799(.A1(new_n883), .A2(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(G217), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT60), .ZN(new_n988));
  OAI21_X1  g802(.A(KEYINPUT118), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT118), .ZN(new_n990));
  INV_X1    g804(.A(new_n988), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n948), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n989), .A2(new_n992), .A3(new_n596), .A4(new_n599), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n989), .A2(new_n992), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n960), .B1(new_n994), .B2(new_n672), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT119), .B1(new_n994), .B2(new_n672), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n993), .B(new_n995), .C1(new_n996), .C2(KEYINPUT61), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n990), .B1(new_n948), .B2(new_n991), .ZN(new_n998));
  AOI211_X1 g812(.A(KEYINPUT118), .B(new_n988), .C1(new_n886), .C2(new_n897), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n672), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT119), .ZN(new_n1001));
  AOI21_X1  g815(.A(KEYINPUT61), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1000), .A2(new_n993), .A3(new_n959), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n997), .A2(new_n1004), .ZN(G66));
  OAI21_X1  g819(.A(G953), .B1(new_n460), .B2(new_n295), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT120), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n853), .B2(G953), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n953), .B1(G898), .B2(new_n458), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT121), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1008), .B(new_n1010), .ZN(G69));
  OAI21_X1  g825(.A(G953), .B1(new_n190), .B2(new_n684), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n532), .B(KEYINPUT122), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n391), .A2(new_n392), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1013), .B(new_n1014), .Z(new_n1015));
  NAND2_X1  g829(.A1(new_n684), .A2(G953), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT125), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n760), .B1(new_n779), .B2(new_n781), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n825), .A2(new_n1020), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n794), .A2(new_n797), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n833), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n876), .A2(new_n767), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1022), .A2(new_n826), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1019), .B1(new_n1025), .B2(new_n458), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1024), .A2(new_n720), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1029), .B(KEYINPUT123), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n1028), .A2(KEYINPUT62), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n857), .A2(new_n693), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n845), .B(new_n1032), .C1(new_n609), .C2(new_n610), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n826), .A2(new_n1031), .A3(new_n1023), .A4(new_n1033), .ZN(new_n1034));
  OAI211_X1 g848(.A(new_n458), .B(new_n1015), .C1(new_n1030), .C2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(KEYINPUT124), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1012), .B1(new_n1036), .B2(KEYINPUT126), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT126), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1019), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g853(.A(KEYINPUT124), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1015), .A2(new_n458), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1040), .B1(new_n1043), .B2(new_n1026), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1039), .B1(new_n1044), .B2(new_n1038), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1037), .B1(new_n1045), .B2(new_n1012), .ZN(G72));
  AND2_X1   g860(.A1(new_n698), .A2(new_n523), .ZN(new_n1047));
  NOR3_X1   g861(.A1(new_n1025), .A2(new_n852), .A3(new_n847), .ZN(new_n1048));
  NAND2_X1  g862(.A1(G472), .A2(G902), .ZN(new_n1049));
  XOR2_X1   g863(.A(new_n1049), .B(KEYINPUT63), .Z(new_n1050));
  INV_X1    g864(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1047), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1050), .B1(new_n698), .B2(new_n523), .ZN(new_n1053));
  NOR2_X1   g867(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g868(.A(new_n1054), .B(KEYINPUT127), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n881), .A2(new_n884), .A3(new_n1055), .ZN(new_n1056));
  OAI211_X1 g870(.A(new_n1052), .B(new_n1056), .C1(G952), .C2(new_n458), .ZN(new_n1057));
  AOI21_X1  g871(.A(new_n1051), .B1(new_n1041), .B2(new_n853), .ZN(new_n1058));
  NOR3_X1   g872(.A1(new_n1058), .A2(new_n523), .A3(new_n698), .ZN(new_n1059));
  NOR2_X1   g873(.A1(new_n1057), .A2(new_n1059), .ZN(G57));
endmodule


