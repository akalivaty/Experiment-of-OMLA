//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1234, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0004(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n205));
  INV_X1    g0005(.A(G116), .ZN(new_n206));
  INV_X1    g0006(.A(G270), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G97), .A2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n209), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n208), .B(new_n213), .C1(G58), .C2(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  INV_X1    g0019(.A(new_n217), .ZN(new_n220));
  OR3_X1    g0020(.A1(new_n220), .A2(KEYINPUT64), .A3(G13), .ZN(new_n221));
  OAI21_X1  g0021(.A(KEYINPUT64), .B1(new_n220), .B2(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n227), .A2(new_n216), .A3(new_n228), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n219), .A2(new_n225), .A3(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G226), .B(G232), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n207), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n202), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n206), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(G58), .B(G68), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n247), .A2(G20), .B1(G159), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT73), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n250), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n251), .A2(G33), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT73), .ZN(new_n258));
  AOI21_X1  g0058(.A(G20), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT74), .B1(new_n259), .B2(KEYINPUT7), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n256), .A2(new_n257), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT73), .ZN(new_n263));
  AOI21_X1  g0063(.A(KEYINPUT73), .B1(new_n256), .B2(new_n257), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n216), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT74), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT7), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n260), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT75), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n269), .A2(new_n270), .A3(G68), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n270), .B1(new_n269), .B2(G68), .ZN(new_n272));
  OAI211_X1 g0072(.A(KEYINPUT16), .B(new_n249), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n228), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT16), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT3), .B(G33), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n267), .B1(new_n277), .B2(G20), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n211), .B1(new_n278), .B2(new_n262), .ZN(new_n279));
  INV_X1    g0079(.A(new_n249), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n273), .A2(new_n275), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n215), .A2(G13), .A3(G20), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n275), .B1(new_n215), .B2(G20), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n284), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n277), .A2(G226), .A3(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G87), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n277), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G223), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n289), .B(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G41), .ZN(new_n297));
  INV_X1    g0097(.A(G45), .ZN(new_n298));
  AOI21_X1  g0098(.A(G1), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G274), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n295), .A2(new_n299), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G232), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n296), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G190), .B2(new_n303), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n282), .A2(new_n288), .A3(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n307), .A2(KEYINPUT17), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(KEYINPUT17), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n282), .A2(new_n288), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n303), .A2(G169), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT76), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n296), .A2(G179), .A3(new_n300), .A4(new_n302), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n312), .B1(new_n311), .B2(new_n313), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT18), .B1(new_n310), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT18), .ZN(new_n320));
  AOI211_X1 g0120(.A(new_n320), .B(new_n317), .C1(new_n282), .C2(new_n288), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n308), .A2(new_n309), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n277), .A2(G223), .A3(G1698), .ZN(new_n323));
  INV_X1    g0123(.A(G222), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n323), .B1(new_n202), .B2(new_n277), .C1(new_n292), .C2(new_n324), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(KEYINPUT67), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(KEYINPUT67), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n295), .A3(new_n327), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n301), .A2(G226), .B1(G274), .B2(new_n299), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT9), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n248), .A2(G150), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n216), .A2(G33), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n332), .B1(new_n201), .B2(new_n216), .C1(new_n283), .C2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G50), .ZN(new_n335));
  INV_X1    g0135(.A(new_n285), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n334), .A2(new_n275), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n287), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n330), .A2(G200), .B1(new_n331), .B2(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n339), .A2(new_n331), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n328), .A2(G190), .A3(new_n329), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT10), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT10), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n340), .A2(new_n345), .A3(new_n341), .A4(new_n342), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n330), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(new_n339), .C1(G179), .C2(new_n330), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n261), .B1(G232), .B2(new_n291), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n212), .B2(new_n291), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n353), .B(new_n295), .C1(G107), .C2(new_n277), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n301), .A2(G244), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n300), .A3(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(G179), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G20), .A2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT68), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n283), .B(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n248), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n358), .B1(new_n359), .B2(new_n333), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n275), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n285), .B(KEYINPUT69), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n202), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT69), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n287), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n364), .B(new_n366), .C1(new_n202), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n356), .A2(new_n348), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n357), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n322), .A2(new_n351), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT13), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n256), .A2(new_n257), .A3(G232), .A4(G1698), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT71), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n256), .A2(new_n257), .A3(G226), .A4(new_n291), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT70), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT71), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n277), .A2(new_n379), .A3(G232), .A4(G1698), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G97), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n376), .A2(new_n378), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n377), .A2(KEYINPUT70), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n295), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n301), .A2(G238), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n300), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n374), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(new_n374), .A3(new_n387), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(G190), .A3(new_n390), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n362), .A2(new_n335), .B1(new_n333), .B2(new_n202), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n216), .A2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n275), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  XOR2_X1   g0194(.A(new_n394), .B(KEYINPUT11), .Z(new_n395));
  NAND2_X1  g0195(.A1(new_n368), .A2(KEYINPUT12), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G68), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n336), .A2(KEYINPUT12), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n365), .A2(KEYINPUT12), .A3(new_n211), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT72), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT72), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n397), .A2(new_n402), .A3(new_n398), .A4(new_n399), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n395), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(KEYINPUT70), .A2(new_n377), .B1(new_n375), .B2(KEYINPUT71), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n377), .A2(KEYINPUT70), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n381), .A4(new_n380), .ZN(new_n407));
  AOI211_X1 g0207(.A(KEYINPUT13), .B(new_n386), .C1(new_n407), .C2(new_n295), .ZN(new_n408));
  OAI21_X1  g0208(.A(G200), .B1(new_n408), .B2(new_n388), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n391), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(G169), .B1(new_n408), .B2(new_n388), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT14), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n389), .A2(G179), .A3(new_n390), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(G169), .C1(new_n408), .C2(new_n388), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n404), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n410), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n356), .A2(G200), .ZN(new_n419));
  INV_X1    g0219(.A(G190), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n356), .A2(new_n420), .ZN(new_n421));
  OR3_X1    g0221(.A1(new_n419), .A2(new_n369), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n373), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n278), .A2(new_n262), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G107), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n248), .A2(KEYINPUT77), .A3(G77), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT77), .B1(new_n248), .B2(G77), .ZN(new_n428));
  INV_X1    g0228(.A(G107), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(KEYINPUT6), .A3(G97), .ZN(new_n430));
  AND2_X1   g0230(.A1(G97), .A2(G107), .ZN(new_n431));
  NOR2_X1   g0231(.A1(G97), .A2(G107), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n430), .B1(new_n433), .B2(KEYINPUT6), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n428), .B1(new_n434), .B2(G20), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n426), .A2(new_n427), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n275), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n285), .A2(G97), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n275), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n215), .A2(G33), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n441), .A3(new_n285), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G97), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n437), .A2(new_n439), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT78), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n438), .B1(new_n436), .B2(new_n275), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(KEYINPUT78), .A3(new_n444), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT5), .B(G41), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n298), .A2(G1), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(G274), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n256), .A2(new_n257), .A3(G244), .A4(new_n291), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(KEYINPUT79), .A2(KEYINPUT4), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n277), .A2(G244), .A3(new_n291), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n277), .A2(G250), .A3(G1698), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n456), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n453), .B1(new_n461), .B2(new_n295), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n450), .A2(new_n451), .ZN(new_n463));
  INV_X1    g0263(.A(new_n295), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(G257), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT80), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n295), .B1(new_n451), .B2(new_n450), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT80), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(G257), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n462), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n447), .A2(new_n449), .B1(G190), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(G200), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT81), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n462), .A2(G179), .A3(new_n470), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n348), .B1(new_n462), .B2(new_n470), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n437), .A2(new_n439), .A3(new_n444), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n445), .B(KEYINPUT81), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n473), .A2(new_n474), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT19), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n216), .B1(new_n381), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G87), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n432), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n216), .A2(G33), .A3(G97), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n485), .A2(new_n487), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n277), .A2(new_n216), .A3(G68), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n275), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n365), .A2(new_n359), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(G87), .B2(new_n443), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n277), .A2(G244), .A3(G1698), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G116), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n496), .B(new_n497), .C1(new_n292), .C2(new_n212), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n295), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n464), .B(G250), .C1(G1), .C2(new_n298), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n451), .A2(G274), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G200), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n495), .B(new_n503), .C1(new_n420), .C2(new_n502), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n492), .B(new_n493), .C1(new_n359), .C2(new_n442), .ZN(new_n505));
  INV_X1    g0305(.A(G179), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n499), .A2(new_n506), .A3(new_n500), .A4(new_n501), .ZN(new_n507));
  INV_X1    g0307(.A(new_n502), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n505), .B(new_n507), .C1(new_n508), .C2(G169), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n277), .A2(G257), .A3(G1698), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n277), .A2(G250), .A3(new_n291), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n295), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n467), .A2(G264), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n515), .A2(new_n452), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(new_n304), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n497), .A2(G20), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n256), .A2(new_n257), .A3(new_n216), .A4(G87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT22), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT22), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n277), .A2(new_n522), .A3(new_n216), .A4(G87), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n519), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n216), .A2(G107), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n525), .B(KEYINPUT23), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT24), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT24), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n524), .A2(new_n529), .A3(new_n526), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n440), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT25), .B1(new_n336), .B2(new_n429), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n336), .A2(KEYINPUT25), .A3(new_n429), .ZN(new_n534));
  AOI22_X1  g0334(.A1(G107), .A2(new_n443), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n515), .A2(new_n452), .A3(new_n516), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(new_n420), .ZN(new_n538));
  NOR4_X1   g0338(.A1(new_n518), .A2(new_n531), .A3(new_n536), .A4(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT84), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n528), .A2(new_n530), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n536), .B1(new_n541), .B2(new_n275), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(new_n348), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(G179), .B2(new_n537), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n540), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n537), .A2(G179), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n514), .A2(new_n295), .B1(G264), .B2(new_n467), .ZN(new_n547));
  AOI21_X1  g0347(.A(G169), .B1(new_n547), .B2(new_n452), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n549), .B(KEYINPUT84), .C1(new_n531), .C2(new_n536), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n539), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n285), .B(new_n367), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(G116), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n552), .A2(G116), .A3(new_n441), .A4(new_n440), .ZN(new_n555));
  INV_X1    g0355(.A(G97), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n460), .B(new_n216), .C1(G33), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT83), .ZN(new_n558));
  AOI21_X1  g0358(.A(G20), .B1(new_n253), .B2(G97), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT83), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(new_n460), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n206), .A2(G20), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n275), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT82), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n275), .A2(KEYINPUT82), .A3(new_n563), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n562), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT20), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n275), .A2(KEYINPUT82), .A3(new_n563), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT82), .B1(new_n275), .B2(new_n563), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT20), .B1(new_n573), .B2(new_n562), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n554), .B(new_n555), .C1(new_n570), .C2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n277), .A2(G257), .A3(new_n291), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n277), .A2(G264), .A3(G1698), .ZN(new_n578));
  INV_X1    g0378(.A(G303), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n277), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(new_n295), .B1(G270), .B2(new_n467), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n452), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G200), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n576), .B(new_n583), .C1(new_n420), .C2(new_n582), .ZN(new_n584));
  INV_X1    g0384(.A(new_n582), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n585), .A2(new_n575), .A3(G179), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT21), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n348), .B1(new_n581), .B2(new_n452), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(new_n575), .B2(new_n588), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n575), .A2(new_n588), .A3(new_n587), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n584), .B(new_n586), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n483), .A2(new_n510), .A3(new_n551), .A4(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n424), .A2(new_n593), .ZN(G372));
  INV_X1    g0394(.A(new_n424), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n586), .B1(new_n590), .B2(new_n589), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT85), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n542), .A2(new_n544), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT85), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n600), .B(new_n586), .C1(new_n590), .C2(new_n589), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n597), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT86), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n472), .A2(G190), .ZN(new_n604));
  AND4_X1   g0404(.A1(KEYINPUT78), .A2(new_n437), .A3(new_n439), .A4(new_n444), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT78), .B1(new_n448), .B2(new_n444), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n474), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n482), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n476), .B1(new_n472), .B2(new_n348), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT81), .B1(new_n609), .B2(new_n445), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n607), .B(new_n510), .C1(new_n608), .C2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n611), .A2(new_n539), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT86), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n597), .A2(new_n613), .A3(new_n599), .A4(new_n601), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n603), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n509), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n510), .A2(new_n481), .A3(new_n482), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n616), .B1(new_n617), .B2(KEYINPUT26), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n605), .A2(new_n606), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT26), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n510), .A2(new_n619), .A3(new_n620), .A4(new_n609), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n595), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n307), .B(KEYINPUT17), .ZN(new_n625));
  INV_X1    g0425(.A(new_n410), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n416), .A2(new_n417), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n371), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n311), .A2(new_n313), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n310), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n320), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n310), .A2(KEYINPUT18), .A3(new_n630), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n347), .B1(new_n629), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(new_n350), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n624), .A2(new_n637), .ZN(G369));
  NAND2_X1  g0438(.A1(new_n597), .A2(new_n601), .ZN(new_n639));
  INV_X1    g0439(.A(G13), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G20), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n215), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n575), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n639), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n591), .B(KEYINPUT87), .Z(new_n650));
  AOI21_X1  g0450(.A(new_n649), .B1(new_n650), .B2(new_n648), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G330), .ZN(new_n652));
  INV_X1    g0452(.A(new_n551), .ZN(new_n653));
  INV_X1    g0453(.A(new_n542), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(new_n647), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n598), .B2(new_n647), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n647), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n596), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n598), .B2(new_n658), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n657), .A2(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n223), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G41), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n487), .A2(G116), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n664), .A2(new_n215), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n226), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n664), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT28), .Z(new_n670));
  NAND2_X1  g0470(.A1(new_n623), .A2(new_n658), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT29), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n617), .A2(KEYINPUT26), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n616), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n510), .A2(new_n619), .A3(new_n609), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n676));
  INV_X1    g0476(.A(new_n611), .ZN(new_n677));
  OR4_X1    g0477(.A1(new_n531), .A2(new_n518), .A3(new_n536), .A4(new_n538), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n545), .A2(new_n550), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n596), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n674), .B(new_n676), .C1(new_n679), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n658), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n672), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n472), .A2(new_n585), .A3(new_n517), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n506), .A3(new_n502), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n462), .A2(new_n581), .A3(G179), .A4(new_n470), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n502), .A2(new_n537), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n689), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR4_X1   g0493(.A1(new_n690), .A2(KEYINPUT30), .A3(new_n502), .A4(new_n537), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n688), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT31), .B1(new_n593), .B2(new_n647), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT88), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n688), .B(KEYINPUT88), .C1(new_n693), .C2(new_n694), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n647), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n697), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G330), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT89), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n589), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n575), .A2(new_n588), .A3(new_n587), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n585), .A2(new_n575), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n706), .A2(new_n707), .B1(new_n708), .B2(G179), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n680), .A2(new_n709), .A3(new_n678), .A4(new_n584), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n710), .A2(new_n611), .A3(new_n647), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n702), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n696), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT89), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(G330), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n705), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n686), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n670), .B1(new_n718), .B2(G1), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT90), .Z(G364));
  AOI21_X1  g0520(.A(new_n215), .B1(new_n641), .B2(G45), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n664), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n223), .A2(G355), .A3(new_n277), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n263), .A2(new_n264), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n663), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(G45), .B2(new_n227), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n242), .A2(new_n298), .ZN(new_n729));
  OAI221_X1 g0529(.A(new_n725), .B1(G116), .B2(new_n223), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G13), .A2(G33), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n228), .B1(G20), .B2(new_n348), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n724), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n733), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n216), .A2(new_n506), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n420), .A3(G200), .ZN(new_n739));
  XOR2_X1   g0539(.A(KEYINPUT33), .B(G317), .Z(new_n740));
  OAI21_X1  g0540(.A(new_n261), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n216), .A2(new_n420), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n506), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n216), .A2(G190), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n304), .A2(G179), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(G322), .A2(new_n745), .B1(new_n749), .B2(G283), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n742), .A2(new_n747), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n750), .B1(new_n579), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G179), .A2(G200), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n746), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n741), .B(new_n752), .C1(G329), .C2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n738), .A2(G190), .A3(G200), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT95), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G326), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n216), .B1(new_n754), .B2(G190), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n764), .A2(KEYINPUT94), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(KEYINPUT94), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n746), .A2(new_n743), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n762), .B1(new_n763), .B2(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n755), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT32), .Z(new_n773));
  INV_X1    g0573(.A(G58), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n744), .A2(new_n774), .B1(new_n769), .B2(new_n202), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT92), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n751), .A2(new_n486), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n739), .A2(new_n211), .B1(new_n758), .B2(new_n335), .ZN(new_n778));
  NOR4_X1   g0578(.A1(new_n773), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n779), .B1(new_n556), .B2(new_n767), .C1(new_n429), .C2(new_n748), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n770), .B1(new_n780), .B2(new_n261), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT96), .Z(new_n782));
  INV_X1    g0582(.A(new_n734), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n736), .B1(new_n651), .B2(new_n737), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT97), .Z(new_n785));
  OR2_X1    g0585(.A1(new_n651), .A2(G330), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n786), .A2(new_n652), .A3(new_n724), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT91), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n785), .A2(new_n788), .ZN(G396));
  AOI21_X1  g0589(.A(new_n647), .B1(new_n615), .B2(new_n622), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT101), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n371), .B(new_n791), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n792), .A2(new_n422), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n369), .A2(new_n647), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n793), .A2(new_n795), .B1(new_n372), .B2(new_n647), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n794), .B1(new_n671), .B2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(new_n717), .Z(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n724), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n751), .A2(new_n335), .B1(new_n748), .B2(new_n211), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT99), .ZN(new_n801));
  INV_X1    g0601(.A(new_n726), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n774), .B2(new_n767), .ZN(new_n804));
  INV_X1    g0604(.A(new_n758), .ZN(new_n805));
  INV_X1    g0605(.A(new_n769), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n805), .A2(G137), .B1(new_n806), .B2(G159), .ZN(new_n807));
  INV_X1    g0607(.A(G150), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n739), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G143), .B2(new_n745), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT98), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n804), .B1(new_n811), .B2(KEYINPUT34), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(KEYINPUT34), .B2(new_n811), .C1(new_n813), .C2(new_n755), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n486), .A2(new_n748), .B1(new_n769), .B2(new_n206), .ZN(new_n815));
  INV_X1    g0615(.A(new_n739), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n277), .B1(new_n816), .B2(G283), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n817), .B1(new_n429), .B2(new_n751), .C1(new_n579), .C2(new_n758), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n815), .B(new_n818), .C1(G311), .C2(new_n756), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n819), .B1(new_n556), .B2(new_n767), .C1(new_n763), .C2(new_n744), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n783), .B1(new_n814), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n734), .A2(new_n731), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n724), .B(new_n821), .C1(new_n202), .C2(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT100), .Z(new_n824));
  INV_X1    g0624(.A(new_n796), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n732), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n799), .A2(new_n826), .ZN(G384));
  INV_X1    g0627(.A(KEYINPUT104), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n627), .A2(new_n658), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n417), .A2(new_n647), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n627), .A2(new_n626), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(KEYINPUT102), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT102), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n418), .B2(new_n831), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n830), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT103), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n832), .A2(KEYINPUT102), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n418), .A2(new_n834), .A3(new_n831), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(KEYINPUT103), .A3(new_n830), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n796), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n677), .A2(new_n551), .A3(new_n592), .A4(new_n658), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n700), .A2(new_n701), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n844), .A2(KEYINPUT31), .B1(new_n845), .B2(new_n647), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n702), .A2(new_n712), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n828), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  INV_X1    g0651(.A(new_n645), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n310), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n634), .B2(new_n625), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n853), .A2(new_n855), .A3(new_n307), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n310), .A2(new_n318), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n631), .A2(new_n853), .A3(new_n307), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n856), .A2(new_n857), .B1(new_n858), .B2(KEYINPUT37), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n851), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n288), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n269), .A2(G68), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT75), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n269), .A2(new_n270), .A3(G68), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n280), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n440), .B1(new_n865), .B2(KEYINPUT16), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n249), .B1(new_n271), .B2(new_n272), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n276), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n861), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n307), .B1(new_n869), .B2(new_n645), .ZN(new_n870));
  INV_X1    g0670(.A(new_n630), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n857), .A2(new_n853), .A3(new_n855), .A4(new_n307), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n869), .A2(new_n645), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n322), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(new_n877), .A3(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n860), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT40), .B1(new_n850), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT103), .B1(new_n841), .B2(new_n830), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n837), .B(new_n829), .C1(new_n839), .C2(new_n840), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n884), .A2(new_n796), .A3(new_n848), .ZN(new_n885));
  NAND2_X1  g0685(.A1(KEYINPUT104), .A2(KEYINPUT40), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n875), .A2(new_n877), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n851), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n878), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n885), .B(new_n886), .C1(KEYINPUT40), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n595), .A2(new_n849), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n891), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(G330), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n627), .A2(new_n647), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n875), .A2(new_n877), .A3(KEYINPUT38), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n875), .B2(new_n877), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT39), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n860), .A2(new_n900), .A3(new_n878), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n896), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n635), .A2(new_n645), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n897), .A2(new_n898), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n838), .A2(new_n842), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n792), .A2(new_n647), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n905), .B1(new_n794), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n903), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n686), .A2(new_n595), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n637), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n909), .B(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n894), .B(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n215), .B2(new_n641), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n206), .B1(new_n434), .B2(KEYINPUT35), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n228), .A2(new_n216), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n915), .B(new_n916), .C1(KEYINPUT35), .C2(new_n434), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT36), .ZN(new_n918));
  OAI21_X1  g0718(.A(G77), .B1(new_n774), .B2(new_n211), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n919), .A2(new_n226), .B1(G50), .B2(new_n211), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(G1), .A3(new_n640), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n914), .A2(new_n918), .A3(new_n921), .ZN(G367));
  INV_X1    g0722(.A(new_n727), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n923), .A2(new_n238), .B1(new_n223), .B2(new_n359), .ZN(new_n924));
  INV_X1    g0724(.A(new_n735), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n723), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT108), .ZN(new_n927));
  INV_X1    g0727(.A(new_n767), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(G107), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n802), .B1(new_n763), .B2(new_n739), .ZN(new_n930));
  INV_X1    g0730(.A(G317), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n755), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n748), .A2(new_n556), .ZN(new_n933));
  INV_X1    g0733(.A(G283), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n744), .A2(new_n579), .B1(new_n769), .B2(new_n934), .ZN(new_n935));
  NOR4_X1   g0735(.A1(new_n930), .A2(new_n932), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n760), .A2(G311), .ZN(new_n937));
  INV_X1    g0737(.A(new_n751), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(G116), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT46), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n929), .A2(new_n936), .A3(new_n937), .A4(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n277), .B1(new_n739), .B2(new_n771), .ZN(new_n942));
  AOI22_X1  g0742(.A1(G150), .A2(new_n745), .B1(new_n806), .B2(G50), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n202), .B2(new_n748), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n942), .B(new_n944), .C1(G137), .C2(new_n756), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n928), .A2(G68), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n760), .A2(G143), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n751), .A2(new_n774), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n941), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT47), .Z(new_n951));
  OAI21_X1  g0751(.A(new_n927), .B1(new_n951), .B2(new_n783), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT109), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n495), .A2(new_n658), .ZN(new_n954));
  MUX2_X1   g0754(.A(new_n510), .B(new_n616), .S(new_n954), .Z(new_n955));
  OAI21_X1  g0755(.A(new_n953), .B1(new_n737), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n657), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n605), .A2(new_n606), .A3(new_n658), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n609), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT105), .ZN(new_n961));
  INV_X1    g0761(.A(new_n959), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n483), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n660), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT42), .Z(new_n967));
  AOI22_X1  g0767(.A1(new_n964), .A2(new_n681), .B1(new_n481), .B2(new_n482), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n647), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n965), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n965), .A3(new_n970), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n974), .B(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n660), .B1(new_n656), .B2(new_n659), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(new_n652), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n718), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  OR3_X1    g0781(.A1(new_n661), .A2(new_n964), .A3(KEYINPUT106), .ZN(new_n982));
  OAI21_X1  g0782(.A(KEYINPUT106), .B1(new_n661), .B2(new_n964), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT44), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n661), .A2(new_n964), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT45), .Z(new_n988));
  NAND3_X1  g0788(.A1(new_n982), .A2(KEYINPUT44), .A3(new_n983), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n958), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n986), .A2(new_n988), .A3(new_n657), .A4(new_n989), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n981), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n718), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n664), .B(KEYINPUT41), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n722), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT107), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n977), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n997), .B1(new_n977), .B2(new_n996), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n957), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT110), .ZN(G387));
  NAND2_X1  g0802(.A1(new_n979), .A2(new_n722), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n361), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n335), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT50), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(KEYINPUT50), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n666), .B1(G68), .B2(G77), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1006), .A2(new_n298), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n235), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n923), .B1(G45), .B2(new_n1010), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n663), .A2(new_n261), .A3(new_n665), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n663), .A2(new_n429), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n925), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n816), .A2(G311), .B1(new_n806), .B2(G303), .ZN(new_n1016));
  INV_X1    g0816(.A(G322), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n931), .B2(new_n744), .C1(new_n759), .C2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT48), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n934), .B2(new_n767), .C1(new_n763), .C2(new_n751), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT49), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n726), .B1(new_n756), .B2(G326), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(new_n206), .C2(new_n748), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n744), .A2(new_n335), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n767), .A2(new_n359), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n938), .A2(G77), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n211), .B2(new_n769), .C1(new_n556), .C2(new_n748), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G150), .B2(new_n756), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n726), .B1(new_n771), .B2(new_n758), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n284), .B2(new_n816), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1025), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1023), .B1(new_n1024), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1015), .B1(new_n1032), .B2(new_n734), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n656), .A2(new_n733), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n723), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n664), .B1(new_n718), .B2(new_n979), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1003), .B(new_n1035), .C1(new_n981), .C2(new_n1036), .ZN(G393));
  NAND3_X1  g0837(.A1(new_n991), .A2(new_n722), .A3(new_n992), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n735), .B1(new_n556), .B2(new_n223), .C1(new_n923), .C2(new_n245), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n277), .B1(new_n749), .B2(G107), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n934), .B2(new_n751), .C1(new_n579), .C2(new_n739), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n758), .A2(new_n931), .B1(new_n744), .B2(new_n768), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT52), .Z(new_n1043));
  AOI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(G322), .C2(new_n756), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n206), .B2(new_n767), .C1(new_n763), .C2(new_n769), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n928), .A2(G77), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n739), .A2(new_n335), .B1(new_n748), .B2(new_n486), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n726), .B1(new_n211), .B2(new_n751), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n1004), .C2(new_n806), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n756), .A2(G143), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n758), .A2(new_n808), .B1(new_n744), .B2(new_n771), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT51), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1045), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n724), .B1(new_n1054), .B2(new_n734), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1039), .B(new_n1055), .C1(new_n964), .C2(new_n737), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n1038), .A2(KEYINPUT111), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT111), .B1(new_n1038), .B2(new_n1056), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n664), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n991), .A2(new_n992), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1060), .B1(new_n1061), .B2(new_n980), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1062), .A2(new_n993), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(G390));
  INV_X1    g0865(.A(KEYINPUT112), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n906), .B1(new_n790), .B2(new_n793), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n896), .B1(new_n884), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n899), .A2(new_n1068), .A3(new_n901), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n683), .A2(new_n658), .A3(new_n793), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1070), .A2(new_n906), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n879), .B(new_n896), .C1(new_n1071), .C2(new_n884), .ZN(new_n1072));
  AOI221_X4 g0872(.A(new_n796), .B1(new_n838), .B2(new_n842), .C1(new_n705), .C2(new_n716), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1069), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n825), .B(G330), .C1(new_n846), .C2(new_n847), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n884), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n595), .A2(G330), .A3(new_n849), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n910), .A2(new_n637), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n905), .B1(new_n717), .B2(new_n825), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1081), .A2(new_n1076), .B1(new_n794), .B2(new_n906), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n715), .B1(new_n714), .B2(G330), .ZN(new_n1083));
  AOI211_X1 g0883(.A(KEYINPUT89), .B(new_n704), .C1(new_n713), .C2(new_n696), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n825), .B(new_n905), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n884), .A2(new_n1075), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n1071), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1080), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1066), .B1(new_n1078), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1078), .A2(new_n1088), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n825), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1076), .B1(new_n1092), .B2(new_n884), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1087), .B1(new_n1093), .B2(new_n1067), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1080), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1091), .A2(KEYINPUT112), .A3(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1089), .A2(new_n664), .A3(new_n1090), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n899), .A2(new_n731), .A3(new_n901), .ZN(new_n1099));
  INV_X1    g0899(.A(G137), .ZN(new_n1100));
  INV_X1    g0900(.A(G128), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n739), .A2(new_n1100), .B1(new_n758), .B2(new_n1101), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n277), .B1(new_n748), .B2(new_n335), .C1(new_n813), .C2(new_n744), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(G125), .C2(new_n756), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n751), .A2(new_n808), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n1106));
  XNOR2_X1  g0906(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT54), .B(G143), .Z(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1108), .B1(new_n771), .B2(new_n767), .C1(new_n769), .C2(new_n1110), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n211), .A2(new_n748), .B1(new_n769), .B2(new_n556), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n777), .B1(G283), .B2(new_n805), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n261), .C1(new_n429), .C2(new_n739), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1112), .B(new_n1114), .C1(G294), .C2(new_n756), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1115), .B(new_n1046), .C1(new_n206), .C2(new_n744), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n783), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n283), .B2(new_n822), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1099), .A2(new_n723), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n1091), .B2(new_n721), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT114), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT114), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1122), .B(new_n1119), .C1(new_n1091), .C2(new_n721), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1098), .A2(new_n1124), .ZN(G378));
  OAI21_X1  g0925(.A(new_n1095), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n339), .A2(new_n852), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n347), .A2(new_n350), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1127), .B1(new_n347), .B2(new_n350), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT55), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1130), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT55), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n1128), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT56), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT119), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1131), .A2(new_n1134), .A3(KEYINPUT56), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(G330), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n881), .B2(new_n890), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n899), .A2(new_n901), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n895), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n884), .A2(new_n1067), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n889), .A2(new_n1145), .B1(new_n635), .B2(new_n645), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1137), .A2(KEYINPUT118), .A3(new_n1139), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(KEYINPUT119), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1147), .A2(KEYINPUT119), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n902), .B2(new_n908), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1142), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1141), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n891), .A2(new_n1153), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1150), .A2(new_n902), .A3(new_n908), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1148), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1126), .A2(KEYINPUT57), .A3(new_n1152), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT120), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT57), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1080), .B1(new_n1078), .B2(new_n1088), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1157), .A2(new_n1152), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1142), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1149), .A2(new_n1151), .B1(new_n891), .B2(new_n1153), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1167), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n1126), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1160), .A2(new_n664), .A3(new_n1164), .A4(new_n1168), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1110), .A2(new_n751), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n739), .A2(new_n813), .B1(new_n769), .B2(new_n1100), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT116), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(G125), .C2(new_n805), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n1101), .B2(new_n744), .C1(new_n808), .C2(new_n767), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT59), .Z(new_n1176));
  AOI21_X1  g0976(.A(G41), .B1(new_n756), .B2(G124), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G33), .B1(new_n749), .B2(G159), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1026), .B1(new_n556), .B2(new_n739), .C1(new_n206), .C2(new_n758), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n748), .A2(new_n774), .ZN(new_n1181));
  NOR4_X1   g0981(.A1(new_n1180), .A2(G41), .A3(new_n726), .A4(new_n1181), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n744), .A2(new_n429), .B1(new_n769), .B2(new_n359), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n756), .B2(G283), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n946), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT115), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n297), .B1(new_n802), .B2(new_n253), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n335), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1187), .B(new_n1188), .C1(new_n1189), .C2(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1179), .B(new_n1192), .C1(new_n1189), .C2(new_n1191), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1170), .A2(new_n731), .B1(new_n734), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n724), .B1(new_n335), .B2(new_n822), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT117), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1167), .A2(new_n722), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1169), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT121), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1169), .A2(KEYINPUT121), .A3(new_n1197), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(G375));
  NAND3_X1  g1002(.A1(new_n1082), .A2(new_n1080), .A3(new_n1087), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1096), .A2(new_n1203), .A3(new_n995), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT122), .Z(new_n1205));
  NAND2_X1  g1005(.A1(new_n884), .A2(new_n731), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n802), .A2(new_n1181), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT124), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n755), .A2(new_n1101), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n1110), .A2(new_n739), .B1(new_n813), .B2(new_n758), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n744), .A2(new_n1100), .B1(new_n769), .B2(new_n808), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n335), .B2(new_n767), .C1(new_n771), .C2(new_n751), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n744), .A2(new_n934), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n739), .A2(new_n206), .B1(new_n758), .B2(new_n763), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G107), .B2(new_n806), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT123), .Z(new_n1217));
  OAI221_X1 g1017(.A(new_n261), .B1(new_n748), .B2(new_n202), .C1(new_n556), .C2(new_n751), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G303), .B2(new_n756), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1025), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1213), .B1(new_n1214), .B2(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1221), .A2(new_n734), .B1(new_n211), .B2(new_n822), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1206), .A2(new_n723), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n1094), .B2(new_n722), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1205), .A2(new_n1224), .ZN(G381));
  INV_X1    g1025(.A(G384), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1064), .A2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(G387), .A2(new_n1227), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1169), .A2(KEYINPUT121), .A3(new_n1197), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT121), .B1(new_n1169), .B2(new_n1197), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1230), .A2(new_n1231), .A3(G378), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1228), .A2(new_n1229), .A3(new_n1232), .ZN(G407));
  INV_X1    g1033(.A(G378), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1200), .A2(new_n1234), .A3(new_n1201), .ZN(new_n1235));
  OAI211_X1 g1035(.A(G407), .B(G213), .C1(G343), .C2(new_n1235), .ZN(G409));
  XOR2_X1   g1036(.A(G393), .B(G396), .Z(new_n1237));
  OR2_X1    g1037(.A1(new_n1064), .A2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1064), .B1(new_n1237), .B2(KEYINPUT110), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1001), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1000), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n956), .B1(new_n1242), .B2(new_n998), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n1239), .A3(new_n1238), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT61), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1241), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1234), .B1(new_n1169), .B2(new_n1197), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n646), .A2(G213), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1167), .A2(new_n995), .A3(new_n1126), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1197), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1250), .B2(G378), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1203), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT125), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1060), .B1(new_n1254), .B2(KEYINPUT60), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT125), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1257), .B(new_n1203), .C1(new_n1088), .C2(new_n1252), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1224), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1226), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(G384), .A3(new_n1224), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1247), .A2(new_n1251), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1246), .B1(KEYINPUT63), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT63), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1259), .A2(G384), .A3(new_n1224), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G384), .B1(new_n1259), .B2(new_n1224), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT126), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n646), .A2(G213), .A3(G2897), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1270), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1263), .A2(KEYINPUT126), .A3(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1198), .A2(G378), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1251), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1263), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1275), .A2(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1266), .B1(new_n1274), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1265), .B1(new_n1280), .B2(new_n1264), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n1247), .A2(new_n1251), .B1(KEYINPUT126), .B2(new_n1263), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT62), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n1283), .A2(new_n1284), .B1(new_n1264), .B2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1275), .A2(new_n1277), .A3(new_n1276), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1245), .B1(new_n1287), .B2(KEYINPUT62), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1282), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1281), .A2(new_n1289), .ZN(G405));
  AND3_X1   g1090(.A1(new_n1235), .A2(new_n1263), .A3(new_n1275), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1263), .B1(new_n1235), .B2(new_n1275), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1282), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1282), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1277), .B1(new_n1232), .B2(new_n1247), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1235), .A2(new_n1263), .A3(new_n1275), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1294), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1293), .A2(new_n1297), .ZN(G402));
endmodule


