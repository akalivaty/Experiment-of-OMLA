//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT65), .B1(new_n189), .B2(G134), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G137), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(new_n192), .A3(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n189), .A2(KEYINPUT11), .A3(G134), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n193), .A3(new_n195), .A4(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT81), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G104), .ZN(new_n202));
  OR2_X1    g016(.A1(new_n202), .A2(KEYINPUT80), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(KEYINPUT80), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n207), .A2(G101), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n205), .A2(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT77), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n202), .A2(new_n212), .A3(KEYINPUT3), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n206), .B1(new_n202), .B2(KEYINPUT3), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT78), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n211), .B2(new_n213), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT78), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(new_n215), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n208), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G143), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n224), .B1(new_n226), .B2(KEYINPUT1), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n229));
  INV_X1    g043(.A(G143), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G146), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n225), .A2(KEYINPUT64), .A3(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(G146), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n226), .A2(new_n233), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n228), .A2(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n223), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n207), .A2(G101), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n236), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n241), .B1(new_n227), .B2(new_n235), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n220), .A2(new_n221), .A3(new_n215), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n221), .B1(new_n220), .B2(new_n215), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n240), .B(new_n242), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n200), .B1(new_n239), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT12), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT10), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n237), .A2(new_n249), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n245), .A2(new_n249), .B1(new_n223), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n214), .A2(new_n217), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(G101), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n243), .B2(new_n244), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n253), .A2(new_n252), .A3(G101), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n234), .A2(new_n259), .B1(new_n235), .B2(new_n257), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT79), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT4), .B1(new_n220), .B2(new_n215), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(new_n219), .B2(new_n222), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT79), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n256), .A2(new_n260), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n251), .B(new_n199), .C1(new_n262), .C2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT12), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n269), .B(new_n200), .C1(new_n239), .C2(new_n246), .ZN(new_n270));
  AND2_X1   g084(.A1(KEYINPUT67), .A2(G953), .ZN(new_n271));
  NOR2_X1   g085(.A1(KEYINPUT67), .A2(G953), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G227), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n248), .A2(new_n268), .A3(new_n270), .A4(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n251), .B1(new_n262), .B2(new_n267), .ZN(new_n279));
  INV_X1    g093(.A(new_n199), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n276), .B1(new_n281), .B2(new_n268), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n187), .B(new_n188), .C1(new_n278), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT82), .ZN(new_n284));
  INV_X1    g098(.A(new_n276), .ZN(new_n285));
  INV_X1    g099(.A(new_n268), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n265), .B1(new_n264), .B2(new_n266), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n255), .A2(new_n261), .A3(KEYINPUT79), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n199), .B1(new_n289), .B2(new_n251), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n285), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n291), .B2(new_n277), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT82), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n187), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n281), .A2(new_n268), .A3(new_n276), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n248), .A2(new_n268), .A3(new_n270), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(new_n276), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n188), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n284), .A2(new_n294), .B1(G469), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G140), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G125), .ZN(new_n301));
  INV_X1    g115(.A(G125), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT74), .ZN(new_n305));
  XNOR2_X1  g119(.A(G125), .B(G140), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n308), .A3(new_n225), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n225), .B2(new_n306), .ZN(new_n310));
  OR2_X1    g124(.A1(KEYINPUT67), .A2(G953), .ZN(new_n311));
  INV_X1    g125(.A(G237), .ZN(new_n312));
  NAND2_X1  g126(.A1(KEYINPUT67), .A2(G953), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n311), .A2(G214), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n230), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n273), .A2(G143), .A3(G214), .A4(new_n312), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT18), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n315), .B(new_n316), .C1(new_n317), .C2(new_n198), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n316), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G131), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n310), .B(new_n318), .C1(new_n320), .C2(new_n317), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n198), .B1(new_n315), .B2(new_n316), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT17), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n301), .A2(new_n303), .A3(KEYINPUT16), .ZN(new_n324));
  OR3_X1    g138(.A1(new_n302), .A2(KEYINPUT16), .A3(G140), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G146), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(G146), .B1(new_n324), .B2(new_n325), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT87), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n328), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT87), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(new_n326), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n323), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n315), .A2(new_n316), .A3(new_n198), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n334), .A2(new_n322), .A3(KEYINPUT17), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n321), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G113), .B(G122), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(new_n205), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n338), .B(new_n321), .C1(new_n333), .C2(new_n335), .ZN(new_n341));
  AOI21_X1  g155(.A(G902), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G475), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT20), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT19), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n304), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n305), .A2(new_n308), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(new_n346), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n326), .B1(new_n349), .B2(G146), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n334), .A2(new_n322), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n321), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n339), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n341), .ZN(new_n354));
  NOR2_X1   g168(.A1(G475), .A2(G902), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n345), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n355), .ZN(new_n358));
  AOI211_X1 g172(.A(KEYINPUT20), .B(new_n358), .C1(new_n353), .C2(new_n341), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n344), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT9), .B(G234), .ZN(new_n362));
  INV_X1    g176(.A(G217), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n362), .A2(new_n363), .A3(G953), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n230), .A2(G128), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n224), .A2(G143), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n192), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT88), .B(G122), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G116), .ZN(new_n371));
  INV_X1    g185(.A(G116), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G122), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n371), .A2(new_n201), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n201), .B1(new_n371), .B2(new_n373), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n369), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT13), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT89), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT89), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT13), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n366), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT90), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n367), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT90), .B1(new_n384), .B2(new_n366), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT91), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT92), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n384), .B2(new_n366), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n378), .A2(new_n380), .ZN(new_n389));
  INV_X1    g203(.A(new_n366), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(KEYINPUT92), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n381), .A2(new_n382), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n384), .A2(KEYINPUT90), .A3(new_n366), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT91), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .A4(new_n367), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n386), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n376), .B1(new_n398), .B2(G134), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n368), .B(new_n192), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n371), .A2(new_n201), .A3(new_n373), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XOR2_X1   g216(.A(new_n373), .B(KEYINPUT14), .Z(new_n403));
  AOI21_X1  g217(.A(new_n201), .B1(new_n403), .B2(new_n371), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n365), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n402), .A2(new_n404), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n394), .A2(new_n395), .A3(new_n367), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n392), .B1(new_n408), .B2(KEYINPUT91), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n192), .B1(new_n409), .B2(new_n397), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n407), .B(new_n364), .C1(new_n410), .C2(new_n376), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G478), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(KEYINPUT15), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(KEYINPUT93), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n406), .A2(new_n411), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT93), .A3(new_n188), .ZN(new_n417));
  INV_X1    g231(.A(new_n414), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n412), .A2(KEYINPUT93), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n415), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G953), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G952), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(G234), .B2(G237), .ZN(new_n424));
  AOI211_X1 g238(.A(new_n188), .B(new_n273), .C1(G234), .C2(G237), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(G898), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n361), .A2(new_n421), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  OAI21_X1  g244(.A(G210), .B1(G237), .B2(G902), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT86), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n260), .A2(G125), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(G125), .B2(new_n237), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n422), .A2(G224), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n436), .B(new_n437), .Z(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT83), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n440), .A2(KEYINPUT84), .ZN(new_n441));
  XOR2_X1   g255(.A(G116), .B(G119), .Z(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT2), .B(G113), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n256), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n255), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n442), .A2(new_n443), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G113), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n372), .A2(G119), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(new_n448), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n447), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n223), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n441), .B1(new_n446), .B2(new_n454), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n455), .A2(KEYINPUT6), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n255), .A2(new_n445), .B1(new_n223), .B2(new_n453), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n455), .A2(KEYINPUT6), .B1(new_n457), .B2(new_n439), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n438), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n439), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n437), .A2(KEYINPUT7), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n436), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n436), .A2(KEYINPUT7), .A3(new_n437), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n240), .B1(new_n243), .B2(new_n244), .ZN(new_n465));
  INV_X1    g279(.A(new_n453), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n454), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n439), .B(KEYINPUT85), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT8), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n188), .B1(new_n464), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n434), .B1(new_n459), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n438), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n455), .A2(KEYINPUT6), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n460), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n455), .A2(KEYINPUT6), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n462), .A2(new_n463), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n457), .B2(new_n439), .ZN(new_n481));
  AOI21_X1  g295(.A(G902), .B1(new_n481), .B2(new_n471), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n482), .A3(new_n433), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n474), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n429), .A2(new_n430), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G221), .B1(new_n362), .B2(G902), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT76), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n299), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n190), .A2(new_n195), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n189), .A2(KEYINPUT11), .A3(G134), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT11), .B1(new_n189), .B2(G134), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n198), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n197), .A2(G131), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n260), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n192), .A2(G137), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n189), .A2(G134), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n198), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n238), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n260), .B(KEYINPUT66), .C1(new_n493), .C2(new_n494), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n497), .A2(new_n498), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n495), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n237), .A2(new_n494), .A3(new_n501), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT30), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n444), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n273), .A2(G210), .A3(new_n312), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT27), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT26), .B(G101), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n506), .A2(new_n507), .ZN(new_n515));
  INV_X1    g329(.A(new_n444), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT68), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT68), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n510), .A2(new_n520), .A3(new_n514), .A4(new_n517), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(KEYINPUT31), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n514), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT28), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT69), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n517), .A2(KEYINPUT69), .A3(new_n524), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n497), .A2(new_n503), .A3(new_n504), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n444), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n524), .B1(new_n531), .B2(new_n517), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n523), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n518), .A2(KEYINPUT31), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n522), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G472), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n188), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT32), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT32), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n535), .A2(new_n539), .A3(new_n536), .A4(new_n188), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OR3_X1    g355(.A1(new_n529), .A2(new_n523), .A3(new_n532), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n514), .B1(new_n510), .B2(new_n517), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT70), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT29), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n543), .A2(KEYINPUT70), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n542), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n517), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n515), .A2(new_n516), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n529), .B1(KEYINPUT28), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n523), .A2(new_n545), .ZN(new_n552));
  AOI21_X1  g366(.A(G902), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n536), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n541), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT24), .B(G110), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n224), .A2(G119), .ZN(new_n560));
  INV_X1    g374(.A(G119), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G128), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT71), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n560), .A2(new_n562), .A3(KEYINPUT71), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n557), .A2(new_n558), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n559), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT23), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n561), .B2(G128), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n562), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G110), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT73), .B1(new_n572), .B2(G110), .ZN(new_n576));
  OAI221_X1 g390(.A(new_n568), .B1(new_n327), .B2(new_n328), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n559), .A2(new_n567), .B1(new_n565), .B2(new_n566), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n572), .A2(G110), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n326), .B(new_n309), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n273), .A2(G221), .A3(G234), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT22), .B(G137), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n584), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n577), .A2(new_n580), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n588), .B(new_n188), .C1(new_n363), .C2(G234), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT75), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n363), .B1(G234), .B2(new_n188), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT25), .B1(new_n588), .B2(new_n188), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT25), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n593), .B(G902), .C1(new_n585), .C2(new_n587), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n488), .A2(new_n556), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  NOR2_X1   g412(.A1(new_n299), .A2(new_n487), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n535), .A2(new_n188), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n537), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n603), .A3(new_n596), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n412), .A2(new_n413), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT94), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n406), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n416), .A2(new_n608), .A3(KEYINPUT33), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n406), .B(new_n411), .C1(new_n607), .C2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(G902), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n606), .B1(new_n612), .B2(new_n413), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  OAI22_X1  g428(.A1(new_n356), .A2(new_n359), .B1(new_n343), .B2(new_n342), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n427), .ZN(new_n617));
  INV_X1    g431(.A(new_n430), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n432), .B1(new_n459), .B2(new_n473), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n479), .A2(new_n482), .A3(new_n431), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n605), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT95), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  NOR2_X1   g439(.A1(new_n417), .A2(new_n418), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n416), .A2(new_n188), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT93), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n414), .B1(new_n412), .B2(KEYINPUT93), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n631), .A2(new_n428), .A3(new_n361), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT96), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n605), .A2(new_n621), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NOR2_X1   g450(.A1(new_n586), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n581), .B(new_n637), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n638), .B(new_n188), .C1(new_n363), .C2(G234), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n595), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n488), .A2(new_n603), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT98), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n643), .B(new_n645), .ZN(G12));
  NAND2_X1  g460(.A1(new_n631), .A2(new_n361), .ZN(new_n647));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n424), .B1(new_n425), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n650), .A2(new_n642), .A3(new_n621), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n556), .A2(new_n599), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  NOR4_X1   g467(.A1(new_n361), .A2(new_n640), .A3(new_n421), .A4(new_n618), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n484), .B(new_n657), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n649), .B(KEYINPUT39), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n599), .A2(new_n661), .ZN(new_n662));
  AOI211_X1 g476(.A(new_n656), .B(new_n660), .C1(KEYINPUT40), .C2(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(KEYINPUT40), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n550), .A2(new_n523), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(KEYINPUT100), .Z(new_n666));
  NAND2_X1  g480(.A1(new_n519), .A2(new_n521), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n188), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G472), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n541), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT101), .Z(new_n671));
  NOR2_X1   g485(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n230), .ZN(G45));
  NOR3_X1   g487(.A1(new_n613), .A2(new_n361), .A3(new_n649), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n642), .A2(new_n621), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n556), .A2(new_n599), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  NAND2_X1  g491(.A1(new_n284), .A2(new_n294), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n292), .A2(new_n187), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n678), .A2(new_n486), .A3(new_n621), .A4(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n556), .A2(new_n680), .A3(new_n596), .A4(new_n617), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT103), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT41), .B(G113), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NAND4_X1  g498(.A1(new_n556), .A2(new_n680), .A3(new_n633), .A4(new_n596), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NAND4_X1  g500(.A1(new_n678), .A2(new_n486), .A3(new_n621), .A4(new_n679), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n642), .A2(new_n429), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n556), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  NAND4_X1  g505(.A1(new_n678), .A2(new_n486), .A3(new_n428), .A4(new_n679), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n522), .B(new_n534), .C1(new_n551), .C2(new_n514), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n536), .A3(new_n188), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n601), .A2(new_n596), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n631), .B2(new_n615), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n630), .A2(new_n629), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n697), .A2(new_n615), .A3(new_n699), .A4(new_n415), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n621), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT105), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n621), .B(new_n703), .C1(new_n698), .C2(new_n700), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n696), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  NAND4_X1  g521(.A1(new_n601), .A2(new_n640), .A3(new_n694), .A4(new_n674), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n687), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n302), .ZN(G27));
  NAND2_X1  g524(.A1(new_n541), .A2(KEYINPUT106), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n538), .A2(new_n712), .A3(new_n540), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n711), .A2(new_n555), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n674), .A2(KEYINPUT42), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n474), .A2(new_n483), .A3(new_n486), .A4(new_n430), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n299), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n714), .A2(new_n596), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n299), .A2(new_n716), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n556), .A2(new_n596), .A3(new_n674), .A4(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G131), .ZN(G33));
  NAND4_X1  g538(.A1(new_n556), .A2(new_n596), .A3(new_n650), .A4(new_n719), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G134), .ZN(G36));
  NOR2_X1   g540(.A1(new_n613), .A2(new_n615), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT43), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n602), .A3(new_n640), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n729), .B(KEYINPUT44), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n297), .B(KEYINPUT45), .ZN(new_n731));
  OAI21_X1  g545(.A(G469), .B1(new_n731), .B2(G902), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n678), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n486), .A3(new_n661), .ZN(new_n736));
  OR4_X1    g550(.A1(new_n618), .A2(new_n730), .A3(new_n484), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT107), .B(G137), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G39));
  NAND2_X1  g553(.A1(new_n735), .A2(new_n486), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT108), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n741), .A2(KEYINPUT108), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n744), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n740), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n554), .B1(new_n538), .B2(new_n540), .ZN(new_n749));
  INV_X1    g563(.A(new_n596), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n484), .A2(new_n618), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n749), .A2(new_n750), .A3(new_n674), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  INV_X1    g569(.A(new_n487), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n596), .A2(new_n756), .A3(new_n430), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT109), .ZN(new_n758));
  INV_X1    g572(.A(new_n658), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n759), .A3(new_n727), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n678), .A2(new_n679), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n760), .B1(KEYINPUT49), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n762), .B(new_n671), .C1(KEYINPUT49), .C2(new_n761), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n761), .A2(new_n716), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n671), .A2(new_n596), .A3(new_n424), .A4(new_n764), .ZN(new_n765));
  OR3_X1    g579(.A1(new_n765), .A2(new_n615), .A3(new_n614), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n728), .A2(new_n424), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n695), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n678), .A2(new_n486), .A3(new_n679), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n658), .A2(new_n430), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n767), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n769), .A2(KEYINPUT50), .A3(new_n772), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n601), .A2(new_n640), .A3(new_n694), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n764), .A2(new_n424), .A3(new_n728), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n766), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n761), .A2(new_n756), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n751), .B(new_n769), .C1(new_n748), .C2(new_n781), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n780), .A2(KEYINPUT51), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT51), .B1(new_n780), .B2(new_n782), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n423), .B(KEYINPUT114), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n770), .A2(new_n687), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI221_X1 g602(.A(new_n788), .B1(new_n787), .B2(new_n786), .C1(new_n765), .C2(new_n616), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n554), .B1(new_n541), .B2(KEYINPUT106), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n750), .B1(new_n790), .B2(new_n713), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n778), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT48), .Z(new_n793));
  OR2_X1    g607(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n783), .A2(new_n784), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n640), .A2(new_n649), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(KEYINPUT110), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n486), .B1(new_n796), .B2(KEYINPUT110), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n299), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n705), .A2(new_n799), .A3(new_n670), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n680), .A2(new_n776), .A3(new_n674), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n800), .A2(new_n652), .A3(new_n676), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n298), .A2(G469), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n283), .A2(KEYINPUT82), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n293), .B1(new_n292), .B2(new_n187), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n756), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n749), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n709), .B1(new_n810), .B2(new_n651), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(KEYINPUT52), .A3(new_n676), .A4(new_n800), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n804), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n681), .A2(new_n685), .A3(new_n706), .A4(new_n690), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT112), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n705), .A2(new_n696), .B1(new_n689), .B2(new_n556), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n681), .A4(new_n685), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n649), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n361), .A2(new_n642), .A3(new_n421), .A4(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n556), .A2(new_n599), .A3(new_n821), .A4(new_n751), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n719), .A2(new_n776), .A3(new_n674), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n725), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n484), .A2(new_n430), .A3(new_n428), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n616), .B2(new_n647), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n599), .A2(new_n603), .A3(new_n826), .A4(new_n596), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n597), .A2(new_n643), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n723), .A2(new_n824), .A3(KEYINPUT53), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n819), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n597), .A2(new_n643), .A3(new_n827), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n814), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n725), .A2(new_n822), .A3(new_n823), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n722), .B2(new_n718), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n813), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n813), .A2(new_n830), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n835), .A2(new_n836), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n804), .A2(new_n812), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n681), .A2(new_n685), .A3(new_n706), .A4(new_n690), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n723), .A3(new_n828), .A4(new_n824), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n836), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n842), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n835), .A2(KEYINPUT111), .A3(new_n836), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT54), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n795), .A2(new_n841), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(G952), .A2(G953), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n763), .B1(new_n852), .B2(new_n853), .ZN(G75));
  AOI22_X1  g668(.A1(new_n791), .A2(new_n717), .B1(new_n720), .B2(new_n721), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n597), .A2(new_n643), .A3(new_n827), .A4(KEYINPUT53), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n855), .A2(new_n833), .A3(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n813), .A3(new_n815), .A4(new_n818), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n847), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n859), .A2(G210), .A3(G902), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT56), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n477), .A2(new_n475), .A3(new_n478), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n459), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n861), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n864), .B1(new_n860), .B2(KEYINPUT56), .ZN(new_n867));
  XOR2_X1   g681(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n868));
  AND3_X1   g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n866), .B2(new_n867), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n273), .A2(G952), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(G51));
  NAND2_X1  g686(.A1(new_n859), .A2(KEYINPUT54), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n839), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(G469), .A2(G902), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT57), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n874), .A2(new_n877), .B1(new_n291), .B2(new_n277), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n878), .A2(KEYINPUT117), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n837), .A2(new_n188), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n880), .A2(G469), .A3(new_n731), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n878), .B2(KEYINPUT117), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n871), .B1(new_n879), .B2(new_n882), .ZN(G54));
  NAND3_X1  g697(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n884));
  INV_X1    g698(.A(new_n354), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n871), .ZN(G60));
  NAND2_X1  g702(.A1(new_n841), .A2(new_n851), .ZN(new_n889));
  NAND2_X1  g703(.A1(G478), .A2(G902), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT59), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n609), .A2(new_n611), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n891), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n839), .B2(new_n873), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT118), .ZN(new_n897));
  OR3_X1    g711(.A1(new_n896), .A2(new_n897), .A3(new_n871), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n897), .B1(new_n896), .B2(new_n871), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n892), .A2(new_n894), .B1(new_n898), .B2(new_n899), .ZN(G63));
  XOR2_X1   g714(.A(new_n588), .B(KEYINPUT121), .Z(new_n901));
  NAND2_X1  g715(.A1(G217), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT120), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT60), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n901), .B1(new_n837), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n847), .B2(new_n858), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n638), .ZN(new_n908));
  INV_X1    g722(.A(new_n871), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n906), .A2(new_n908), .A3(KEYINPUT61), .A4(new_n909), .ZN(new_n910));
  XOR2_X1   g724(.A(KEYINPUT119), .B(KEYINPUT61), .Z(new_n911));
  INV_X1    g725(.A(new_n901), .ZN(new_n912));
  OAI211_X1 g726(.A(KEYINPUT122), .B(new_n909), .C1(new_n907), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n908), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT122), .B1(new_n906), .B2(new_n909), .ZN(new_n915));
  OAI211_X1 g729(.A(KEYINPUT123), .B(new_n911), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n909), .B1(new_n907), .B2(new_n912), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n913), .A3(new_n908), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT123), .B1(new_n921), .B2(new_n911), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n910), .B1(new_n917), .B2(new_n922), .ZN(G66));
  INV_X1    g737(.A(G224), .ZN(new_n924));
  OAI21_X1  g738(.A(G953), .B1(new_n426), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n273), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n832), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n456), .B(new_n458), .C1(G898), .C2(new_n273), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(G69));
  XNOR2_X1  g743(.A(new_n509), .B(new_n349), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n616), .A2(new_n647), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n751), .ZN(new_n932));
  NOR4_X1   g746(.A1(new_n662), .A2(new_n749), .A3(new_n750), .A4(new_n932), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT124), .Z(new_n934));
  NAND3_X1  g748(.A1(new_n754), .A2(new_n737), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n811), .A2(new_n676), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n672), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n930), .B1(new_n940), .B2(new_n926), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n754), .A2(new_n737), .A3(new_n723), .ZN(new_n942));
  INV_X1    g756(.A(new_n705), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n736), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n791), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n945), .A2(new_n676), .A3(new_n725), .A4(new_n811), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n273), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n273), .A2(G900), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT125), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n930), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n941), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n273), .B1(G227), .B2(G900), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n930), .B2(KEYINPUT126), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n953), .B(new_n956), .ZN(G72));
  AND3_X1   g771(.A1(new_n510), .A2(new_n523), .A3(new_n517), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n523), .B1(new_n510), .B2(new_n517), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT63), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT127), .Z(new_n963));
  AOI21_X1  g777(.A(new_n871), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n942), .A2(new_n946), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n940), .A2(new_n959), .B1(new_n965), .B2(new_n958), .ZN(new_n966));
  INV_X1    g780(.A(new_n832), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n546), .A2(new_n544), .ZN(new_n969));
  INV_X1    g783(.A(new_n667), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n962), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n968), .B1(new_n850), .B2(new_n971), .ZN(G57));
endmodule


