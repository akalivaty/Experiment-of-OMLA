//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XOR2_X1   g0008(.A(KEYINPUT66), .B(G244), .Z(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G107), .A2(G264), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n208), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  INV_X1    g0018(.A(new_n208), .ZN(new_n219));
  INV_X1    g0019(.A(G13), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n219), .A2(KEYINPUT65), .A3(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT65), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n222), .B1(new_n208), .B2(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n204), .A2(new_n205), .ZN(new_n230));
  INV_X1    g0030(.A(G50), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n218), .B(new_n226), .C1(new_n229), .C2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT67), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n231), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n203), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G45), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n254), .A2(new_n255), .A3(G274), .A4(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n266), .A2(G223), .B1(new_n269), .B2(G77), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n264), .A2(new_n265), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G222), .A3(new_n261), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n260), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OR2_X1    g0075(.A1(KEYINPUT68), .A2(G1), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT68), .A2(G1), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n258), .A3(new_n277), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n278), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n279));
  AOI21_X1  g0079(.A(KEYINPUT69), .B1(new_n278), .B2(new_n254), .ZN(new_n280));
  OAI21_X1  g0080(.A(G226), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G200), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT75), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT10), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(new_n285), .B2(new_n284), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n227), .B1(new_n208), .B2(new_n263), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT70), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(new_n263), .B2(G20), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n228), .A2(KEYINPUT70), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT8), .B(G58), .ZN(new_n294));
  INV_X1    g0094(.A(G150), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n228), .A2(new_n263), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n228), .B1(new_n230), .B2(new_n231), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n288), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n276), .A2(G13), .A3(G20), .A4(new_n277), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT71), .ZN(new_n301));
  AND2_X1   g0101(.A1(KEYINPUT68), .A2(G1), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT68), .A2(G1), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT71), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(G13), .A4(G20), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n231), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n301), .A2(new_n306), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n276), .A2(new_n277), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n228), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n288), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n309), .A2(G50), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n299), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n299), .A2(new_n308), .A3(new_n314), .A4(KEYINPUT74), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT9), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(KEYINPUT9), .A3(new_n318), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n275), .A2(G190), .A3(new_n281), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n287), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(KEYINPUT76), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT76), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n321), .A2(new_n327), .A3(new_n322), .A4(new_n323), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n328), .A3(new_n283), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n325), .B1(new_n329), .B2(KEYINPUT10), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n301), .A2(new_n306), .A3(new_n203), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT12), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n210), .B1(new_n290), .B2(new_n291), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n296), .A2(new_n231), .B1(new_n228), .B2(G68), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n288), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT77), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT77), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(new_n288), .C1(new_n333), .C2(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT11), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT11), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(new_n341), .A3(new_n338), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n332), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G238), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT69), .ZN(new_n345));
  NOR2_X1   g0145(.A1(G41), .A2(G45), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n302), .A2(new_n303), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n345), .B1(new_n347), .B2(new_n274), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n278), .A2(KEYINPUT69), .A3(new_n254), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(G226), .A2(G1698), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n236), .B2(G1698), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n271), .B1(G33), .B2(G97), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n259), .B1(new_n353), .B2(new_n254), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT13), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(G238), .B1(new_n279), .B2(new_n280), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G97), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n236), .A2(G1698), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G226), .B2(G1698), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n358), .B1(new_n360), .B2(new_n269), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n260), .B1(new_n361), .B2(new_n274), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n356), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G200), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT73), .B1(new_n309), .B2(new_n313), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT73), .ZN(new_n367));
  AOI211_X1 g0167(.A(new_n367), .B(new_n288), .C1(new_n301), .C2(new_n306), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n311), .A2(new_n203), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n355), .A2(G190), .A3(new_n363), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n343), .A2(new_n365), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n209), .B1(new_n348), .B2(new_n349), .ZN(new_n374));
  INV_X1    g0174(.A(G107), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n269), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(G232), .A2(G1698), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n344), .B2(G1698), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n376), .B(new_n274), .C1(new_n269), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n259), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n374), .A2(new_n380), .A3(G179), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n374), .A2(new_n380), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G169), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n309), .A2(new_n313), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n367), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n309), .A2(KEYINPUT73), .A3(new_n313), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n387), .A2(G77), .A3(new_n312), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n294), .ZN(new_n390));
  INV_X1    g0190(.A(new_n296), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n390), .A2(new_n391), .B1(G20), .B2(G77), .ZN(new_n392));
  XOR2_X1   g0192(.A(KEYINPUT15), .B(G87), .Z(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n292), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n313), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n307), .A2(KEYINPUT72), .A3(new_n210), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT72), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n309), .B2(G77), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n395), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n389), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n385), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n383), .A2(G200), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n382), .A2(G190), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n389), .A4(new_n399), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n282), .A2(new_n384), .ZN(new_n405));
  INV_X1    g0205(.A(G179), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n275), .A2(new_n406), .A3(new_n281), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n405), .A2(new_n315), .A3(new_n407), .ZN(new_n408));
  AND4_X1   g0208(.A1(new_n373), .A2(new_n401), .A3(new_n404), .A4(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n274), .B1(new_n304), .B2(new_n258), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n260), .B1(G232), .B2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(G223), .B(new_n261), .C1(new_n267), .C2(new_n268), .ZN(new_n412));
  OAI211_X1 g0212(.A(G226), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n413));
  INV_X1    g0213(.A(G87), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n412), .B(new_n413), .C1(new_n263), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n274), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n411), .A2(G179), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n384), .B1(new_n411), .B2(new_n416), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G58), .A2(G68), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n204), .A2(new_n205), .A3(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(G20), .B1(G159), .B2(new_n391), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n264), .A2(new_n228), .A3(new_n265), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT7), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n228), .A4(new_n265), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n203), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT78), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n423), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI211_X1 g0230(.A(KEYINPUT78), .B(new_n203), .C1(new_n426), .C2(new_n427), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n420), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n422), .A2(G20), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n391), .A2(G159), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n313), .B1(new_n436), .B2(KEYINPUT16), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n386), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n311), .A2(new_n294), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n439), .A2(new_n440), .B1(new_n307), .B2(new_n294), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n419), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT18), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT7), .B1(new_n269), .B2(new_n228), .ZN(new_n445));
  INV_X1    g0245(.A(new_n427), .ZN(new_n446));
  OAI21_X1  g0246(.A(G68), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n435), .B1(new_n447), .B2(KEYINPUT78), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n428), .A2(new_n429), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT16), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(KEYINPUT16), .A3(new_n423), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n288), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n441), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n419), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n453), .A2(new_n454), .A3(new_n443), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n444), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G190), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n411), .A2(new_n457), .A3(new_n416), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n411), .A2(new_n416), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(G200), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n438), .A2(new_n460), .A3(new_n441), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT17), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n343), .A2(new_n371), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT14), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n350), .A2(new_n354), .A3(KEYINPUT13), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n357), .B1(new_n356), .B2(new_n362), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n464), .B(G169), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n355), .A2(G179), .A3(new_n363), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n464), .B1(new_n364), .B2(G169), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n409), .A2(new_n456), .A3(new_n462), .A4(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT79), .B1(new_n330), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n472), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT79), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT10), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n284), .B1(new_n324), .B2(KEYINPUT76), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(new_n328), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n474), .B(new_n475), .C1(new_n478), .C2(new_n325), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n304), .A2(G33), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n439), .A2(G97), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT6), .ZN(new_n484));
  INV_X1    g0284(.A(G97), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n484), .A2(new_n485), .A3(G107), .ZN(new_n486));
  XNOR2_X1  g0286(.A(G97), .B(G107), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n488), .A2(new_n228), .B1(new_n210), .B2(new_n296), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n375), .B1(new_n426), .B2(new_n427), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n288), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n307), .A2(new_n485), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n483), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n310), .A2(new_n257), .ZN(new_n494));
  XOR2_X1   g0294(.A(KEYINPUT5), .B(G41), .Z(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n494), .A2(new_n496), .A3(G274), .A4(new_n254), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n304), .A2(G45), .ZN(new_n498));
  OAI211_X1 g0298(.A(G257), .B(new_n254), .C1(new_n498), .C2(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(G244), .B(new_n261), .C1(new_n267), .C2(new_n268), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT80), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT80), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(G250), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G283), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT81), .ZN(new_n511));
  OAI21_X1  g0311(.A(G244), .B1(new_n267), .B2(new_n268), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n502), .A2(G1698), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n511), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n271), .A2(KEYINPUT81), .A3(G244), .A4(new_n513), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT82), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n254), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n507), .A2(KEYINPUT82), .A3(new_n517), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n500), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n493), .B1(new_n522), .B2(G190), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT83), .ZN(new_n524));
  OAI21_X1  g0324(.A(G200), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n515), .A2(new_n516), .ZN(new_n526));
  INV_X1    g0326(.A(new_n510), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n501), .A2(new_n505), .A3(new_n502), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n505), .B1(new_n501), .B2(new_n502), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n519), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n274), .A3(new_n521), .ZN(new_n533));
  INV_X1    g0333(.A(new_n500), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(KEYINPUT83), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n523), .B1(new_n525), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n384), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n522), .A2(new_n406), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n539), .A3(new_n493), .ZN(new_n540));
  INV_X1    g0340(.A(new_n393), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n307), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n309), .A2(G87), .A3(new_n313), .A4(new_n482), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT19), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n228), .B1(new_n358), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n414), .A2(new_n485), .A3(new_n375), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n271), .A2(new_n228), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(new_n203), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n485), .B1(new_n290), .B2(new_n291), .ZN(new_n550));
  OR3_X1    g0350(.A1(new_n550), .A2(KEYINPUT84), .A3(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT84), .B1(new_n550), .B2(KEYINPUT19), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n542), .B(new_n543), .C1(new_n553), .C2(new_n313), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G200), .ZN(new_n556));
  OAI211_X1 g0356(.A(G238), .B(new_n261), .C1(new_n267), .C2(new_n268), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G116), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n558), .C1(new_n512), .C2(new_n261), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n274), .ZN(new_n560));
  INV_X1    g0360(.A(G274), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n304), .A2(G45), .A3(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n254), .B(new_n562), .C1(new_n494), .C2(G250), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n556), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n560), .A2(new_n563), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(G190), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n309), .A2(new_n313), .A3(new_n393), .A4(new_n482), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n542), .B(new_n567), .C1(new_n553), .C2(new_n313), .ZN(new_n568));
  AOI21_X1  g0368(.A(G169), .B1(new_n560), .B2(new_n563), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n406), .B2(new_n565), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n555), .A2(new_n566), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n537), .A2(new_n540), .A3(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n509), .B(new_n228), .C1(G33), .C2(new_n485), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n573), .B(new_n288), .C1(new_n228), .C2(G116), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT20), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(G116), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n307), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n577), .B1(new_n304), .B2(G33), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n579), .B1(new_n369), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G264), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n582));
  OAI211_X1 g0382(.A(G257), .B(new_n261), .C1(new_n267), .C2(new_n268), .ZN(new_n583));
  XNOR2_X1  g0383(.A(KEYINPUT85), .B(G303), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n583), .C1(new_n271), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n274), .ZN(new_n586));
  OAI211_X1 g0386(.A(G270), .B(new_n254), .C1(new_n498), .C2(new_n495), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(G179), .A3(new_n497), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n497), .A3(new_n587), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(KEYINPUT21), .A3(G169), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n581), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(G169), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n387), .A2(new_n388), .A3(new_n580), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n576), .A2(new_n578), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT86), .B1(new_n595), .B2(KEYINPUT21), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT86), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(new_n598), .C1(new_n581), .C2(new_n592), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n591), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g0400(.A(KEYINPUT87), .B(KEYINPUT22), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n548), .B2(new_n414), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT22), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(KEYINPUT87), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n271), .A2(new_n228), .A3(G87), .A4(new_n604), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n263), .A2(new_n577), .A3(G20), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT23), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n228), .B2(G107), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n375), .A2(KEYINPUT23), .A3(G20), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n606), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n602), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT24), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT24), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n602), .A2(new_n613), .A3(new_n605), .A4(new_n610), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n313), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n386), .B1(G33), .B2(new_n304), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT25), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n309), .B2(G107), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n307), .A2(KEYINPUT25), .A3(new_n375), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n617), .A2(G107), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(G257), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n622));
  OAI211_X1 g0422(.A(G250), .B(new_n261), .C1(new_n267), .C2(new_n268), .ZN(new_n623));
  INV_X1    g0423(.A(G294), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n622), .B(new_n623), .C1(new_n263), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n274), .ZN(new_n626));
  OAI211_X1 g0426(.A(G264), .B(new_n254), .C1(new_n498), .C2(new_n495), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n497), .A3(new_n627), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n628), .A2(new_n457), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(G200), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n616), .A2(new_n621), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n384), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n628), .A2(G179), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n620), .A2(new_n619), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n439), .A2(new_n482), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(new_n375), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n632), .B(new_n633), .C1(new_n636), .C2(new_n615), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n589), .A2(G200), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n581), .B(new_n639), .C1(new_n457), .C2(new_n589), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n600), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n481), .A2(new_n572), .A3(new_n641), .ZN(G372));
  INV_X1    g0442(.A(new_n408), .ZN(new_n643));
  INV_X1    g0443(.A(new_n330), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT89), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n401), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n385), .A2(new_n400), .A3(KEYINPUT89), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n373), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n648), .A2(new_n471), .ZN(new_n649));
  INV_X1    g0449(.A(new_n462), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n456), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n643), .B1(new_n644), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n537), .A2(new_n540), .A3(new_n571), .ZN(new_n653));
  INV_X1    g0453(.A(new_n631), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n600), .B2(new_n637), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n653), .A2(new_n655), .B1(new_n568), .B2(new_n570), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n571), .A2(new_n538), .A3(new_n539), .A4(new_n493), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT88), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n658), .B1(new_n657), .B2(new_n659), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n661), .A2(new_n662), .B1(new_n659), .B2(new_n657), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n652), .B1(new_n481), .B2(new_n665), .ZN(G369));
  NAND2_X1  g0466(.A1(new_n596), .A2(new_n599), .ZN(new_n667));
  INV_X1    g0467(.A(new_n591), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n220), .A2(G20), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT27), .B1(new_n310), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n304), .A2(new_n673), .A3(new_n670), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n672), .A2(G213), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G343), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT90), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n581), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n669), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n680), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n600), .A2(new_n640), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT91), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT91), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n681), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n678), .B1(new_n636), .B2(new_n615), .ZN(new_n688));
  INV_X1    g0488(.A(new_n637), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n638), .A2(new_n688), .B1(new_n689), .B2(new_n678), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n685), .A2(G330), .A3(new_n687), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n631), .A2(new_n637), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n600), .A2(new_n693), .A3(new_n678), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n637), .A2(new_n678), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT92), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n669), .A2(new_n638), .A3(new_n679), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT92), .ZN(new_n698));
  INV_X1    g0498(.A(new_n695), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n692), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n224), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n546), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n232), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n707), .B(KEYINPUT93), .C1(new_n708), .C2(new_n705), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(KEYINPUT93), .B2(new_n707), .ZN(new_n710));
  XOR2_X1   g0510(.A(new_n710), .B(KEYINPUT28), .Z(new_n711));
  OAI21_X1  g0511(.A(new_n631), .B1(new_n669), .B2(new_n689), .ZN(new_n712));
  INV_X1    g0512(.A(new_n568), .ZN(new_n713));
  INV_X1    g0513(.A(new_n570), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n712), .A2(new_n572), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT96), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n657), .A2(new_n716), .A3(new_n659), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n657), .A2(new_n659), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n716), .B1(new_n657), .B2(new_n659), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT29), .B(new_n679), .C1(new_n715), .C2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n678), .B1(new_n656), .B2(new_n663), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(KEYINPUT29), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(G179), .B1(new_n560), .B2(new_n563), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n628), .A3(new_n589), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT95), .B1(new_n522), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n626), .A2(new_n560), .A3(new_n563), .A4(new_n627), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n588), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n533), .A2(new_n534), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT95), .ZN(new_n733));
  INV_X1    g0533(.A(new_n726), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n535), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n522), .A2(KEYINPUT30), .A3(new_n729), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n727), .A2(new_n732), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n678), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n535), .A2(new_n734), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n732), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n679), .A2(new_n739), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n738), .A2(new_n739), .B1(new_n743), .B2(KEYINPUT94), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n743), .A2(KEYINPUT94), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n572), .A2(new_n641), .A3(new_n678), .ZN(new_n747));
  OAI21_X1  g0547(.A(G330), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n724), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n711), .B1(new_n750), .B2(G1), .ZN(G364));
  NAND2_X1  g0551(.A1(new_n685), .A2(new_n687), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n255), .B1(new_n670), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OR3_X1    g0558(.A1(new_n704), .A2(KEYINPUT97), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT97), .B1(new_n704), .B2(new_n758), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n224), .A2(G355), .A3(new_n271), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n703), .A2(new_n271), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G45), .B2(new_n708), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n251), .A2(new_n257), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n762), .B1(G116), .B2(new_n224), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n227), .B1(G20), .B2(new_n384), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n755), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n761), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n767), .ZN(new_n770));
  NAND3_X1  g0570(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G179), .A2(G200), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n228), .B1(new_n774), .B2(G190), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n773), .A2(new_n203), .B1(new_n775), .B2(new_n485), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n228), .A2(new_n457), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n406), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n269), .B1(new_n779), .B2(G87), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT32), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n228), .A2(G190), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n774), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(new_n406), .A3(G200), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT99), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n780), .B1(new_n781), .B2(new_n785), .C1(new_n788), .C2(new_n375), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n776), .B(new_n789), .C1(new_n781), .C2(new_n785), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n406), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n777), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n782), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G58), .A2(new_n793), .B1(new_n795), .B2(G77), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n771), .A2(new_n457), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n796), .B1(new_n231), .B2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT98), .Z(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n269), .B1(new_n775), .B2(new_n624), .C1(new_n778), .C2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G326), .B2(new_n797), .ZN(new_n803));
  INV_X1    g0603(.A(G322), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n792), .A2(new_n804), .B1(new_n794), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n783), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(G329), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n773), .B1(KEYINPUT100), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(KEYINPUT100), .B2(new_n810), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G283), .B2(new_n787), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n790), .A2(new_n800), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n756), .B(new_n769), .C1(new_n770), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G330), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n752), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n685), .A2(G330), .A3(new_n687), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n818), .A2(new_n819), .A3(new_n761), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n816), .A2(new_n820), .ZN(G396));
  NAND2_X1  g0621(.A1(new_n400), .A2(new_n678), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n646), .B2(new_n647), .ZN(new_n823));
  INV_X1    g0623(.A(new_n822), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(new_n401), .B2(new_n404), .ZN(new_n825));
  OAI21_X1  g0625(.A(KEYINPUT102), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n647), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT89), .B1(new_n385), .B2(new_n400), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n401), .ZN(new_n830));
  INV_X1    g0630(.A(new_n404), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n822), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT102), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n829), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n826), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n657), .A2(new_n659), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT88), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n719), .B1(new_n838), .B2(new_n660), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n836), .B(new_n679), .C1(new_n715), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n723), .B2(new_n836), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n761), .B1(new_n841), .B2(new_n748), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n748), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(KEYINPUT103), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(KEYINPUT103), .B2(new_n843), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n767), .A2(new_n753), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n761), .B1(new_n210), .B2(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G143), .A2(new_n793), .B1(new_n795), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n798), .B2(new_n849), .C1(new_n295), .C2(new_n773), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT34), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n788), .A2(new_n203), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n775), .A2(new_n202), .ZN(new_n854));
  INV_X1    g0654(.A(G132), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n271), .B1(new_n783), .B2(new_n855), .C1(new_n778), .C2(new_n231), .ZN(new_n856));
  NOR4_X1   g0656(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n850), .A2(new_n851), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n792), .A2(new_n624), .B1(new_n775), .B2(new_n485), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT101), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n788), .A2(new_n414), .ZN(new_n861));
  INV_X1    g0661(.A(G283), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n773), .A2(new_n862), .B1(new_n798), .B2(new_n801), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n269), .B1(new_n783), .B2(new_n805), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n778), .A2(new_n375), .B1(new_n794), .B2(new_n577), .ZN(new_n865));
  NOR4_X1   g0665(.A1(new_n861), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n857), .A2(new_n858), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n847), .B1(new_n770), .B2(new_n867), .C1(new_n836), .C2(new_n754), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n845), .A2(new_n868), .ZN(G384));
  NOR2_X1   g0669(.A1(new_n436), .A2(KEYINPUT16), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n441), .B1(new_n452), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n675), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n456), .B2(new_n462), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n453), .A2(new_n454), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n453), .A2(new_n675), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n461), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n878), .A2(KEYINPUT108), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(KEYINPUT108), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n871), .B1(new_n454), .B2(new_n675), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n877), .B1(new_n882), .B2(new_n461), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n874), .B(KEYINPUT38), .C1(new_n881), .C2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n438), .A2(new_n441), .A3(new_n460), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(new_n442), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT108), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(new_n877), .A4(new_n876), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n878), .A2(KEYINPUT108), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n885), .B1(new_n891), .B2(new_n873), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n884), .A2(new_n892), .A3(KEYINPUT39), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n887), .A2(new_n876), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n889), .A2(new_n890), .B1(new_n895), .B2(KEYINPUT37), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n876), .B1(new_n456), .B2(new_n462), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n885), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT39), .B1(new_n884), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n471), .A2(KEYINPUT106), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT106), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n463), .B(new_n902), .C1(new_n469), .C2(new_n470), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n678), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n371), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n332), .A2(new_n340), .A3(new_n342), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n678), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n373), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n901), .A2(new_n903), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT107), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n901), .A2(new_n909), .A3(KEYINPUT107), .A4(new_n903), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n471), .A2(new_n679), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n830), .A2(new_n679), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT105), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n916), .B1(new_n840), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n884), .A2(new_n892), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n456), .A2(new_n675), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n905), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n480), .B(new_n722), .C1(KEYINPUT29), .C2(new_n723), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n652), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n924), .B(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT110), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n738), .A2(KEYINPUT109), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT109), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n737), .A2(new_n930), .A3(new_n678), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n739), .A3(new_n931), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n600), .A2(new_n638), .A3(new_n640), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n653), .A2(new_n933), .A3(new_n679), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n737), .A2(new_n742), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n914), .A2(new_n915), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n937), .A3(new_n836), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n879), .B2(new_n880), .ZN(new_n940));
  INV_X1    g0740(.A(new_n897), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT38), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n891), .A2(new_n885), .A3(new_n873), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT40), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n928), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n884), .B2(new_n898), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n835), .B1(new_n914), .B2(new_n915), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n947), .A2(KEYINPUT110), .A3(new_n936), .A4(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n921), .A2(new_n948), .A3(new_n936), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n945), .A2(new_n949), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n480), .A2(new_n936), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n817), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n927), .A2(new_n954), .B1(new_n310), .B2(new_n671), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n927), .B2(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT35), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n488), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n229), .A2(G116), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n488), .B2(new_n957), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(new_n961), .B2(KEYINPUT104), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(KEYINPUT104), .B2(new_n961), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT36), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n421), .A2(G77), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n247), .B1(new_n708), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(new_n220), .A3(new_n310), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n956), .A2(new_n964), .A3(new_n967), .ZN(G367));
  NAND2_X1  g0768(.A1(new_n678), .A2(new_n554), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n571), .B(new_n969), .Z(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n540), .A2(new_n679), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n535), .A2(KEYINPUT83), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n522), .A2(new_n524), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n976), .A3(G200), .ZN(new_n977));
  INV_X1    g0777(.A(new_n493), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n535), .B2(new_n384), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n977), .A2(new_n523), .B1(new_n979), .B2(new_n539), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n678), .A2(new_n493), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n974), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OR3_X1    g0782(.A1(new_n692), .A2(KEYINPUT111), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT111), .B1(new_n692), .B2(new_n982), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n973), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n973), .A3(new_n984), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n537), .A2(new_n689), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n678), .B1(new_n989), .B2(new_n540), .ZN(new_n990));
  INV_X1    g0790(.A(new_n982), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n694), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n990), .B1(new_n992), .B2(KEYINPUT42), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(KEYINPUT42), .B2(new_n992), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n986), .A2(new_n987), .B1(new_n988), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n987), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n988), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n996), .A2(new_n997), .A3(new_n985), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n704), .B(KEYINPUT41), .Z(new_n1000));
  INV_X1    g0800(.A(KEYINPUT45), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT112), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n701), .B2(new_n991), .ZN(new_n1003));
  AOI211_X1 g0803(.A(KEYINPUT112), .B(new_n982), .C1(new_n696), .C2(new_n700), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n694), .A2(KEYINPUT92), .A3(new_n695), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n698), .B1(new_n697), .B2(new_n699), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n991), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(KEYINPUT112), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n701), .A2(new_n1002), .A3(new_n991), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1009), .A2(KEYINPUT45), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n696), .A2(new_n700), .A3(new_n982), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT44), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1005), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n692), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n600), .A2(new_n678), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n697), .B1(new_n691), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n819), .B(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n749), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1005), .A2(new_n1011), .A3(new_n1014), .A4(new_n692), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1017), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1000), .B1(new_n1023), .B2(new_n750), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n999), .B1(new_n1024), .B2(new_n758), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT113), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g0827(.A(KEYINPUT113), .B(new_n999), .C1(new_n1024), .C2(new_n758), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n970), .A2(new_n755), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n761), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n763), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(new_n242), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n768), .B1(new_n224), .B2(new_n541), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n210), .A2(new_n786), .B1(new_n792), .B2(new_n295), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n271), .B1(new_n778), .B2(new_n202), .C1(new_n784), .C2(new_n773), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n794), .A2(new_n231), .B1(new_n783), .B2(new_n849), .ZN(new_n1038));
  INV_X1    g0838(.A(G143), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n798), .A2(new_n1039), .B1(new_n775), .B2(new_n203), .ZN(new_n1040));
  OR4_X1    g0840(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n269), .B1(new_n792), .B2(new_n584), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G294), .B2(new_n772), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n775), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1044), .A2(G107), .B1(G311), .B2(new_n797), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G283), .A2(new_n795), .B1(new_n807), .B2(G317), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n485), .C2(new_n786), .ZN(new_n1048));
  AOI21_X1  g0848(.A(KEYINPUT114), .B1(new_n779), .B2(G116), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT46), .Z(new_n1050));
  OAI21_X1  g0850(.A(new_n1041), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT47), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1035), .B1(new_n1052), .B2(new_n767), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1030), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1029), .A2(new_n1054), .ZN(G387));
  INV_X1    g0855(.A(new_n1020), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n690), .A2(new_n755), .ZN(new_n1057));
  OR3_X1    g0857(.A1(new_n239), .A2(new_n257), .A3(new_n271), .ZN(new_n1058));
  XOR2_X1   g0858(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(G50), .B2(new_n294), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1060), .B(new_n257), .C1(new_n203), .C2(new_n210), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n1059), .A2(G50), .A3(new_n294), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n269), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n706), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n703), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n768), .B1(new_n224), .B2(new_n375), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1031), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n794), .A2(new_n203), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n778), .A2(new_n210), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(G50), .C2(new_n793), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n271), .B1(new_n783), .B2(new_n295), .C1(new_n773), .C2(new_n294), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n541), .A2(new_n775), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n797), .B2(G159), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n787), .A2(G97), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1070), .A2(new_n1072), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n271), .B1(new_n807), .B2(G326), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n778), .A2(new_n624), .B1(new_n775), .B2(new_n862), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n794), .A2(new_n584), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G317), .B2(new_n793), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n805), .B2(new_n773), .C1(new_n804), .C2(new_n798), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT48), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1078), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT49), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1077), .B1(new_n577), .B2(new_n786), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1076), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1067), .B1(new_n1088), .B2(new_n767), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1056), .A2(new_n758), .B1(new_n1057), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1021), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(KEYINPUT116), .A3(new_n704), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n750), .B2(new_n1056), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT116), .B1(new_n1091), .B2(new_n704), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1090), .B1(new_n1093), .B2(new_n1094), .ZN(G393));
  NAND3_X1  g0895(.A1(new_n1017), .A2(new_n758), .A3(new_n1022), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1032), .A2(new_n246), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n768), .B1(new_n224), .B2(new_n485), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1031), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n861), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n798), .A2(new_n295), .B1(new_n792), .B2(new_n784), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT51), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n778), .A2(new_n203), .B1(new_n783), .B2(new_n1039), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n269), .B(new_n1103), .C1(new_n390), .C2(new_n795), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n775), .A2(new_n210), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n772), .B2(G50), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n269), .B1(new_n794), .B2(new_n624), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n773), .A2(new_n584), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(G116), .C2(new_n1044), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n778), .A2(new_n862), .B1(new_n783), .B2(new_n804), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n787), .A2(G107), .B1(KEYINPUT117), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1110), .B(new_n1112), .C1(KEYINPUT117), .C2(new_n1111), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n793), .A2(G311), .B1(G317), .B2(new_n797), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT52), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1107), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1099), .B1(new_n1116), .B2(new_n767), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n755), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n991), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1096), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1023), .A2(new_n704), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1091), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1120), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(G390));
  INV_X1    g0925(.A(new_n935), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n747), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n817), .B1(new_n1127), .B2(new_n932), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1128), .A2(new_n948), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n826), .A2(new_n834), .A3(new_n679), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n656), .B2(new_n663), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n937), .B1(new_n1131), .B2(new_n918), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n904), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT39), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n942), .B2(new_n943), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1132), .A2(new_n1133), .B1(new_n1135), .B2(new_n893), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n904), .B1(new_n884), .B2(new_n898), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n679), .B(new_n836), .C1(new_n715), .C2(new_n721), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n919), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1138), .B1(new_n1140), .B2(new_n937), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1129), .B1(new_n1136), .B2(new_n1141), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n920), .A2(new_n904), .B1(new_n894), .B2(new_n899), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n720), .A2(new_n719), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n717), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n678), .B1(new_n1145), .B2(new_n656), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n918), .B1(new_n1146), .B2(new_n836), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1137), .B1(new_n1147), .B2(new_n916), .ZN(new_n1148));
  OAI211_X1 g0948(.A(G330), .B(new_n836), .C1(new_n746), .C2(new_n747), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1149), .A2(new_n916), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1143), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1142), .A2(new_n1151), .A3(new_n758), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n761), .B1(new_n294), .B2(new_n846), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n853), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n271), .B(new_n1105), .C1(G87), .C2(new_n779), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G107), .A2(new_n772), .B1(new_n797), .B2(G283), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n792), .A2(new_n577), .B1(new_n783), .B2(new_n624), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G97), .B2(new_n795), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(KEYINPUT54), .B(G143), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n794), .A2(new_n1161), .B1(new_n775), .B2(new_n784), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G137), .B2(new_n772), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT119), .Z(new_n1164));
  AOI22_X1  g0964(.A1(G132), .A2(new_n793), .B1(new_n807), .B2(G125), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1165), .B(new_n271), .C1(new_n231), .C2(new_n786), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1167));
  NAND3_X1  g0967(.A1(new_n779), .A2(G150), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1167), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n778), .B2(new_n295), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1168), .B(new_n1170), .C1(new_n798), .C2(new_n1171), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1166), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1160), .B1(new_n1164), .B2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(KEYINPUT121), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(KEYINPUT121), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n767), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1154), .B1(new_n1175), .B2(new_n1177), .C1(new_n900), .C2(new_n754), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1152), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT122), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT122), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1152), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1128), .A2(new_n480), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n925), .A2(new_n1184), .A3(new_n652), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1128), .A2(new_n948), .B1(new_n1149), .B2(new_n916), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1131), .A2(new_n918), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n937), .B1(new_n1128), .B2(new_n836), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n919), .B(new_n1139), .C1(new_n1149), .C2(new_n916), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n1187), .A2(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1142), .A2(new_n1151), .A3(new_n1186), .A4(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1192), .A2(new_n704), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1142), .A2(new_n1151), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1191), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1194), .B1(new_n1195), .B2(new_n1185), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1183), .A2(new_n1197), .ZN(G378));
  INV_X1    g0998(.A(KEYINPUT124), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1185), .B(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1192), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT57), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n945), .A2(new_n949), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n817), .B1(new_n950), .B2(new_n946), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n319), .A2(new_n675), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n330), .B2(new_n643), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n408), .B(new_n1206), .C1(new_n478), .C2(new_n325), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1210), .B(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1205), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1203), .A2(new_n1212), .A3(new_n1204), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1214), .A2(new_n924), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n924), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1217));
  OAI21_X1  g1017(.A(KEYINPUT125), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1214), .A2(new_n924), .A3(new_n1215), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT125), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1202), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n924), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1203), .A2(new_n1212), .A3(new_n1204), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1212), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1226), .A2(new_n1219), .B1(new_n1192), .B2(new_n1200), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n704), .B1(new_n1227), .B2(KEYINPUT57), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1222), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1213), .A2(new_n754), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n269), .A2(new_n256), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1231), .B(new_n1069), .C1(G68), .C2(new_n1044), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n541), .A2(new_n794), .B1(new_n786), .B2(new_n202), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n792), .A2(new_n375), .B1(new_n783), .B2(new_n862), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(G97), .A2(new_n772), .B1(new_n797), .B2(G116), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1232), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT58), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G50), .B1(new_n263), .B2(new_n256), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1237), .A2(new_n1238), .B1(new_n1231), .B2(new_n1239), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n792), .A2(new_n1171), .B1(new_n794), .B2(new_n849), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n778), .A2(new_n1161), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1242), .A2(KEYINPUT123), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G125), .B2(new_n797), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1044), .A2(G150), .B1(G132), .B2(new_n772), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1241), .B(new_n1246), .C1(KEYINPUT123), .C2(new_n1242), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(KEYINPUT59), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n263), .B(new_n256), .C1(new_n786), .C2(new_n784), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G124), .B2(new_n807), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT59), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1251), .B1(new_n1247), .B2(new_n1252), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1240), .B1(new_n1238), .B2(new_n1237), .C1(new_n1249), .C2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n767), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n761), .B1(new_n231), .B2(new_n846), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1230), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1226), .A2(new_n1219), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1259), .B2(new_n758), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1229), .A2(new_n1260), .ZN(G375));
  AOI21_X1  g1061(.A(new_n761), .B1(new_n203), .B2(new_n846), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G283), .A2(new_n793), .B1(new_n807), .B2(G303), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n485), .B2(new_n778), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(G77), .B2(new_n787), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n773), .A2(new_n577), .B1(new_n798), .B2(new_n624), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n269), .B1(new_n794), .B2(new_n375), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1266), .A2(new_n1073), .A3(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n271), .B1(new_n786), .B2(new_n202), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n855), .A2(new_n798), .B1(new_n773), .B2(new_n1161), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1269), .B(new_n1270), .C1(G50), .C2(new_n1044), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n778), .A2(new_n784), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n792), .A2(new_n849), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n794), .A2(new_n295), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n783), .A2(new_n1171), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1265), .A2(new_n1268), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n1262), .B1(new_n770), .B2(new_n1277), .C1(new_n937), .C2(new_n754), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n757), .B(KEYINPUT126), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1278), .B1(new_n1195), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1191), .A2(new_n1186), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1000), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1195), .B2(new_n1185), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1281), .B1(new_n1282), .B2(new_n1284), .ZN(G381));
  INV_X1    g1085(.A(G375), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1180), .A2(new_n1182), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1287));
  OR2_X1    g1087(.A1(G381), .A2(G384), .ZN(new_n1288));
  NOR4_X1   g1088(.A1(new_n1288), .A2(G396), .A3(G390), .A4(G393), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1290));
  OR2_X1    g1090(.A1(new_n1290), .A2(G387), .ZN(G407));
  OR3_X1    g1091(.A1(G375), .A2(G343), .A3(G378), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G407), .A2(G213), .A3(new_n1292), .ZN(G409));
  XNOR2_X1  g1093(.A(G393), .B(G396), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G387), .A2(new_n1124), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1029), .A2(new_n1054), .A3(G390), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(G390), .B1(new_n1029), .B2(new_n1054), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1054), .ZN(new_n1300));
  AOI211_X1 g1100(.A(new_n1300), .B(new_n1124), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1299), .A2(new_n1301), .A3(new_n1294), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1298), .A2(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G378), .B(new_n1260), .C1(new_n1222), .C2(new_n1228), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1279), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1259), .A2(new_n1283), .A3(new_n1201), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1258), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1287), .B1(new_n1305), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1304), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(G213), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1311), .A2(G343), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(G2897), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(KEYINPUT60), .B1(new_n1195), .B2(new_n1185), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1282), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  OR2_X1    g1119(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1320));
  OR2_X1    g1120(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(KEYINPUT60), .A4(new_n1185), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1319), .A2(new_n704), .A3(new_n1322), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1323), .A2(new_n1281), .A3(G384), .ZN(new_n1324));
  AOI21_X1  g1124(.A(G384), .B1(new_n1323), .B2(new_n1281), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1316), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1323), .A2(new_n1281), .ZN(new_n1327));
  INV_X1    g1127(.A(G384), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1323), .A2(new_n1281), .A3(G384), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(new_n1330), .A3(new_n1315), .ZN(new_n1331));
  AND2_X1   g1131(.A1(new_n1326), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT61), .B1(new_n1314), .B2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1312), .B1(new_n1304), .B2(new_n1309), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1334), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1335), .B1(new_n1334), .B2(new_n1336), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1303), .B(new_n1333), .C1(new_n1337), .C2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT62), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1334), .A2(new_n1340), .A3(new_n1336), .ZN(new_n1341));
  XNOR2_X1  g1141(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1326), .A2(new_n1331), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1342), .B1(new_n1334), .B2(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1340), .B1(new_n1334), .B2(new_n1336), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1341), .A2(new_n1344), .A3(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1339), .B1(new_n1346), .B2(new_n1303), .ZN(G405));
  NAND2_X1  g1147(.A1(G375), .A2(new_n1287), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1336), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1348), .A2(new_n1304), .A3(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1349), .B1(new_n1348), .B2(new_n1304), .ZN(new_n1352));
  OAI22_X1  g1152(.A1(new_n1351), .A2(new_n1352), .B1(new_n1302), .B2(new_n1298), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1352), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1354), .A2(new_n1303), .A3(new_n1350), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1353), .A2(new_n1355), .ZN(G402));
endmodule


