//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT65), .B(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n207), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n201), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT64), .Z(new_n227));
  OAI221_X1 g0027(.A(new_n212), .B1(KEYINPUT1), .B2(new_n221), .C1(new_n224), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT67), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT69), .ZN(new_n242));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G41), .ZN(new_n250));
  OAI211_X1 g0050(.A(G1), .B(G13), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  MUX2_X1   g0051(.A(G222), .B(G223), .S(G1698), .Z(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n254), .B1(new_n255), .B2(new_n253), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n251), .B1(new_n256), .B2(KEYINPUT71), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(KEYINPUT71), .B2(new_n256), .ZN(new_n258));
  AND2_X1   g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n222), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(new_n222), .B2(new_n259), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT70), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT70), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n251), .A2(new_n266), .A3(new_n262), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n263), .B1(new_n268), .B2(G226), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n258), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G200), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n258), .A2(G190), .A3(new_n269), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT9), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n222), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n203), .A2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT8), .ZN(new_n281));
  INV_X1    g0081(.A(G58), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(KEYINPUT72), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT72), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(KEYINPUT8), .A3(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n207), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n275), .B1(new_n280), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT73), .ZN(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n291), .A2(new_n207), .A3(G1), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G50), .ZN(new_n294));
  INV_X1    g0094(.A(new_n275), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n206), .A2(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n294), .B1(new_n298), .B2(G50), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n290), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n289), .A2(KEYINPUT73), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n273), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n300), .A2(KEYINPUT9), .A3(new_n302), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n271), .B(new_n272), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n300), .A2(new_n302), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n270), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n258), .A2(new_n313), .A3(new_n269), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n293), .A2(new_n286), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n298), .B2(new_n286), .ZN(new_n318));
  INV_X1    g0118(.A(G68), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT65), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT65), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G68), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT3), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G33), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT7), .B1(new_n327), .B2(new_n207), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT7), .ZN(new_n329));
  AOI211_X1 g0129(.A(new_n329), .B(G20), .C1(new_n324), .C2(new_n326), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n323), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G159), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n279), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n225), .B1(new_n213), .B2(new_n282), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(G20), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n295), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT80), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n324), .A2(new_n326), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n249), .A2(KEYINPUT80), .A3(KEYINPUT3), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT81), .ZN(new_n342));
  AOI21_X1  g0142(.A(G20), .B1(new_n342), .B2(new_n329), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(KEYINPUT81), .A2(KEYINPUT7), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n340), .A2(new_n341), .A3(new_n343), .A4(new_n345), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(G68), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT82), .ZN(new_n350));
  AOI211_X1 g0150(.A(new_n350), .B(new_n333), .C1(new_n334), .C2(G20), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n282), .B1(new_n320), .B2(new_n322), .ZN(new_n352));
  OAI21_X1  g0152(.A(G20), .B1(new_n352), .B2(new_n201), .ZN(new_n353));
  INV_X1    g0153(.A(new_n333), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT82), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT16), .B(new_n349), .C1(new_n351), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT83), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n338), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n357), .B1(new_n338), .B2(new_n356), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n318), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n260), .A2(new_n261), .ZN(new_n361));
  INV_X1    g0161(.A(new_n262), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n251), .A2(G232), .A3(new_n262), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(G1698), .B1(new_n340), .B2(new_n341), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G223), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n340), .A2(new_n341), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(G226), .A3(G1698), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G87), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT84), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n365), .B1(new_n372), .B2(new_n260), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT85), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n363), .A2(new_n375), .A3(new_n364), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n375), .B1(new_n363), .B2(new_n364), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n377), .A2(new_n378), .A3(G179), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n372), .A2(new_n260), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n374), .A2(new_n311), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n360), .A2(KEYINPUT18), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT18), .B1(new_n360), .B2(new_n381), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G226), .A2(G1698), .ZN(new_n385));
  INV_X1    g0185(.A(G232), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(G1698), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(new_n253), .B1(G33), .B2(G97), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n363), .B1(new_n388), .B2(new_n251), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n214), .B1(new_n265), .B2(new_n267), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n389), .A2(KEYINPUT13), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT13), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(G1698), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(G226), .B2(G1698), .ZN(new_n394));
  INV_X1    g0194(.A(G97), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n394), .A2(new_n327), .B1(new_n249), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n263), .B1(new_n396), .B2(new_n260), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n264), .A2(KEYINPUT70), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n266), .B1(new_n251), .B2(new_n262), .ZN(new_n399));
  OAI21_X1  g0199(.A(G238), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n392), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(G169), .B1(new_n391), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT14), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT13), .B1(new_n389), .B2(new_n390), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n397), .A2(new_n400), .A3(new_n392), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(G179), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT14), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(G169), .C1(new_n391), .C2(new_n401), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n292), .A2(new_n275), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT78), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n292), .B2(new_n275), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n411), .A2(G68), .A3(new_n296), .A4(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT12), .B1(new_n292), .B2(new_n319), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n323), .A2(new_n207), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n291), .A2(G1), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n417), .A2(KEYINPUT12), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n415), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n278), .A2(G50), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n420), .B1(new_n255), .B2(new_n287), .C1(new_n323), .C2(new_n207), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT11), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n421), .A2(new_n422), .A3(new_n275), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n422), .B1(new_n421), .B2(new_n275), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n414), .B(new_n419), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n404), .A2(new_n405), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G200), .ZN(new_n427));
  INV_X1    g0227(.A(new_n425), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n404), .A2(G190), .A3(new_n405), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n409), .A2(new_n425), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n411), .A2(G77), .A3(new_n296), .A4(new_n413), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT79), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n292), .A2(new_n255), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT8), .B(G58), .Z(new_n435));
  NAND2_X1  g0235(.A1(new_n279), .A2(KEYINPUT76), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT76), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n278), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT77), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G20), .A2(G77), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n440), .B1(new_n439), .B2(new_n441), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT15), .B(G87), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(new_n287), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n433), .B(new_n434), .C1(new_n446), .C2(new_n295), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n327), .A2(G107), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G238), .A2(G1698), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n386), .B2(G1698), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n253), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n251), .B1(new_n452), .B2(KEYINPUT74), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(KEYINPUT74), .B2(new_n452), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n263), .B1(new_n268), .B2(G244), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n454), .A2(KEYINPUT75), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT75), .B1(new_n454), .B2(new_n455), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n447), .B1(G200), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(G190), .B1(new_n456), .B2(new_n457), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n311), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n313), .B1(new_n456), .B2(new_n457), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n447), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n431), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n380), .ZN(new_n466));
  INV_X1    g0266(.A(new_n378), .ZN(new_n467));
  INV_X1    g0267(.A(G190), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(new_n376), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n466), .A2(new_n469), .B1(new_n373), .B2(G200), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(new_n318), .C1(new_n358), .C2(new_n359), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT17), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NOR4_X1   g0273(.A1(new_n316), .A2(new_n384), .A3(new_n465), .A4(new_n473), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(G257), .A3(new_n251), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n475), .A2(new_n251), .A3(G274), .A4(new_n477), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G250), .A2(G1698), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT4), .A2(G244), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(G1698), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n253), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G1698), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n368), .A2(G244), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n482), .B1(new_n492), .B2(new_n251), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT6), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n494), .A2(new_n395), .A3(G107), .ZN(new_n495));
  XNOR2_X1  g0295(.A(G97), .B(G107), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n497), .A2(new_n207), .B1(new_n255), .B2(new_n279), .ZN(new_n498));
  INV_X1    g0298(.A(G107), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n329), .B1(new_n253), .B2(G20), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n327), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n275), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n293), .A2(G97), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n206), .A2(G33), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n410), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n505), .B1(new_n507), .B2(new_n395), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n493), .A2(new_n311), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT86), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n492), .B2(new_n251), .ZN(new_n512));
  INV_X1    g0312(.A(G244), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n340), .B2(new_n341), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT4), .B1(new_n514), .B2(new_n489), .ZN(new_n515));
  OAI211_X1 g0315(.A(KEYINPUT86), .B(new_n260), .C1(new_n515), .C2(new_n488), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT87), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n481), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n479), .A2(KEYINPUT87), .A3(new_n480), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n512), .A2(new_n313), .A3(new_n516), .A4(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n510), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n477), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n523), .A2(G250), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n251), .ZN(new_n525));
  INV_X1    g0325(.A(new_n361), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(new_n523), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n514), .A2(G1698), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n368), .A2(G238), .A3(new_n489), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G116), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n527), .B1(new_n531), .B2(new_n260), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n313), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n366), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n251), .B1(new_n534), .B2(new_n528), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n311), .B1(new_n535), .B2(new_n527), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n340), .A2(new_n341), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n207), .A2(G68), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n207), .B1(new_n249), .B2(new_n395), .ZN(new_n540));
  INV_X1    g0340(.A(G87), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(new_n395), .A3(new_n499), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n539), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n287), .A2(KEYINPUT19), .A3(new_n395), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n537), .A2(new_n538), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n275), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n444), .A2(new_n292), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n546), .B(new_n547), .C1(new_n444), .C2(new_n507), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n533), .A2(new_n536), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(G200), .B1(new_n535), .B2(new_n527), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n531), .A2(new_n260), .ZN(new_n551));
  INV_X1    g0351(.A(new_n527), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(G190), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n410), .A2(G87), .A3(new_n506), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n546), .A2(new_n547), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n550), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(G200), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n260), .B1(new_n515), .B2(new_n488), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(new_n511), .B1(new_n518), .B2(new_n519), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n558), .B1(new_n560), .B2(new_n516), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n496), .A2(new_n494), .ZN(new_n562));
  INV_X1    g0362(.A(new_n495), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(G20), .B1(G77), .B2(new_n278), .ZN(new_n565));
  OAI21_X1  g0365(.A(G107), .B1(new_n328), .B2(new_n330), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n508), .B1(new_n567), .B2(new_n275), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n559), .A2(G190), .A3(new_n482), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT88), .B1(new_n561), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n512), .A2(new_n516), .A3(new_n520), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G200), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n568), .A2(new_n569), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT88), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n522), .B(new_n557), .C1(new_n571), .C2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n368), .A2(G264), .A3(G1698), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT89), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT89), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n368), .A2(new_n580), .A3(G264), .A4(G1698), .ZN(new_n581));
  INV_X1    g0381(.A(G303), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n253), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(G257), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n340), .B2(new_n341), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n583), .B1(new_n585), .B2(new_n489), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n579), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n260), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n260), .B1(new_n477), .B2(new_n475), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G270), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n480), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n411), .A2(G116), .A3(new_n413), .A4(new_n506), .ZN(new_n593));
  INV_X1    g0393(.A(G116), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n417), .A2(G20), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n487), .B(new_n207), .C1(G33), .C2(new_n395), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n596), .B(new_n275), .C1(new_n207), .C2(G116), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT20), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n593), .B(new_n595), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n588), .A2(G179), .A3(new_n592), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT90), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n591), .B1(new_n587), .B2(new_n260), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT90), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(G179), .A4(new_n601), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n601), .A2(G169), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(G190), .ZN(new_n611));
  INV_X1    g0411(.A(new_n601), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n611), .B(new_n612), .C1(new_n558), .C2(new_n604), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n588), .A2(new_n592), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n614), .A2(KEYINPUT21), .A3(G169), .A4(new_n601), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n607), .A2(new_n610), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n585), .A2(G1698), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n368), .A2(G250), .A3(new_n489), .ZN(new_n618));
  NAND2_X1  g0418(.A1(G33), .A2(G294), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n620), .A2(new_n260), .B1(G264), .B2(new_n589), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(G179), .A3(new_n480), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n260), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n589), .A2(G264), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n623), .A2(new_n480), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n622), .B1(new_n625), .B2(new_n311), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT22), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n207), .A2(G87), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n627), .B1(new_n327), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT23), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n630), .A2(new_n499), .A3(KEYINPUT92), .A4(G20), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n499), .A3(G20), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT92), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n499), .A2(G20), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n632), .A2(new_n633), .B1(new_n634), .B2(KEYINPUT23), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT91), .B1(new_n530), .B2(G20), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT91), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n637), .A2(new_n207), .A3(G33), .A4(G116), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n629), .A2(new_n631), .A3(new_n635), .A4(new_n639), .ZN(new_n640));
  AOI211_X1 g0440(.A(new_n627), .B(new_n628), .C1(new_n340), .C2(new_n341), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT24), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n628), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n368), .A2(KEYINPUT22), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n253), .A2(new_n643), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n645), .A2(new_n627), .B1(new_n636), .B2(new_n638), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n635), .A2(new_n631), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT24), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n644), .A2(new_n646), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n295), .B1(new_n642), .B2(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n292), .A2(KEYINPUT25), .A3(new_n499), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT25), .B1(new_n292), .B2(new_n499), .ZN(new_n652));
  OAI22_X1  g0452(.A1(new_n507), .A2(new_n499), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n626), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n621), .A2(new_n480), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G200), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n621), .A2(G190), .A3(new_n480), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n654), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n616), .A2(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n474), .A2(new_n577), .A3(new_n662), .ZN(G372));
  INV_X1    g0463(.A(new_n315), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT93), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n382), .B2(new_n383), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT18), .ZN(new_n667));
  INV_X1    g0467(.A(new_n318), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n338), .A2(new_n356), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT83), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n338), .A2(new_n356), .A3(new_n357), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n381), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n667), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n360), .A2(KEYINPUT18), .A3(new_n381), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(KEYINPUT93), .A3(new_n675), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n666), .A2(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n462), .A2(new_n447), .A3(new_n463), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n430), .A2(new_n427), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n678), .A2(new_n679), .B1(new_n425), .B2(new_n409), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n677), .B1(new_n473), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n664), .B1(new_n681), .B2(new_n309), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n615), .A2(new_n610), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(new_n607), .A3(new_n656), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n522), .B1(new_n571), .B2(new_n576), .ZN(new_n685));
  INV_X1    g0485(.A(new_n557), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .A4(new_n660), .ZN(new_n687));
  INV_X1    g0487(.A(new_n549), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(KEYINPUT26), .A3(new_n522), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n510), .A2(new_n521), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n557), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n688), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n474), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n682), .A2(new_n695), .ZN(G369));
  INV_X1    g0496(.A(new_n417), .ZN(new_n697));
  OR3_X1    g0497(.A1(new_n697), .A2(KEYINPUT27), .A3(G20), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT27), .B1(new_n697), .B2(G20), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G343), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n655), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n656), .A2(new_n660), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n657), .A2(G169), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n654), .B1(new_n705), .B2(new_n622), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT95), .B1(new_n706), .B2(new_n702), .ZN(new_n707));
  AND4_X1   g0507(.A1(KEYINPUT95), .A2(new_n626), .A3(new_n655), .A4(new_n702), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT94), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n683), .A2(new_n607), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n601), .A2(new_n702), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n683), .A2(new_n607), .A3(new_n613), .A4(new_n712), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n710), .B1(new_n716), .B2(G330), .ZN(new_n717));
  INV_X1    g0517(.A(G330), .ZN(new_n718));
  AOI211_X1 g0518(.A(KEYINPUT94), .B(new_n718), .C1(new_n714), .C2(new_n715), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n709), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n656), .A2(new_n702), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n702), .B1(new_n683), .B2(new_n607), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n709), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(new_n723), .ZN(G399));
  INV_X1    g0524(.A(new_n210), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G41), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n542), .A2(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n226), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n702), .B1(new_n687), .B2(new_n693), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT29), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(KEYINPUT96), .B(KEYINPUT31), .Z(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n572), .A2(new_n657), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n551), .A2(new_n552), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n614), .A2(KEYINPUT97), .A3(new_n313), .A4(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT97), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n313), .B1(new_n535), .B2(new_n527), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n743), .B1(new_n744), .B2(new_n604), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n740), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n604), .A2(G179), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n621), .A2(new_n532), .A3(new_n559), .A4(new_n482), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n741), .A2(new_n493), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n313), .B(new_n591), .C1(new_n587), .C2(new_n260), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n751), .A2(new_n752), .A3(KEYINPUT30), .A4(new_n621), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n702), .B(new_n739), .C1(new_n746), .C2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n702), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n750), .A2(new_n753), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n740), .A2(new_n742), .A3(new_n745), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n755), .B1(new_n759), .B2(KEYINPUT31), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n561), .A2(KEYINPUT88), .A3(new_n570), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n575), .B1(new_n573), .B2(new_n574), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n686), .B(new_n691), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NOR4_X1   g0563(.A1(new_n763), .A2(new_n616), .A3(new_n661), .A4(new_n702), .ZN(new_n764));
  OAI21_X1  g0564(.A(G330), .B1(new_n760), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n737), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n731), .B1(new_n767), .B2(G1), .ZN(G364));
  NAND2_X1  g0568(.A1(new_n716), .A2(G330), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(KEYINPUT94), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n716), .A2(new_n710), .A3(G330), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n291), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n206), .B1(new_n774), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n726), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n773), .B(new_n778), .C1(G330), .C2(new_n716), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n468), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n207), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n395), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n207), .A2(new_n313), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n558), .A2(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n782), .B1(new_n789), .B2(G68), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT101), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n207), .A2(G179), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n784), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G107), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G190), .A2(G200), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(KEYINPUT32), .B1(new_n797), .B2(new_n332), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n795), .A2(new_n253), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n468), .A2(new_n558), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n783), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n783), .A2(new_n796), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n801), .A2(new_n202), .B1(new_n802), .B2(new_n255), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n783), .A2(G190), .A3(new_n558), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n800), .A2(new_n792), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n804), .A2(new_n282), .B1(new_n805), .B2(new_n541), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n797), .A2(KEYINPUT32), .A3(new_n332), .ZN(new_n807));
  NOR4_X1   g0607(.A1(new_n799), .A2(new_n803), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n327), .B1(new_n805), .B2(new_n582), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT102), .ZN(new_n810));
  INV_X1    g0610(.A(new_n804), .ZN(new_n811));
  INV_X1    g0611(.A(new_n797), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n811), .A2(G322), .B1(new_n812), .B2(G329), .ZN(new_n813));
  INV_X1    g0613(.A(G294), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n814), .B2(new_n781), .ZN(new_n815));
  INV_X1    g0615(.A(new_n801), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G326), .A2(new_n816), .B1(new_n794), .B2(G283), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n818), .B2(new_n802), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT33), .B(G317), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n815), .B(new_n819), .C1(new_n789), .C2(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n791), .A2(new_n808), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n222), .B1(G20), .B2(new_n311), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n777), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n725), .A2(new_n327), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n826), .A2(G355), .B1(new_n594), .B2(new_n725), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n244), .A2(G45), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT98), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n725), .A2(new_n368), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n227), .B2(G45), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n827), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(G13), .A2(G33), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(G20), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n823), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT99), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n825), .B1(new_n832), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n835), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n716), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n779), .A2(new_n841), .ZN(G396));
  NAND4_X1  g0642(.A1(new_n462), .A2(new_n447), .A3(new_n463), .A4(new_n756), .ZN(new_n843));
  INV_X1    g0643(.A(new_n446), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n844), .A2(new_n275), .B1(new_n255), .B2(new_n292), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n756), .B1(new_n845), .B2(new_n433), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n459), .B2(new_n460), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n843), .B1(new_n847), .B2(new_n678), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n732), .B(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(new_n765), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT105), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n777), .B1(new_n850), .B2(new_n765), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n789), .A2(G283), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n327), .B1(new_n805), .B2(new_n499), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT103), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n804), .A2(new_n814), .B1(new_n801), .B2(new_n582), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G311), .B2(new_n812), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n802), .A2(new_n594), .B1(new_n793), .B2(new_n541), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(new_n782), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n855), .A2(new_n857), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n794), .A2(G68), .ZN(new_n863));
  INV_X1    g0663(.A(G132), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n863), .B1(new_n202), .B2(new_n805), .C1(new_n864), .C2(new_n797), .ZN(new_n865));
  INV_X1    g0665(.A(new_n781), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n537), .B(new_n865), .C1(G58), .C2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n802), .ZN(new_n868));
  AOI22_X1  g0668(.A1(G137), .A2(new_n816), .B1(new_n868), .B2(G159), .ZN(new_n869));
  INV_X1    g0669(.A(G143), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n869), .B1(new_n870), .B2(new_n804), .C1(new_n788), .C2(new_n277), .ZN(new_n871));
  XOR2_X1   g0671(.A(KEYINPUT104), .B(KEYINPUT34), .Z(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n867), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n871), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(new_n872), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n862), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n823), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n823), .A2(new_n833), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n778), .B1(new_n255), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n848), .B2(new_n833), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n854), .A2(new_n882), .ZN(G384));
  NOR2_X1   g0683(.A1(new_n774), .A2(new_n206), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n662), .A2(new_n577), .A3(new_n756), .ZN(new_n885));
  OAI211_X1 g0685(.A(KEYINPUT31), .B(new_n702), .C1(new_n746), .C2(new_n754), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n702), .B1(new_n746), .B2(new_n754), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n738), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n408), .A2(new_n406), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n407), .B1(new_n426), .B2(G169), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n425), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n425), .A2(new_n702), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n679), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT106), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n892), .A2(new_n679), .A3(KEYINPUT106), .A4(new_n893), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n430), .A2(new_n427), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n425), .B(new_n702), .C1(new_n899), .C2(new_n409), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n848), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n889), .A2(new_n901), .A3(KEYINPUT40), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT108), .B(KEYINPUT38), .Z(new_n903));
  XNOR2_X1  g0703(.A(new_n471), .B(KEYINPUT17), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n666), .A2(new_n904), .A3(new_n676), .ZN(new_n905));
  INV_X1    g0705(.A(new_n700), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n360), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n360), .A2(KEYINPUT93), .A3(new_n381), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n471), .A3(new_n907), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT93), .B1(new_n360), .B2(new_n381), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT37), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT109), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n471), .B1(new_n672), .B2(new_n700), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT37), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n672), .B2(new_n673), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT37), .B1(new_n360), .B2(new_n381), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n919), .A2(KEYINPUT109), .A3(new_n471), .A4(new_n907), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n913), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n903), .B1(new_n909), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n915), .A2(new_n917), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n356), .A2(new_n275), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n353), .A2(new_n354), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n350), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n335), .A2(KEYINPUT82), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT16), .B1(new_n928), .B2(new_n349), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n318), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n381), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n471), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT107), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n471), .A3(KEYINPUT107), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n930), .A2(new_n906), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n923), .B1(new_n937), .B2(KEYINPUT37), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT38), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n674), .A2(new_n675), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n936), .B1(new_n904), .B2(new_n940), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n902), .B1(new_n922), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT110), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT110), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n902), .B(new_n945), .C1(new_n922), .C2(new_n942), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT40), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n889), .A2(new_n901), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n935), .A2(new_n936), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT107), .B1(new_n931), .B2(new_n471), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT37), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n923), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n941), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT38), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n948), .B1(new_n942), .B2(new_n955), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n944), .A2(new_n946), .B1(new_n947), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n474), .A2(new_n889), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n718), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT39), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n922), .B2(new_n942), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n409), .A2(new_n425), .A3(new_n756), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n939), .B1(new_n938), .B2(new_n941), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT38), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT39), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n962), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n677), .A2(new_n906), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n732), .A2(new_n849), .B1(new_n678), .B2(new_n756), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT106), .B1(new_n431), .B2(new_n893), .ZN(new_n971));
  INV_X1    g0771(.A(new_n897), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n900), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n965), .A2(new_n966), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n969), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n968), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n474), .B1(new_n734), .B2(new_n736), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n682), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n978), .B(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n884), .B1(new_n960), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n981), .B2(new_n960), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n594), .B(new_n224), .C1(new_n564), .C2(KEYINPUT35), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(KEYINPUT35), .B2(new_n564), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT36), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n352), .A2(new_n226), .A3(new_n255), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n319), .A2(G50), .ZN(new_n988));
  OAI211_X1 g0788(.A(G1), .B(new_n291), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n983), .A2(new_n986), .A3(new_n989), .ZN(G367));
  OR2_X1    g0790(.A1(new_n555), .A2(new_n756), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n686), .A2(KEYINPUT111), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n549), .B2(new_n991), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT111), .B1(new_n686), .B2(new_n991), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n835), .ZN(new_n996));
  INV_X1    g0796(.A(new_n830), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n838), .B1(new_n210), .B2(new_n444), .C1(new_n239), .C2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n778), .B1(new_n998), .B2(KEYINPUT115), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(KEYINPUT115), .B2(new_n998), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n805), .A2(new_n594), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n1001), .A2(KEYINPUT46), .B1(new_n499), .B2(new_n781), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT46), .B2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n789), .A2(G294), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(KEYINPUT116), .B(G311), .ZN(new_n1005));
  INV_X1    g0805(.A(G283), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n801), .A2(new_n1005), .B1(new_n802), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n793), .A2(new_n395), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(G317), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n804), .A2(new_n582), .B1(new_n797), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1011), .A2(new_n368), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1003), .A2(new_n1004), .A3(new_n1009), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n789), .A2(G159), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n805), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G58), .A2(new_n1015), .B1(new_n812), .B2(G137), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n794), .A2(G77), .ZN(new_n1017));
  AND3_X1   g0817(.A1(new_n1016), .A2(new_n253), .A3(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n781), .A2(new_n319), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n804), .A2(new_n277), .B1(new_n801), .B2(new_n870), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G50), .B2(new_n868), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1014), .A2(new_n1018), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1013), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT47), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1000), .B1(new_n823), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n996), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n726), .B(KEYINPUT41), .Z(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n709), .A2(new_n722), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT95), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n656), .B2(new_n756), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n706), .A2(KEYINPUT95), .A3(new_n702), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n654), .A2(new_n659), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1035), .A2(new_n658), .B1(new_n626), .B2(new_n655), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1033), .A2(new_n1034), .B1(new_n1036), .B2(new_n703), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n722), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n772), .A2(new_n1031), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1031), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n770), .A2(new_n771), .A3(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n737), .A2(new_n1040), .A3(new_n765), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT114), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT44), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n691), .B1(new_n568), .B2(new_n756), .C1(new_n761), .C2(new_n762), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n522), .A2(new_n702), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1045), .B1(new_n723), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n721), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1048), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(KEYINPUT44), .A3(new_n1052), .ZN(new_n1053));
  AND3_X1   g0853(.A1(new_n1049), .A2(new_n1053), .A3(KEYINPUT113), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT113), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1055), .B(new_n1045), .C1(new_n723), .C2(new_n1048), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n723), .A2(KEYINPUT45), .A3(new_n1048), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT45), .B1(new_n723), .B2(new_n1048), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1044), .B(new_n720), .C1(new_n1054), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT45), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n723), .A2(KEYINPUT45), .A3(new_n1048), .ZN(new_n1063));
  AOI21_X1  g0863(.A(KEYINPUT44), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1062), .A2(new_n1063), .B1(new_n1064), .B2(new_n1055), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n720), .A2(new_n1044), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n772), .A2(KEYINPUT114), .A3(new_n709), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1049), .A2(new_n1053), .A3(KEYINPUT113), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1043), .B1(new_n1060), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1030), .B1(new_n1070), .B2(new_n766), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n775), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1048), .A2(new_n709), .A3(new_n722), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1073), .A2(KEYINPUT42), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n691), .B1(new_n1046), .B2(new_n656), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n756), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1073), .A2(KEYINPUT42), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT43), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n995), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(KEYINPUT43), .B1(new_n993), .B2(new_n994), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1077), .A2(new_n1076), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1083), .A2(new_n1079), .A3(new_n995), .A4(new_n1074), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n772), .A2(new_n709), .A3(new_n1048), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1086), .A2(KEYINPUT112), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(KEYINPUT112), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1085), .A2(KEYINPUT112), .A3(new_n1086), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1028), .B1(new_n1072), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(G387));
  NAND2_X1  g0894(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n766), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n726), .A3(new_n1043), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n435), .A2(new_n202), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT50), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n728), .B(new_n476), .C1(new_n319), .C2(new_n255), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n830), .B1(new_n1099), .B2(new_n1100), .C1(new_n235), .C2(new_n476), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n826), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1101), .B1(G107), .B2(new_n210), .C1(new_n728), .C2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n778), .B1(new_n1103), .B2(new_n838), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n804), .A2(new_n1010), .B1(new_n802), .B2(new_n582), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n816), .A2(G322), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(new_n788), .C2(new_n1005), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT48), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n866), .A2(G283), .B1(new_n1015), .B2(G294), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT118), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT49), .ZN(new_n1115));
  OR2_X1    g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n793), .A2(new_n594), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n368), .B(new_n1118), .C1(G326), .C2(new_n812), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1116), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n286), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n789), .A2(new_n1121), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n781), .A2(new_n444), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n805), .A2(new_n255), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n537), .A2(new_n1124), .A3(new_n1008), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n801), .A2(new_n332), .B1(new_n802), .B2(new_n319), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n804), .A2(new_n202), .B1(new_n797), .B2(new_n277), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .A4(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1120), .A2(new_n1129), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1104), .B1(new_n709), .B2(new_n840), .C1(new_n1130), .C2(new_n824), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1040), .A2(new_n1042), .A3(new_n776), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1097), .A2(new_n1133), .ZN(G393));
  AOI21_X1  g0934(.A(new_n837), .B1(G97), .B2(new_n725), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n830), .A2(new_n247), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n778), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n795), .B(new_n327), .C1(new_n594), .C2(new_n781), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G294), .A2(new_n868), .B1(new_n812), .B2(G322), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n1006), .B2(new_n805), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1138), .B(new_n1140), .C1(G303), .C2(new_n789), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n804), .A2(new_n818), .B1(new_n801), .B2(new_n1010), .ZN(new_n1142));
  XOR2_X1   g0942(.A(KEYINPUT119), .B(KEYINPUT52), .Z(new_n1143));
  XNOR2_X1  g0943(.A(new_n1142), .B(new_n1143), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n804), .A2(new_n332), .B1(new_n801), .B2(new_n277), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT51), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n788), .A2(new_n202), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n866), .A2(G77), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n368), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n793), .A2(new_n541), .B1(new_n797), .B2(new_n870), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n435), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1151), .A2(new_n802), .B1(new_n213), .B2(new_n805), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1147), .A2(new_n1149), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1141), .A2(new_n1144), .B1(new_n1146), .B2(new_n1153), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1137), .B1(new_n824), .B2(new_n1154), .C1(new_n1048), .C2(new_n840), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1060), .A2(new_n1069), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n776), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1043), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1060), .A2(new_n1069), .A3(new_n1043), .ZN(new_n1161));
  AND4_X1   g0961(.A1(KEYINPUT120), .A2(new_n1160), .A3(new_n726), .A4(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n727), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT120), .B1(new_n1163), .B2(new_n1161), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1158), .B1(new_n1162), .B2(new_n1164), .ZN(G390));
  NAND3_X1  g0965(.A1(new_n694), .A2(new_n756), .A3(new_n849), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n843), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT121), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n886), .B1(new_n759), .B2(new_n739), .ZN(new_n1169));
  OAI21_X1  g0969(.A(G330), .B1(new_n1169), .B2(new_n764), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n973), .A2(new_n849), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1168), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n889), .A2(new_n901), .A3(KEYINPUT121), .A4(G330), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g0974(.A(G330), .B(new_n849), .C1(new_n760), .C2(new_n764), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1175), .A2(new_n974), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1167), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1175), .A2(new_n974), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n974), .B1(new_n1170), .B2(new_n848), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n970), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n474), .A2(G330), .A3(new_n889), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n979), .A2(new_n1183), .A3(new_n682), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1174), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n962), .A2(new_n967), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n963), .B1(new_n970), .B2(new_n974), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n964), .B1(new_n1167), .B2(new_n973), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n918), .A2(new_n920), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1192), .A2(new_n913), .B1(new_n905), .B2(new_n908), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n966), .B1(new_n1193), .B2(new_n903), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1187), .B1(new_n1190), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1191), .B1(new_n962), .B2(new_n967), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n922), .A2(new_n942), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(new_n1189), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1197), .A2(new_n1199), .A3(new_n1178), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1186), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1190), .A2(new_n1195), .A3(new_n1179), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1174), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1202), .A2(new_n1203), .A3(new_n1185), .A4(new_n1182), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1201), .A2(new_n726), .A3(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n776), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1188), .A2(new_n833), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n879), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n777), .B1(new_n1121), .B2(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n805), .A2(new_n277), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT53), .ZN(new_n1211));
  INV_X1    g1011(.A(G137), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n788), .ZN(new_n1213));
  INV_X1    g1013(.A(G128), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n253), .B1(new_n801), .B2(new_n1214), .C1(new_n781), .C2(new_n332), .ZN(new_n1215));
  INV_X1    g1015(.A(G125), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n793), .A2(new_n202), .B1(new_n797), .B2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(KEYINPUT54), .B(G143), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n804), .A2(new_n864), .B1(new_n802), .B2(new_n1218), .ZN(new_n1219));
  OR3_X1    g1019(.A1(new_n1215), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G283), .A2(new_n816), .B1(new_n868), .B2(G97), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n594), .B2(new_n804), .C1(new_n788), .C2(new_n499), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n253), .B1(new_n1015), .B2(G87), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n812), .A2(G294), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1223), .A2(new_n1148), .A3(new_n863), .A4(new_n1224), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n1213), .A2(new_n1220), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1209), .B1(new_n1226), .B2(new_n823), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1207), .A2(new_n1227), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1206), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1205), .A2(new_n1229), .ZN(G378));
  AOI21_X1  g1030(.A(new_n718), .B1(new_n956), .B2(new_n947), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n310), .A2(new_n700), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n664), .B1(new_n307), .B2(new_n308), .ZN(new_n1233));
  XOR2_X1   g1033(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1232), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n316), .A2(new_n1234), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1240), .B(new_n1236), .C1(new_n310), .C2(new_n700), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(KEYINPUT124), .B(KEYINPUT55), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1239), .A2(new_n1241), .A3(new_n1243), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n946), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n945), .B1(new_n1194), .B2(new_n902), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1231), .B(new_n1247), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n944), .A2(new_n946), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1247), .B1(new_n1252), .B2(new_n1231), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n978), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1231), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1247), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n978), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n1250), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n775), .B1(new_n1254), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1256), .A2(new_n833), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n777), .B1(G50), .B2(new_n1208), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT122), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n368), .A2(G41), .ZN(new_n1264));
  AOI211_X1 g1064(.A(G50), .B(new_n1264), .C1(new_n249), .C2(new_n250), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1124), .B(new_n1019), .C1(G107), .C2(new_n811), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n789), .A2(G97), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n801), .A2(new_n594), .B1(new_n793), .B2(new_n282), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n802), .A2(new_n444), .B1(new_n797), .B2(new_n1006), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1266), .A2(new_n1267), .A3(new_n1270), .A4(new_n1264), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT58), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1265), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n1212), .A2(new_n802), .B1(new_n805), .B2(new_n1218), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n804), .A2(new_n1214), .B1(new_n801), .B2(new_n1216), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n1274), .B(new_n1275), .C1(G150), .C2(new_n866), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n864), .B2(new_n788), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT59), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n249), .B(new_n250), .C1(new_n793), .C2(new_n332), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(G124), .B2(new_n812), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1277), .A2(KEYINPUT59), .ZN(new_n1282));
  OAI221_X1 g1082(.A(new_n1273), .B1(new_n1272), .B2(new_n1271), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1263), .B1(new_n1283), .B2(new_n823), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1261), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1260), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1204), .A2(new_n1185), .ZN(new_n1288));
  NOR3_X1   g1088(.A1(new_n1251), .A2(new_n1253), .A3(new_n978), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1258), .B1(new_n1257), .B2(new_n1250), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1288), .B(KEYINPUT57), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n726), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1254), .A2(new_n1259), .B1(new_n1185), .B2(new_n1204), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1293), .A2(KEYINPUT57), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1287), .B1(new_n1292), .B2(new_n1294), .ZN(G375));
  INV_X1    g1095(.A(new_n1182), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1184), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(new_n1030), .A3(new_n1186), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n778), .B1(new_n319), .B2(new_n879), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n816), .A2(G294), .B1(new_n812), .B2(G303), .ZN(new_n1300));
  AND4_X1   g1100(.A1(new_n327), .A2(new_n1300), .A3(new_n1017), .A4(new_n1123), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n811), .A2(G283), .B1(new_n868), .B2(G107), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n395), .B2(new_n805), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1303), .B1(G116), .B2(new_n789), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n788), .A2(new_n1218), .ZN(new_n1305));
  OAI22_X1  g1105(.A1(new_n804), .A2(new_n1212), .B1(new_n805), .B2(new_n332), .ZN(new_n1306));
  OAI22_X1  g1106(.A1(new_n801), .A2(new_n864), .B1(new_n802), .B2(new_n277), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1305), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n793), .A2(new_n282), .B1(new_n797), .B2(new_n1214), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n537), .B(new_n1309), .C1(G50), .C2(new_n866), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1301), .A2(new_n1304), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  OAI221_X1 g1111(.A(new_n1299), .B1(new_n824), .B2(new_n1311), .C1(new_n973), .C2(new_n834), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1296), .B2(new_n775), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1298), .A2(new_n1314), .ZN(G381));
  INV_X1    g1115(.A(G396), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1097), .A2(new_n1133), .A3(new_n1316), .ZN(new_n1317));
  OR4_X1    g1117(.A1(G384), .A2(G387), .A3(G381), .A4(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n776), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1285), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n727), .B1(new_n1293), .B2(KEYINPUT57), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1288), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT57), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1320), .B1(new_n1321), .B2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(G378), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  OR3_X1    g1127(.A1(new_n1318), .A2(new_n1327), .A3(G390), .ZN(G407));
  OAI211_X1 g1128(.A(G407), .B(G213), .C1(G343), .C2(new_n1327), .ZN(G409));
  INV_X1    g1129(.A(G213), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1330), .A2(G343), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(G2897), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1186), .A2(KEYINPUT60), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1297), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1177), .A2(new_n1184), .A3(KEYINPUT60), .A4(new_n1181), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n726), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1335), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(G384), .B1(new_n1339), .B2(new_n1314), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1337), .B1(new_n1334), .B2(new_n1297), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n854), .A2(new_n882), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1313), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1333), .B1(new_n1340), .B2(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1339), .A2(G384), .A3(new_n1314), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1342), .B1(new_n1341), .B2(new_n1313), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1345), .A2(new_n1346), .A3(new_n1332), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1344), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(G375), .A2(G378), .ZN(new_n1349));
  NOR3_X1   g1149(.A1(G378), .A2(new_n1260), .A3(new_n1286), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1293), .A2(new_n1030), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1331), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1348), .B1(new_n1349), .B2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT126), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1160), .A2(new_n726), .A3(new_n1161), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT120), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1163), .A2(KEYINPUT120), .A3(new_n1161), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1360), .B1(new_n775), .B2(new_n1071), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n1359), .B(new_n1158), .C1(new_n1361), .C2(new_n1028), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1316), .B1(new_n1097), .B2(new_n1133), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1364), .A2(KEYINPUT125), .A3(new_n1317), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT125), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1317), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1366), .B1(new_n1367), .B2(new_n1363), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1365), .A2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(G390), .A2(new_n1093), .ZN(new_n1370));
  AND4_X1   g1170(.A1(new_n1354), .A2(new_n1362), .A3(new_n1369), .A4(new_n1370), .ZN(new_n1371));
  OAI21_X1  g1171(.A(KEYINPUT126), .B1(G390), .B2(new_n1093), .ZN(new_n1372));
  AOI22_X1  g1172(.A1(new_n1372), .A2(new_n1369), .B1(new_n1362), .B2(new_n1370), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1371), .A2(new_n1373), .ZN(new_n1374));
  NOR3_X1   g1174(.A1(new_n1353), .A2(new_n1374), .A3(KEYINPUT61), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1340), .A2(new_n1343), .ZN(new_n1376));
  OAI211_X1 g1176(.A(new_n1352), .B(new_n1376), .C1(new_n1326), .C2(new_n1325), .ZN(new_n1377));
  INV_X1    g1177(.A(KEYINPUT63), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  OAI21_X1  g1179(.A(KEYINPUT127), .B1(new_n1377), .B2(new_n1378), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1287), .A2(new_n1326), .A3(new_n1351), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1331), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1381), .A2(new_n1382), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1383), .B1(G378), .B2(G375), .ZN(new_n1384));
  INV_X1    g1184(.A(KEYINPUT127), .ZN(new_n1385));
  NAND4_X1  g1185(.A1(new_n1384), .A2(new_n1385), .A3(KEYINPUT63), .A4(new_n1376), .ZN(new_n1386));
  NAND4_X1  g1186(.A1(new_n1375), .A2(new_n1379), .A3(new_n1380), .A4(new_n1386), .ZN(new_n1387));
  OAI211_X1 g1187(.A(new_n1382), .B(new_n1381), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1388));
  INV_X1    g1188(.A(new_n1348), .ZN(new_n1389));
  AOI21_X1  g1189(.A(KEYINPUT61), .B1(new_n1388), .B2(new_n1389), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1377), .A2(KEYINPUT62), .ZN(new_n1391));
  INV_X1    g1191(.A(KEYINPUT62), .ZN(new_n1392));
  NAND4_X1  g1192(.A1(new_n1349), .A2(new_n1392), .A3(new_n1352), .A4(new_n1376), .ZN(new_n1393));
  NAND3_X1  g1193(.A1(new_n1390), .A2(new_n1391), .A3(new_n1393), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1394), .A2(new_n1374), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1387), .A2(new_n1395), .ZN(G405));
  NAND2_X1  g1196(.A1(new_n1327), .A2(new_n1349), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1397), .A2(new_n1374), .ZN(new_n1398));
  INV_X1    g1198(.A(new_n1398), .ZN(new_n1399));
  NOR2_X1   g1199(.A1(new_n1397), .A2(new_n1374), .ZN(new_n1400));
  OAI22_X1  g1200(.A1(new_n1399), .A2(new_n1400), .B1(new_n1340), .B2(new_n1343), .ZN(new_n1401));
  INV_X1    g1201(.A(new_n1400), .ZN(new_n1402));
  NAND3_X1  g1202(.A1(new_n1402), .A2(new_n1376), .A3(new_n1398), .ZN(new_n1403));
  NAND2_X1  g1203(.A1(new_n1401), .A2(new_n1403), .ZN(G402));
endmodule


