

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584;

  AND2_X1 U324 ( .A1(n515), .A2(n292), .ZN(n516) );
  NOR2_X1 U325 ( .A1(n570), .A2(n574), .ZN(n292) );
  NOR2_X1 U326 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U327 ( .A(n366), .B(n293), .ZN(n335) );
  INV_X1 U328 ( .A(KEYINPUT47), .ZN(n509) );
  XOR2_X1 U329 ( .A(KEYINPUT101), .B(n441), .Z(n552) );
  XNOR2_X1 U330 ( .A(n347), .B(n346), .ZN(n507) );
  AND2_X1 U331 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  INV_X1 U332 ( .A(KEYINPUT73), .ZN(n295) );
  XNOR2_X1 U333 ( .A(G99GAT), .B(KEYINPUT74), .ZN(n294) );
  XNOR2_X1 U334 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U335 ( .A(n335), .B(n427), .ZN(n339) );
  XNOR2_X1 U336 ( .A(n342), .B(n297), .ZN(n301) );
  XNOR2_X1 U337 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U338 ( .A(n345), .B(n407), .ZN(n346) );
  XNOR2_X1 U339 ( .A(n313), .B(n312), .ZN(n574) );
  XNOR2_X1 U340 ( .A(n555), .B(KEYINPUT55), .ZN(n556) );
  XNOR2_X1 U341 ( .A(n480), .B(KEYINPUT41), .ZN(n539) );
  XNOR2_X1 U342 ( .A(n294), .B(G106GAT), .ZN(n342) );
  NAND2_X1 U343 ( .A1(G230GAT), .A2(G233GAT), .ZN(n296) );
  XOR2_X1 U344 ( .A(KEYINPUT32), .B(KEYINPUT76), .Z(n299) );
  XNOR2_X1 U345 ( .A(KEYINPUT33), .B(KEYINPUT78), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U347 ( .A(n301), .B(n300), .Z(n313) );
  XOR2_X1 U348 ( .A(KEYINPUT75), .B(KEYINPUT31), .Z(n303) );
  XNOR2_X1 U349 ( .A(G176GAT), .B(G148GAT), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U351 ( .A(G92GAT), .B(G57GAT), .Z(n305) );
  XNOR2_X1 U352 ( .A(G120GAT), .B(G85GAT), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n311) );
  XNOR2_X1 U355 ( .A(G64GAT), .B(KEYINPUT77), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n308), .B(G204GAT), .ZN(n425) );
  XNOR2_X1 U357 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n309), .B(G78GAT), .ZN(n354) );
  XNOR2_X1 U359 ( .A(n425), .B(n354), .ZN(n310) );
  XOR2_X1 U360 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n345) );
  XNOR2_X1 U361 ( .A(G8GAT), .B(G22GAT), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n314), .B(G15GAT), .ZN(n355) );
  XOR2_X1 U363 ( .A(n345), .B(n355), .Z(n316) );
  NAND2_X1 U364 ( .A1(G229GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n332) );
  XOR2_X1 U366 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n318) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(KEYINPUT69), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n330) );
  XOR2_X1 U369 ( .A(G43GAT), .B(G36GAT), .Z(n320) );
  XNOR2_X1 U370 ( .A(G50GAT), .B(G29GAT), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n328) );
  XOR2_X1 U372 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n322) );
  XNOR2_X1 U373 ( .A(KEYINPUT70), .B(KEYINPUT68), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U375 ( .A(G141GAT), .B(G1GAT), .Z(n324) );
  XNOR2_X1 U376 ( .A(G169GAT), .B(G113GAT), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U378 ( .A(n326), .B(n325), .Z(n327) );
  XNOR2_X1 U379 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U380 ( .A(n330), .B(n329), .Z(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n537) );
  NOR2_X1 U382 ( .A1(n574), .A2(n537), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n333), .B(KEYINPUT79), .ZN(n467) );
  XOR2_X1 U384 ( .A(G29GAT), .B(G85GAT), .Z(n366) );
  XNOR2_X1 U385 ( .A(G36GAT), .B(G190GAT), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n334), .B(G92GAT), .ZN(n427) );
  XOR2_X1 U387 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n337) );
  XNOR2_X1 U388 ( .A(KEYINPUT10), .B(KEYINPUT81), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U390 ( .A(n339), .B(n338), .Z(n344) );
  XOR2_X1 U391 ( .A(KEYINPUT80), .B(G218GAT), .Z(n341) );
  XNOR2_X1 U392 ( .A(G50GAT), .B(G162GAT), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n384) );
  XNOR2_X1 U394 ( .A(n342), .B(n384), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n347) );
  XNOR2_X1 U396 ( .A(G43GAT), .B(G134GAT), .ZN(n407) );
  XOR2_X1 U397 ( .A(KEYINPUT82), .B(n507), .Z(n565) );
  XOR2_X1 U398 ( .A(G1GAT), .B(G57GAT), .Z(n365) );
  XOR2_X1 U399 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n349) );
  XNOR2_X1 U400 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U402 ( .A(G211GAT), .B(G155GAT), .Z(n351) );
  XNOR2_X1 U403 ( .A(G127GAT), .B(G183GAT), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U405 ( .A(n353), .B(n352), .Z(n357) );
  XNOR2_X1 U406 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U407 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U408 ( .A(n365), .B(n358), .Z(n360) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U410 ( .A(n360), .B(n359), .ZN(n578) );
  INV_X1 U411 ( .A(n578), .ZN(n543) );
  NOR2_X1 U412 ( .A1(n565), .A2(n543), .ZN(n361) );
  XNOR2_X1 U413 ( .A(n361), .B(KEYINPUT16), .ZN(n450) );
  XOR2_X1 U414 ( .A(KEYINPUT3), .B(G155GAT), .Z(n363) );
  XNOR2_X1 U415 ( .A(KEYINPUT2), .B(G148GAT), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U417 ( .A(G141GAT), .B(n364), .Z(n391) );
  XOR2_X1 U418 ( .A(G162GAT), .B(n365), .Z(n368) );
  XNOR2_X1 U419 ( .A(G134GAT), .B(n366), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U421 ( .A(n391), .B(n369), .Z(n371) );
  NAND2_X1 U422 ( .A1(G225GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U423 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U424 ( .A(KEYINPUT97), .B(KEYINPUT6), .Z(n373) );
  XNOR2_X1 U425 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U427 ( .A(n375), .B(n374), .Z(n383) );
  XOR2_X1 U428 ( .A(KEYINPUT0), .B(G127GAT), .Z(n377) );
  XNOR2_X1 U429 ( .A(KEYINPUT83), .B(G120GAT), .ZN(n376) );
  XNOR2_X1 U430 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U431 ( .A(G113GAT), .B(n378), .Z(n422) );
  XOR2_X1 U432 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n380) );
  XNOR2_X1 U433 ( .A(KEYINPUT5), .B(KEYINPUT100), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n422), .B(n381), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n383), .B(n382), .ZN(n441) );
  XOR2_X1 U437 ( .A(n384), .B(G106GAT), .Z(n386) );
  NAND2_X1 U438 ( .A1(G228GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U440 ( .A(n387), .B(G204GAT), .Z(n393) );
  XOR2_X1 U441 ( .A(KEYINPUT21), .B(KEYINPUT93), .Z(n389) );
  XNOR2_X1 U442 ( .A(KEYINPUT92), .B(G211GAT), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U444 ( .A(G197GAT), .B(n390), .Z(n428) );
  XNOR2_X1 U445 ( .A(n391), .B(n428), .ZN(n392) );
  XNOR2_X1 U446 ( .A(n393), .B(n392), .ZN(n401) );
  XOR2_X1 U447 ( .A(KEYINPUT22), .B(KEYINPUT95), .Z(n395) );
  XNOR2_X1 U448 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U450 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n397) );
  XNOR2_X1 U451 ( .A(G22GAT), .B(G78GAT), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U453 ( .A(n399), .B(n398), .Z(n400) );
  XNOR2_X1 U454 ( .A(n401), .B(n400), .ZN(n554) );
  XOR2_X1 U455 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n403) );
  XNOR2_X1 U456 ( .A(KEYINPUT17), .B(KEYINPUT87), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U458 ( .A(n404), .B(G183GAT), .Z(n406) );
  XNOR2_X1 U459 ( .A(G169GAT), .B(G176GAT), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n432) );
  XOR2_X1 U461 ( .A(G190GAT), .B(G99GAT), .Z(n409) );
  XOR2_X1 U462 ( .A(n407), .B(KEYINPUT88), .Z(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U464 ( .A(n432), .B(n410), .Z(n412) );
  NAND2_X1 U465 ( .A1(G227GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n412), .B(n411), .ZN(n420) );
  XOR2_X1 U467 ( .A(KEYINPUT86), .B(KEYINPUT84), .Z(n414) );
  XNOR2_X1 U468 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U470 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n416) );
  XNOR2_X1 U471 ( .A(G15GAT), .B(G71GAT), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U473 ( .A(n418), .B(n417), .Z(n419) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n557) );
  XOR2_X1 U476 ( .A(G218GAT), .B(G8GAT), .Z(n424) );
  NAND2_X1 U477 ( .A1(G226GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U479 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U482 ( .A(n432), .B(n431), .ZN(n547) );
  NOR2_X1 U483 ( .A1(n557), .A2(n547), .ZN(n433) );
  NOR2_X1 U484 ( .A1(n554), .A2(n433), .ZN(n434) );
  XOR2_X1 U485 ( .A(KEYINPUT25), .B(n434), .Z(n438) );
  NAND2_X1 U486 ( .A1(n554), .A2(n557), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n435), .B(KEYINPUT26), .ZN(n569) );
  XOR2_X1 U488 ( .A(KEYINPUT27), .B(n547), .Z(n442) );
  INV_X1 U489 ( .A(n442), .ZN(n436) );
  NOR2_X1 U490 ( .A1(n569), .A2(n436), .ZN(n437) );
  NOR2_X1 U491 ( .A1(n438), .A2(n437), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n439), .B(KEYINPUT104), .ZN(n440) );
  NOR2_X1 U493 ( .A1(n441), .A2(n440), .ZN(n448) );
  NAND2_X1 U494 ( .A1(n442), .A2(n552), .ZN(n443) );
  XOR2_X1 U495 ( .A(KEYINPUT102), .B(n443), .Z(n535) );
  XNOR2_X1 U496 ( .A(KEYINPUT67), .B(KEYINPUT28), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n444), .B(n554), .ZN(n458) );
  NAND2_X1 U498 ( .A1(n535), .A2(n458), .ZN(n519) );
  XNOR2_X1 U499 ( .A(KEYINPUT91), .B(n557), .ZN(n445) );
  NOR2_X1 U500 ( .A1(n519), .A2(n445), .ZN(n446) );
  XOR2_X1 U501 ( .A(KEYINPUT103), .B(n446), .Z(n447) );
  NOR2_X1 U502 ( .A1(n448), .A2(n447), .ZN(n463) );
  INV_X1 U503 ( .A(n463), .ZN(n449) );
  NAND2_X1 U504 ( .A1(n450), .A2(n449), .ZN(n481) );
  NOR2_X1 U505 ( .A1(n467), .A2(n481), .ZN(n451) );
  XOR2_X1 U506 ( .A(KEYINPUT105), .B(n451), .Z(n459) );
  NAND2_X1 U507 ( .A1(n459), .A2(n552), .ZN(n454) );
  XNOR2_X1 U508 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n452), .B(KEYINPUT106), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(G1324GAT) );
  INV_X1 U511 ( .A(n547), .ZN(n497) );
  NAND2_X1 U512 ( .A1(n459), .A2(n497), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n455), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U514 ( .A(G15GAT), .B(KEYINPUT35), .Z(n457) );
  INV_X1 U515 ( .A(n557), .ZN(n520) );
  NAND2_X1 U516 ( .A1(n459), .A2(n520), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n457), .B(n456), .ZN(G1326GAT) );
  XOR2_X1 U518 ( .A(G22GAT), .B(KEYINPUT107), .Z(n461) );
  INV_X1 U519 ( .A(n458), .ZN(n501) );
  NAND2_X1 U520 ( .A1(n459), .A2(n501), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n461), .B(n460), .ZN(G1327GAT) );
  XOR2_X1 U522 ( .A(G29GAT), .B(KEYINPUT108), .Z(n470) );
  XNOR2_X1 U523 ( .A(KEYINPUT110), .B(KEYINPUT37), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n462), .B(KEYINPUT109), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n565), .B(KEYINPUT36), .ZN(n511) );
  NOR2_X1 U526 ( .A1(n578), .A2(n463), .ZN(n464) );
  NAND2_X1 U527 ( .A1(n511), .A2(n464), .ZN(n465) );
  XNOR2_X1 U528 ( .A(n466), .B(n465), .ZN(n494) );
  NOR2_X1 U529 ( .A1(n467), .A2(n494), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n468), .B(KEYINPUT38), .ZN(n478) );
  NAND2_X1 U531 ( .A1(n552), .A2(n478), .ZN(n469) );
  XNOR2_X1 U532 ( .A(n470), .B(n469), .ZN(n472) );
  XOR2_X1 U533 ( .A(KEYINPUT111), .B(KEYINPUT39), .Z(n471) );
  XNOR2_X1 U534 ( .A(n472), .B(n471), .ZN(G1328GAT) );
  XNOR2_X1 U535 ( .A(G36GAT), .B(KEYINPUT112), .ZN(n474) );
  NAND2_X1 U536 ( .A1(n497), .A2(n478), .ZN(n473) );
  XNOR2_X1 U537 ( .A(n474), .B(n473), .ZN(G1329GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT113), .B(KEYINPUT40), .Z(n476) );
  NAND2_X1 U539 ( .A1(n478), .A2(n520), .ZN(n475) );
  XNOR2_X1 U540 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U541 ( .A(G43GAT), .B(n477), .ZN(G1330GAT) );
  NAND2_X1 U542 ( .A1(n478), .A2(n501), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n479), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U544 ( .A(n574), .B(KEYINPUT64), .ZN(n480) );
  INV_X1 U545 ( .A(n539), .ZN(n559) );
  NAND2_X1 U546 ( .A1(n537), .A2(n559), .ZN(n493) );
  NOR2_X1 U547 ( .A1(n493), .A2(n481), .ZN(n482) );
  XNOR2_X1 U548 ( .A(n482), .B(KEYINPUT114), .ZN(n489) );
  NAND2_X1 U549 ( .A1(n489), .A2(n552), .ZN(n486) );
  XOR2_X1 U550 ( .A(KEYINPUT115), .B(KEYINPUT42), .Z(n484) );
  XNOR2_X1 U551 ( .A(G57GAT), .B(KEYINPUT116), .ZN(n483) );
  XNOR2_X1 U552 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U553 ( .A(n486), .B(n485), .ZN(G1332GAT) );
  NAND2_X1 U554 ( .A1(n489), .A2(n497), .ZN(n487) );
  XNOR2_X1 U555 ( .A(n487), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U556 ( .A1(n489), .A2(n520), .ZN(n488) );
  XNOR2_X1 U557 ( .A(n488), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT43), .B(KEYINPUT117), .Z(n491) );
  NAND2_X1 U559 ( .A1(n501), .A2(n489), .ZN(n490) );
  XNOR2_X1 U560 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U561 ( .A(G78GAT), .B(n492), .Z(G1335GAT) );
  XNOR2_X1 U562 ( .A(G85GAT), .B(KEYINPUT118), .ZN(n496) );
  NOR2_X1 U563 ( .A1(n494), .A2(n493), .ZN(n502) );
  NAND2_X1 U564 ( .A1(n552), .A2(n502), .ZN(n495) );
  XNOR2_X1 U565 ( .A(n496), .B(n495), .ZN(G1336GAT) );
  NAND2_X1 U566 ( .A1(n502), .A2(n497), .ZN(n498) );
  XNOR2_X1 U567 ( .A(n498), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U568 ( .A(G99GAT), .B(KEYINPUT119), .Z(n500) );
  NAND2_X1 U569 ( .A1(n502), .A2(n520), .ZN(n499) );
  XNOR2_X1 U570 ( .A(n500), .B(n499), .ZN(G1338GAT) );
  NAND2_X1 U571 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U572 ( .A(n503), .B(KEYINPUT44), .ZN(n504) );
  XNOR2_X1 U573 ( .A(G106GAT), .B(n504), .ZN(G1339GAT) );
  NOR2_X1 U574 ( .A1(n537), .A2(n539), .ZN(n505) );
  XNOR2_X1 U575 ( .A(n505), .B(KEYINPUT46), .ZN(n506) );
  NOR2_X1 U576 ( .A1(n578), .A2(n506), .ZN(n508) );
  AND2_X1 U577 ( .A1(n508), .A2(n507), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(n517) );
  INV_X1 U579 ( .A(n537), .ZN(n570) );
  NAND2_X1 U580 ( .A1(n511), .A2(n578), .ZN(n514) );
  XOR2_X1 U581 ( .A(KEYINPUT66), .B(KEYINPUT120), .Z(n512) );
  XNOR2_X1 U582 ( .A(KEYINPUT45), .B(n512), .ZN(n513) );
  XNOR2_X1 U583 ( .A(n514), .B(n513), .ZN(n515) );
  NOR2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n518), .B(KEYINPUT48), .ZN(n548) );
  NOR2_X1 U586 ( .A1(n548), .A2(n519), .ZN(n521) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n530) );
  NOR2_X1 U588 ( .A1(n537), .A2(n530), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G113GAT), .B(KEYINPUT121), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(G1340GAT) );
  NOR2_X1 U591 ( .A1(n539), .A2(n530), .ZN(n525) );
  XNOR2_X1 U592 ( .A(KEYINPUT49), .B(KEYINPUT122), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U594 ( .A(G120GAT), .B(n526), .ZN(G1341GAT) );
  NOR2_X1 U595 ( .A1(n543), .A2(n530), .ZN(n528) );
  XNOR2_X1 U596 ( .A(KEYINPUT123), .B(KEYINPUT50), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n529), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT124), .B(KEYINPUT51), .Z(n533) );
  INV_X1 U600 ( .A(n530), .ZN(n531) );
  NAND2_X1 U601 ( .A1(n531), .A2(n565), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(n534), .ZN(G1343GAT) );
  NOR2_X1 U604 ( .A1(n569), .A2(n548), .ZN(n536) );
  NAND2_X1 U605 ( .A1(n536), .A2(n535), .ZN(n545) );
  NOR2_X1 U606 ( .A1(n537), .A2(n545), .ZN(n538) );
  XOR2_X1 U607 ( .A(G141GAT), .B(n538), .Z(G1344GAT) );
  NOR2_X1 U608 ( .A1(n539), .A2(n545), .ZN(n541) );
  XNOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(n542), .ZN(G1345GAT) );
  NOR2_X1 U612 ( .A1(n543), .A2(n545), .ZN(n544) );
  XOR2_X1 U613 ( .A(G155GAT), .B(n544), .Z(G1346GAT) );
  NOR2_X1 U614 ( .A1(n507), .A2(n545), .ZN(n546) );
  XOR2_X1 U615 ( .A(G162GAT), .B(n546), .Z(G1347GAT) );
  NOR2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n550) );
  INV_X1 U617 ( .A(KEYINPUT54), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT65), .ZN(n568) );
  NOR2_X1 U620 ( .A1(n568), .A2(n554), .ZN(n555) );
  NOR2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n570), .A2(n564), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n561) );
  NAND2_X1 U625 ( .A1(n564), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n564), .A2(n578), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n581) );
  NAND2_X1 U635 ( .A1(n581), .A2(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n576) );
  NAND2_X1 U639 ( .A1(n581), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  NAND2_X1 U642 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U643 ( .A(n579), .B(KEYINPUT126), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n583) );
  NAND2_X1 U646 ( .A1(n581), .A2(n511), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

