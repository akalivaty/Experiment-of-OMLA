

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U562 ( .A1(n723), .A2(n722), .ZN(n724) );
  INV_X1 U563 ( .A(n677), .ZN(n647) );
  BUF_X1 U564 ( .A(n591), .Z(n544) );
  OR2_X1 U565 ( .A1(n661), .A2(n976), .ZN(n658) );
  XNOR2_X1 U566 ( .A(KEYINPUT96), .B(KEYINPUT30), .ZN(n604) );
  XNOR2_X1 U567 ( .A(n600), .B(KEYINPUT64), .ZN(n691) );
  NOR2_X1 U568 ( .A1(n715), .A2(n717), .ZN(n528) );
  XNOR2_X1 U569 ( .A(n658), .B(KEYINPUT95), .ZN(n659) );
  XNOR2_X1 U570 ( .A(n605), .B(n604), .ZN(n606) );
  XNOR2_X1 U571 ( .A(KEYINPUT31), .B(KEYINPUT97), .ZN(n613) );
  XNOR2_X1 U572 ( .A(n614), .B(n613), .ZN(n670) );
  NAND2_X1 U573 ( .A1(G8), .A2(n677), .ZN(n717) );
  NOR2_X1 U574 ( .A1(n763), .A2(G1384), .ZN(n600) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  INV_X1 U576 ( .A(G651), .ZN(n534) );
  NOR2_X1 U577 ( .A1(G543), .A2(n534), .ZN(n529) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n529), .Z(n800) );
  NAND2_X1 U579 ( .A1(n800), .A2(G62), .ZN(n530) );
  XOR2_X1 U580 ( .A(KEYINPUT81), .B(n530), .Z(n532) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n576) );
  NOR2_X2 U582 ( .A1(n576), .A2(G651), .ZN(n808) );
  NAND2_X1 U583 ( .A1(n808), .A2(G50), .ZN(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U585 ( .A(KEYINPUT82), .B(n533), .ZN(n538) );
  NOR2_X1 U586 ( .A1(G543), .A2(G651), .ZN(n804) );
  NAND2_X1 U587 ( .A1(G88), .A2(n804), .ZN(n536) );
  NOR2_X1 U588 ( .A1(n576), .A2(n534), .ZN(n801) );
  NAND2_X1 U589 ( .A1(G75), .A2(n801), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n538), .A2(n537), .ZN(G166) );
  INV_X1 U592 ( .A(G166), .ZN(G303) );
  NAND2_X1 U593 ( .A1(n881), .A2(G113), .ZN(n541) );
  INV_X1 U594 ( .A(G2105), .ZN(n543) );
  AND2_X1 U595 ( .A1(n543), .A2(G2104), .ZN(n885) );
  NAND2_X1 U596 ( .A1(G101), .A2(n885), .ZN(n539) );
  XOR2_X1 U597 ( .A(KEYINPUT23), .B(n539), .Z(n540) );
  NAND2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n548) );
  NOR2_X1 U599 ( .A1(G2104), .A2(G2105), .ZN(n542) );
  XOR2_X1 U600 ( .A(KEYINPUT17), .B(n542), .Z(n590) );
  BUF_X1 U601 ( .A(n590), .Z(n887) );
  NAND2_X1 U602 ( .A1(G137), .A2(n887), .ZN(n546) );
  NOR2_X1 U603 ( .A1(G2104), .A2(n543), .ZN(n591) );
  NAND2_X1 U604 ( .A1(G125), .A2(n544), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U606 ( .A1(n548), .A2(n547), .ZN(G160) );
  NAND2_X1 U607 ( .A1(G63), .A2(n800), .ZN(n550) );
  NAND2_X1 U608 ( .A1(G51), .A2(n808), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U610 ( .A(KEYINPUT6), .B(n551), .ZN(n558) );
  NAND2_X1 U611 ( .A1(n804), .A2(G89), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U613 ( .A1(G76), .A2(n801), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U615 ( .A(KEYINPUT74), .B(n555), .Z(n556) );
  XNOR2_X1 U616 ( .A(KEYINPUT5), .B(n556), .ZN(n557) );
  NOR2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U618 ( .A(KEYINPUT7), .B(n559), .Z(G168) );
  NAND2_X1 U619 ( .A1(G90), .A2(n804), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G77), .A2(n801), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n563) );
  XOR2_X1 U622 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n562) );
  XNOR2_X1 U623 ( .A(n563), .B(n562), .ZN(n568) );
  NAND2_X1 U624 ( .A1(G64), .A2(n800), .ZN(n565) );
  NAND2_X1 U625 ( .A1(G52), .A2(n808), .ZN(n564) );
  NAND2_X1 U626 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U627 ( .A(KEYINPUT65), .B(n566), .Z(n567) );
  NOR2_X1 U628 ( .A1(n568), .A2(n567), .ZN(G171) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G61), .A2(n800), .ZN(n570) );
  NAND2_X1 U631 ( .A1(G86), .A2(n804), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U633 ( .A1(n801), .A2(G73), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT2), .B(n571), .Z(n572) );
  NOR2_X1 U635 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n808), .A2(G48), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(G305) );
  NAND2_X1 U638 ( .A1(G87), .A2(n576), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G49), .A2(n808), .ZN(n578) );
  NAND2_X1 U640 ( .A1(G74), .A2(G651), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U642 ( .A1(n800), .A2(n579), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U644 ( .A(n582), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U645 ( .A1(G85), .A2(n804), .ZN(n584) );
  NAND2_X1 U646 ( .A1(G72), .A2(n801), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U648 ( .A1(G60), .A2(n800), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G47), .A2(n808), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  OR2_X1 U651 ( .A1(n588), .A2(n587), .ZN(G290) );
  NOR2_X1 U652 ( .A1(G2090), .A2(G303), .ZN(n589) );
  NAND2_X1 U653 ( .A1(G8), .A2(n589), .ZN(n690) );
  NAND2_X1 U654 ( .A1(G160), .A2(G40), .ZN(n692) );
  INV_X1 U655 ( .A(n692), .ZN(n601) );
  NAND2_X1 U656 ( .A1(G138), .A2(n590), .ZN(n598) );
  NAND2_X1 U657 ( .A1(G114), .A2(n881), .ZN(n593) );
  NAND2_X1 U658 ( .A1(G126), .A2(n591), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U660 ( .A(KEYINPUT88), .B(n594), .ZN(n596) );
  AND2_X1 U661 ( .A1(G102), .A2(n885), .ZN(n595) );
  NOR2_X1 U662 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U663 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U664 ( .A(n599), .B(KEYINPUT89), .ZN(n763) );
  NAND2_X2 U665 ( .A1(n601), .A2(n691), .ZN(n677) );
  NOR2_X1 U666 ( .A1(n677), .A2(G2084), .ZN(n602) );
  NAND2_X1 U667 ( .A1(G8), .A2(n602), .ZN(n675) );
  NOR2_X1 U668 ( .A1(G1966), .A2(n717), .ZN(n673) );
  NOR2_X1 U669 ( .A1(n673), .A2(n602), .ZN(n603) );
  NAND2_X1 U670 ( .A1(n603), .A2(G8), .ZN(n605) );
  NOR2_X1 U671 ( .A1(G168), .A2(n606), .ZN(n612) );
  NAND2_X1 U672 ( .A1(n677), .A2(G1961), .ZN(n609) );
  XOR2_X1 U673 ( .A(G2078), .B(KEYINPUT25), .Z(n607) );
  XNOR2_X1 U674 ( .A(KEYINPUT92), .B(n607), .ZN(n963) );
  NAND2_X1 U675 ( .A1(n647), .A2(n963), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U677 ( .A(n610), .B(KEYINPUT93), .ZN(n666) );
  NOR2_X1 U678 ( .A1(G171), .A2(n666), .ZN(n611) );
  NOR2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U680 ( .A1(G79), .A2(n801), .ZN(n621) );
  NAND2_X1 U681 ( .A1(G66), .A2(n800), .ZN(n616) );
  NAND2_X1 U682 ( .A1(G92), .A2(n804), .ZN(n615) );
  NAND2_X1 U683 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U684 ( .A1(n808), .A2(G54), .ZN(n617) );
  XOR2_X1 U685 ( .A(KEYINPUT72), .B(n617), .Z(n618) );
  NOR2_X1 U686 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U688 ( .A(n622), .B(KEYINPUT15), .ZN(n623) );
  XOR2_X1 U689 ( .A(KEYINPUT73), .B(n623), .Z(n988) );
  NAND2_X1 U690 ( .A1(G1348), .A2(n677), .ZN(n625) );
  NAND2_X1 U691 ( .A1(G2067), .A2(n647), .ZN(n624) );
  NAND2_X1 U692 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U693 ( .A(KEYINPUT94), .B(n626), .Z(n644) );
  OR2_X1 U694 ( .A1(n988), .A2(n644), .ZN(n643) );
  XOR2_X1 U695 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n628) );
  NAND2_X1 U696 ( .A1(G56), .A2(n800), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n628), .B(n627), .ZN(n636) );
  NAND2_X1 U698 ( .A1(n804), .A2(G81), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n629), .B(KEYINPUT12), .ZN(n631) );
  NAND2_X1 U700 ( .A1(G68), .A2(n801), .ZN(n630) );
  NAND2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U702 ( .A(n632), .B(KEYINPUT13), .ZN(n634) );
  NAND2_X1 U703 ( .A1(G43), .A2(n808), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U706 ( .A(KEYINPUT71), .B(n637), .ZN(n994) );
  INV_X1 U707 ( .A(G1996), .ZN(n746) );
  NOR2_X1 U708 ( .A1(n677), .A2(n746), .ZN(n638) );
  XOR2_X1 U709 ( .A(n638), .B(KEYINPUT26), .Z(n640) );
  NAND2_X1 U710 ( .A1(n677), .A2(G1341), .ZN(n639) );
  NAND2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U712 ( .A1(n994), .A2(n641), .ZN(n642) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U714 ( .A1(n644), .A2(n988), .ZN(n645) );
  NAND2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n660) );
  NAND2_X1 U716 ( .A1(n647), .A2(G2072), .ZN(n648) );
  XOR2_X1 U717 ( .A(KEYINPUT27), .B(n648), .Z(n650) );
  NAND2_X1 U718 ( .A1(G1956), .A2(n677), .ZN(n649) );
  NAND2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n661) );
  NAND2_X1 U720 ( .A1(G65), .A2(n800), .ZN(n652) );
  NAND2_X1 U721 ( .A1(G78), .A2(n801), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U723 ( .A1(n804), .A2(G91), .ZN(n653) );
  XOR2_X1 U724 ( .A(KEYINPUT68), .B(n653), .Z(n654) );
  NOR2_X1 U725 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n808), .A2(G53), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n976) );
  NOR2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U729 ( .A1(n976), .A2(n661), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT28), .B(n662), .Z(n663) );
  NOR2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U732 ( .A(n665), .B(KEYINPUT29), .ZN(n668) );
  NAND2_X1 U733 ( .A1(n666), .A2(G171), .ZN(n667) );
  NAND2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U735 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U736 ( .A(n671), .B(KEYINPUT98), .ZN(n676) );
  INV_X1 U737 ( .A(n676), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n688) );
  NAND2_X1 U740 ( .A1(n676), .A2(G286), .ZN(n684) );
  INV_X1 U741 ( .A(G8), .ZN(n682) );
  NOR2_X1 U742 ( .A1(G1971), .A2(n717), .ZN(n679) );
  NOR2_X1 U743 ( .A1(G2090), .A2(n677), .ZN(n678) );
  NOR2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U745 ( .A1(G303), .A2(n680), .ZN(n681) );
  OR2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U747 ( .A1(n684), .A2(n683), .ZN(n686) );
  XOR2_X1 U748 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n685) );
  XNOR2_X1 U749 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U751 ( .A(KEYINPUT100), .B(n689), .ZN(n714) );
  NAND2_X1 U752 ( .A1(n690), .A2(n714), .ZN(n703) );
  NOR2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n759) );
  XNOR2_X1 U754 ( .A(G2067), .B(KEYINPUT37), .ZN(n756) );
  NAND2_X1 U755 ( .A1(G116), .A2(n881), .ZN(n694) );
  NAND2_X1 U756 ( .A1(G128), .A2(n544), .ZN(n693) );
  NAND2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U758 ( .A(n695), .B(KEYINPUT35), .ZN(n700) );
  NAND2_X1 U759 ( .A1(G104), .A2(n885), .ZN(n697) );
  NAND2_X1 U760 ( .A1(G140), .A2(n887), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U762 ( .A(KEYINPUT34), .B(n698), .Z(n699) );
  NAND2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U764 ( .A(n701), .B(KEYINPUT36), .Z(n896) );
  NOR2_X1 U765 ( .A1(n756), .A2(n896), .ZN(n935) );
  NAND2_X1 U766 ( .A1(n759), .A2(n935), .ZN(n753) );
  AND2_X1 U767 ( .A1(n717), .A2(n753), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n708) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n704) );
  XOR2_X1 U770 ( .A(n704), .B(KEYINPUT24), .Z(n705) );
  NOR2_X1 U771 ( .A1(n717), .A2(n705), .ZN(n706) );
  NAND2_X1 U772 ( .A1(n753), .A2(n706), .ZN(n707) );
  AND2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n725) );
  NOR2_X1 U774 ( .A1(G288), .A2(G1976), .ZN(n989) );
  INV_X1 U775 ( .A(n989), .ZN(n974) );
  NOR2_X1 U776 ( .A1(G1971), .A2(G303), .ZN(n709) );
  XNOR2_X1 U777 ( .A(n709), .B(KEYINPUT101), .ZN(n710) );
  AND2_X1 U778 ( .A1(n974), .A2(n710), .ZN(n712) );
  INV_X1 U779 ( .A(KEYINPUT33), .ZN(n711) );
  AND2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n713) );
  AND2_X1 U781 ( .A1(n714), .A2(n713), .ZN(n723) );
  NAND2_X1 U782 ( .A1(G288), .A2(G1976), .ZN(n990) );
  INV_X1 U783 ( .A(n990), .ZN(n715) );
  NOR2_X1 U784 ( .A1(KEYINPUT33), .A2(n528), .ZN(n719) );
  NAND2_X1 U785 ( .A1(n989), .A2(KEYINPUT33), .ZN(n716) );
  NOR2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U787 ( .A1(n719), .A2(n718), .ZN(n721) );
  XOR2_X1 U788 ( .A(G1981), .B(G305), .Z(n985) );
  AND2_X1 U789 ( .A1(n985), .A2(n753), .ZN(n720) );
  NAND2_X1 U790 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n725), .A2(n724), .ZN(n744) );
  XOR2_X1 U792 ( .A(G1986), .B(G290), .Z(n978) );
  XOR2_X1 U793 ( .A(KEYINPUT90), .B(G1991), .Z(n954) );
  NAND2_X1 U794 ( .A1(G95), .A2(n885), .ZN(n727) );
  NAND2_X1 U795 ( .A1(G107), .A2(n881), .ZN(n726) );
  NAND2_X1 U796 ( .A1(n727), .A2(n726), .ZN(n731) );
  NAND2_X1 U797 ( .A1(G131), .A2(n887), .ZN(n729) );
  NAND2_X1 U798 ( .A1(G119), .A2(n544), .ZN(n728) );
  NAND2_X1 U799 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U800 ( .A1(n731), .A2(n730), .ZN(n865) );
  NOR2_X1 U801 ( .A1(n954), .A2(n865), .ZN(n741) );
  NAND2_X1 U802 ( .A1(G105), .A2(n885), .ZN(n732) );
  XNOR2_X1 U803 ( .A(n732), .B(KEYINPUT38), .ZN(n735) );
  NAND2_X1 U804 ( .A1(G129), .A2(n544), .ZN(n733) );
  XOR2_X1 U805 ( .A(KEYINPUT91), .B(n733), .Z(n734) );
  NAND2_X1 U806 ( .A1(n735), .A2(n734), .ZN(n739) );
  NAND2_X1 U807 ( .A1(G117), .A2(n881), .ZN(n737) );
  NAND2_X1 U808 ( .A1(G141), .A2(n887), .ZN(n736) );
  NAND2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U810 ( .A1(n739), .A2(n738), .ZN(n867) );
  NOR2_X1 U811 ( .A1(n867), .A2(n746), .ZN(n740) );
  NOR2_X1 U812 ( .A1(n741), .A2(n740), .ZN(n749) );
  NAND2_X1 U813 ( .A1(n978), .A2(n749), .ZN(n742) );
  NAND2_X1 U814 ( .A1(n742), .A2(n759), .ZN(n743) );
  NAND2_X1 U815 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U816 ( .A(n745), .B(KEYINPUT102), .ZN(n761) );
  AND2_X1 U817 ( .A1(n746), .A2(n867), .ZN(n931) );
  AND2_X1 U818 ( .A1(n954), .A2(n865), .ZN(n927) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n747) );
  XOR2_X1 U820 ( .A(n747), .B(KEYINPUT103), .Z(n748) );
  NOR2_X1 U821 ( .A1(n927), .A2(n748), .ZN(n750) );
  INV_X1 U822 ( .A(n749), .ZN(n939) );
  NOR2_X1 U823 ( .A1(n750), .A2(n939), .ZN(n751) );
  NOR2_X1 U824 ( .A1(n931), .A2(n751), .ZN(n752) );
  XNOR2_X1 U825 ( .A(n752), .B(KEYINPUT39), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U827 ( .A(n755), .B(KEYINPUT104), .ZN(n757) );
  NAND2_X1 U828 ( .A1(n756), .A2(n896), .ZN(n941) );
  NAND2_X1 U829 ( .A1(n757), .A2(n941), .ZN(n758) );
  NAND2_X1 U830 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U831 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U832 ( .A(n762), .B(KEYINPUT40), .ZN(G329) );
  BUF_X1 U833 ( .A(n763), .Z(G164) );
  XOR2_X1 U834 ( .A(KEYINPUT105), .B(G2435), .Z(n765) );
  XNOR2_X1 U835 ( .A(G2430), .B(G2438), .ZN(n764) );
  XNOR2_X1 U836 ( .A(n765), .B(n764), .ZN(n772) );
  XOR2_X1 U837 ( .A(G2446), .B(G2454), .Z(n767) );
  XNOR2_X1 U838 ( .A(G2451), .B(G2443), .ZN(n766) );
  XNOR2_X1 U839 ( .A(n767), .B(n766), .ZN(n768) );
  XOR2_X1 U840 ( .A(n768), .B(G2427), .Z(n770) );
  XNOR2_X1 U841 ( .A(G1341), .B(G1348), .ZN(n769) );
  XNOR2_X1 U842 ( .A(n770), .B(n769), .ZN(n771) );
  XNOR2_X1 U843 ( .A(n772), .B(n771), .ZN(n773) );
  AND2_X1 U844 ( .A1(n773), .A2(G14), .ZN(G401) );
  INV_X1 U845 ( .A(G57), .ZN(G237) );
  INV_X1 U846 ( .A(G120), .ZN(G236) );
  INV_X1 U847 ( .A(G69), .ZN(G235) );
  NAND2_X1 U848 ( .A1(G94), .A2(G452), .ZN(n774) );
  XNOR2_X1 U849 ( .A(n774), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U850 ( .A1(G7), .A2(G661), .ZN(n775) );
  XNOR2_X1 U851 ( .A(n775), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U852 ( .A(G223), .ZN(n843) );
  NAND2_X1 U853 ( .A1(n843), .A2(G567), .ZN(n776) );
  XOR2_X1 U854 ( .A(KEYINPUT11), .B(n776), .Z(G234) );
  INV_X1 U855 ( .A(n994), .ZN(n777) );
  NAND2_X1 U856 ( .A1(n777), .A2(G860), .ZN(G153) );
  INV_X1 U857 ( .A(G171), .ZN(G301) );
  NAND2_X1 U858 ( .A1(G868), .A2(G301), .ZN(n779) );
  INV_X1 U859 ( .A(n988), .ZN(n783) );
  INV_X1 U860 ( .A(G868), .ZN(n823) );
  NAND2_X1 U861 ( .A1(n783), .A2(n823), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(G284) );
  XOR2_X1 U863 ( .A(KEYINPUT69), .B(n976), .Z(G299) );
  NAND2_X1 U864 ( .A1(G286), .A2(G868), .ZN(n781) );
  NAND2_X1 U865 ( .A1(G299), .A2(n823), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n781), .A2(n780), .ZN(G297) );
  INV_X1 U867 ( .A(G559), .ZN(n785) );
  NOR2_X1 U868 ( .A1(G860), .A2(n785), .ZN(n782) );
  NOR2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U870 ( .A(KEYINPUT16), .B(n784), .Z(G148) );
  NAND2_X1 U871 ( .A1(n785), .A2(n988), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n786), .A2(G868), .ZN(n788) );
  NAND2_X1 U873 ( .A1(n994), .A2(n823), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n788), .A2(n787), .ZN(G282) );
  XOR2_X1 U875 ( .A(KEYINPUT18), .B(KEYINPUT75), .Z(n790) );
  NAND2_X1 U876 ( .A1(G123), .A2(n544), .ZN(n789) );
  XNOR2_X1 U877 ( .A(n790), .B(n789), .ZN(n797) );
  NAND2_X1 U878 ( .A1(G99), .A2(n885), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G111), .A2(n881), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n887), .A2(G135), .ZN(n793) );
  XOR2_X1 U882 ( .A(KEYINPUT76), .B(n793), .Z(n794) );
  NOR2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n928) );
  XOR2_X1 U885 ( .A(n928), .B(G2096), .Z(n799) );
  XNOR2_X1 U886 ( .A(G2100), .B(KEYINPUT77), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(G156) );
  NAND2_X1 U888 ( .A1(G67), .A2(n800), .ZN(n803) );
  NAND2_X1 U889 ( .A1(G80), .A2(n801), .ZN(n802) );
  NAND2_X1 U890 ( .A1(n803), .A2(n802), .ZN(n807) );
  NAND2_X1 U891 ( .A1(G93), .A2(n804), .ZN(n805) );
  XNOR2_X1 U892 ( .A(KEYINPUT79), .B(n805), .ZN(n806) );
  NOR2_X1 U893 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U894 ( .A1(n808), .A2(G55), .ZN(n809) );
  NAND2_X1 U895 ( .A1(n810), .A2(n809), .ZN(n822) );
  NAND2_X1 U896 ( .A1(G559), .A2(n988), .ZN(n811) );
  XNOR2_X1 U897 ( .A(n811), .B(KEYINPUT78), .ZN(n820) );
  XNOR2_X1 U898 ( .A(n820), .B(n994), .ZN(n812) );
  NOR2_X1 U899 ( .A1(G860), .A2(n812), .ZN(n813) );
  XOR2_X1 U900 ( .A(n822), .B(n813), .Z(G145) );
  XNOR2_X1 U901 ( .A(KEYINPUT19), .B(G305), .ZN(n814) );
  XNOR2_X1 U902 ( .A(n814), .B(n822), .ZN(n817) );
  XNOR2_X1 U903 ( .A(G288), .B(n994), .ZN(n815) );
  XNOR2_X1 U904 ( .A(n815), .B(G299), .ZN(n816) );
  XNOR2_X1 U905 ( .A(n817), .B(n816), .ZN(n819) );
  XNOR2_X1 U906 ( .A(G290), .B(G166), .ZN(n818) );
  XNOR2_X1 U907 ( .A(n819), .B(n818), .ZN(n850) );
  XNOR2_X1 U908 ( .A(n820), .B(n850), .ZN(n821) );
  NAND2_X1 U909 ( .A1(n821), .A2(G868), .ZN(n825) );
  NAND2_X1 U910 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U911 ( .A1(n825), .A2(n824), .ZN(G295) );
  NAND2_X1 U912 ( .A1(G2078), .A2(G2084), .ZN(n826) );
  XNOR2_X1 U913 ( .A(n826), .B(KEYINPUT83), .ZN(n827) );
  XNOR2_X1 U914 ( .A(n827), .B(KEYINPUT20), .ZN(n828) );
  NAND2_X1 U915 ( .A1(n828), .A2(G2090), .ZN(n829) );
  XNOR2_X1 U916 ( .A(KEYINPUT21), .B(n829), .ZN(n830) );
  NAND2_X1 U917 ( .A1(n830), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U918 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U919 ( .A1(G132), .A2(G82), .ZN(n831) );
  XNOR2_X1 U920 ( .A(n831), .B(KEYINPUT84), .ZN(n832) );
  XNOR2_X1 U921 ( .A(n832), .B(KEYINPUT22), .ZN(n833) );
  NOR2_X1 U922 ( .A1(G218), .A2(n833), .ZN(n834) );
  NAND2_X1 U923 ( .A1(G96), .A2(n834), .ZN(n924) );
  NAND2_X1 U924 ( .A1(n924), .A2(G2106), .ZN(n839) );
  NOR2_X1 U925 ( .A1(G235), .A2(G236), .ZN(n835) );
  NAND2_X1 U926 ( .A1(G108), .A2(n835), .ZN(n836) );
  NOR2_X1 U927 ( .A1(n836), .A2(G237), .ZN(n837) );
  XNOR2_X1 U928 ( .A(n837), .B(KEYINPUT85), .ZN(n923) );
  NAND2_X1 U929 ( .A1(n923), .A2(G567), .ZN(n838) );
  NAND2_X1 U930 ( .A1(n839), .A2(n838), .ZN(n849) );
  NAND2_X1 U931 ( .A1(G661), .A2(G483), .ZN(n840) );
  XNOR2_X1 U932 ( .A(KEYINPUT86), .B(n840), .ZN(n841) );
  NOR2_X1 U933 ( .A1(n849), .A2(n841), .ZN(n846) );
  NAND2_X1 U934 ( .A1(n846), .A2(G36), .ZN(n842) );
  XOR2_X1 U935 ( .A(KEYINPUT87), .B(n842), .Z(G176) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U938 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n845) );
  XNOR2_X1 U940 ( .A(KEYINPUT106), .B(n845), .ZN(n847) );
  NAND2_X1 U941 ( .A1(n847), .A2(n846), .ZN(n848) );
  XOR2_X1 U942 ( .A(KEYINPUT107), .B(n848), .Z(G188) );
  INV_X1 U943 ( .A(n849), .ZN(G319) );
  XOR2_X1 U944 ( .A(n850), .B(G286), .Z(n852) );
  XNOR2_X1 U945 ( .A(G171), .B(n988), .ZN(n851) );
  XNOR2_X1 U946 ( .A(n852), .B(n851), .ZN(n853) );
  NOR2_X1 U947 ( .A1(G37), .A2(n853), .ZN(G397) );
  NAND2_X1 U948 ( .A1(G100), .A2(n885), .ZN(n854) );
  XNOR2_X1 U949 ( .A(n854), .B(KEYINPUT110), .ZN(n858) );
  XOR2_X1 U950 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n856) );
  NAND2_X1 U951 ( .A1(G124), .A2(n544), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n856), .B(n855), .ZN(n857) );
  NAND2_X1 U953 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U954 ( .A1(G112), .A2(n881), .ZN(n860) );
  NAND2_X1 U955 ( .A1(G136), .A2(n887), .ZN(n859) );
  NAND2_X1 U956 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U957 ( .A1(n862), .A2(n861), .ZN(G162) );
  XOR2_X1 U958 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n864) );
  XNOR2_X1 U959 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(n866) );
  XOR2_X1 U961 ( .A(n866), .B(n865), .Z(n869) );
  XNOR2_X1 U962 ( .A(G160), .B(n867), .ZN(n868) );
  XNOR2_X1 U963 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U964 ( .A(G162), .B(n870), .Z(n871) );
  XNOR2_X1 U965 ( .A(n928), .B(n871), .ZN(n880) );
  NAND2_X1 U966 ( .A1(G118), .A2(n881), .ZN(n873) );
  NAND2_X1 U967 ( .A1(G130), .A2(n544), .ZN(n872) );
  NAND2_X1 U968 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U969 ( .A1(G106), .A2(n885), .ZN(n875) );
  NAND2_X1 U970 ( .A1(G142), .A2(n887), .ZN(n874) );
  NAND2_X1 U971 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U972 ( .A(KEYINPUT45), .B(n876), .Z(n877) );
  NOR2_X1 U973 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U974 ( .A(n880), .B(n879), .Z(n895) );
  NAND2_X1 U975 ( .A1(G115), .A2(n881), .ZN(n883) );
  NAND2_X1 U976 ( .A1(G127), .A2(n544), .ZN(n882) );
  NAND2_X1 U977 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U978 ( .A(n884), .B(KEYINPUT47), .ZN(n892) );
  NAND2_X1 U979 ( .A1(n885), .A2(G103), .ZN(n886) );
  XOR2_X1 U980 ( .A(KEYINPUT111), .B(n886), .Z(n889) );
  NAND2_X1 U981 ( .A1(n887), .A2(G139), .ZN(n888) );
  NAND2_X1 U982 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U983 ( .A(KEYINPUT112), .B(n890), .Z(n891) );
  NAND2_X1 U984 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U985 ( .A(n893), .B(KEYINPUT113), .ZN(n945) );
  XNOR2_X1 U986 ( .A(G164), .B(n945), .ZN(n894) );
  XNOR2_X1 U987 ( .A(n895), .B(n894), .ZN(n897) );
  XNOR2_X1 U988 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U989 ( .A1(G37), .A2(n898), .ZN(G395) );
  XOR2_X1 U990 ( .A(G2096), .B(G2100), .Z(n900) );
  XNOR2_X1 U991 ( .A(KEYINPUT42), .B(G2678), .ZN(n899) );
  XNOR2_X1 U992 ( .A(n900), .B(n899), .ZN(n904) );
  XOR2_X1 U993 ( .A(KEYINPUT43), .B(G2072), .Z(n902) );
  XNOR2_X1 U994 ( .A(G2067), .B(G2090), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U996 ( .A(n904), .B(n903), .Z(n906) );
  XNOR2_X1 U997 ( .A(G2078), .B(G2084), .ZN(n905) );
  XNOR2_X1 U998 ( .A(n906), .B(n905), .ZN(G227) );
  XOR2_X1 U999 ( .A(G1976), .B(G1981), .Z(n908) );
  XNOR2_X1 U1000 ( .A(G1961), .B(G1956), .ZN(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1002 ( .A(n909), .B(KEYINPUT41), .Z(n911) );
  XNOR2_X1 U1003 ( .A(G1996), .B(G1991), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1005 ( .A(G2474), .B(G1971), .Z(n913) );
  XNOR2_X1 U1006 ( .A(G1986), .B(G1966), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(n915), .B(n914), .ZN(G229) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n916) );
  XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n916), .Z(n917) );
  XNOR2_X1 U1011 ( .A(KEYINPUT116), .B(n917), .ZN(n922) );
  NOR2_X1 U1012 ( .A1(G397), .A2(G395), .ZN(n918) );
  XOR2_X1 U1013 ( .A(KEYINPUT117), .B(n918), .Z(n919) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n919), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n920), .ZN(n921) );
  NAND2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(G225) );
  XOR2_X1 U1017 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  XNOR2_X1 U1018 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U1020 ( .A(G132), .ZN(G219) );
  INV_X1 U1021 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(KEYINPUT108), .ZN(G325) );
  INV_X1 U1024 ( .A(G325), .ZN(G261) );
  INV_X1 U1025 ( .A(G96), .ZN(G221) );
  XOR2_X1 U1026 ( .A(G160), .B(G2084), .Z(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n934) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(KEYINPUT51), .B(n932), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n937) );
  INV_X1 U1033 ( .A(n935), .ZN(n936) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(n940), .B(KEYINPUT120), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1038 ( .A(KEYINPUT121), .B(n943), .Z(n950) );
  XOR2_X1 U1039 ( .A(G164), .B(G2078), .Z(n944) );
  XNOR2_X1 U1040 ( .A(KEYINPUT122), .B(n944), .ZN(n947) );
  XOR2_X1 U1041 ( .A(G2072), .B(n945), .Z(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1043 ( .A(KEYINPUT50), .B(n948), .Z(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(KEYINPUT52), .B(n951), .ZN(n952) );
  INV_X1 U1046 ( .A(KEYINPUT55), .ZN(n1026) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n1026), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n953), .A2(G29), .ZN(n1035) );
  XNOR2_X1 U1049 ( .A(G2090), .B(G35), .ZN(n968) );
  XNOR2_X1 U1050 ( .A(n954), .B(G25), .ZN(n962) );
  XNOR2_X1 U1051 ( .A(G2067), .B(G26), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G32), .B(G1996), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(G28), .A2(n957), .ZN(n960) );
  XOR2_X1 U1055 ( .A(G33), .B(G2072), .Z(n958) );
  XNOR2_X1 U1056 ( .A(KEYINPUT123), .B(n958), .ZN(n959) );
  NOR2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(G27), .B(n963), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(KEYINPUT53), .B(n966), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n971) );
  XOR2_X1 U1063 ( .A(G2084), .B(G34), .Z(n969) );
  XNOR2_X1 U1064 ( .A(KEYINPUT54), .B(n969), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n1027) );
  NOR2_X1 U1066 ( .A1(G29), .A2(KEYINPUT55), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n1027), .A2(n972), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(G11), .A2(n973), .ZN(n1033) );
  XNOR2_X1 U1069 ( .A(G16), .B(KEYINPUT56), .ZN(n1004) );
  XNOR2_X1 U1070 ( .A(G166), .B(G1971), .ZN(n1002) );
  NAND2_X1 U1071 ( .A1(n990), .A2(n974), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n975), .A2(KEYINPUT126), .ZN(n983) );
  XOR2_X1 U1073 ( .A(G1956), .B(n976), .Z(n977) );
  NAND2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n981) );
  XOR2_X1 U1075 ( .A(G1961), .B(G301), .Z(n979) );
  XNOR2_X1 U1076 ( .A(KEYINPUT125), .B(n979), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n1000) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G168), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(n984), .B(KEYINPUT124), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(n987), .B(KEYINPUT57), .ZN(n998) );
  XNOR2_X1 U1083 ( .A(n988), .B(G1348), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n989), .A2(KEYINPUT126), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(G1341), .B(n994), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1031) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G21), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G5), .B(G1961), .ZN(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1016) );
  XOR2_X1 U1096 ( .A(G1348), .B(KEYINPUT59), .Z(n1007) );
  XNOR2_X1 U1097 ( .A(G4), .B(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(G20), .B(G1956), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G1341), .B(G19), .ZN(n1011) );
  XNOR2_X1 U1101 ( .A(G1981), .B(G6), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1014), .Z(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(G23), .B(G1976), .ZN(n1017) );
  NOR2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1109 ( .A(G1986), .B(G24), .Z(n1019) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1024), .Z(n1025) );
  NOR2_X1 U1114 ( .A1(G16), .A2(n1025), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1120 ( .A(n1036), .B(KEYINPUT62), .ZN(n1037) );
  XNOR2_X1 U1121 ( .A(KEYINPUT127), .B(n1037), .ZN(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

