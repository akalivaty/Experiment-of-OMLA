

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579;

  XNOR2_X1 U320 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U321 ( .A(n392), .B(n391), .ZN(n536) );
  XNOR2_X1 U322 ( .A(n336), .B(n335), .ZN(n340) );
  XNOR2_X1 U323 ( .A(KEYINPUT100), .B(KEYINPUT36), .ZN(n341) );
  XNOR2_X1 U324 ( .A(n390), .B(KEYINPUT48), .ZN(n391) );
  XNOR2_X1 U325 ( .A(n532), .B(n341), .ZN(n479) );
  XNOR2_X1 U326 ( .A(n334), .B(n394), .ZN(n335) );
  XNOR2_X1 U327 ( .A(n376), .B(n375), .ZN(n377) );
  INV_X1 U328 ( .A(G190GAT), .ZN(n447) );
  XNOR2_X1 U329 ( .A(n304), .B(n303), .ZN(n514) );
  XNOR2_X1 U330 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U331 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(G176GAT), .B(G190GAT), .Z(n289) );
  XNOR2_X1 U333 ( .A(G169GAT), .B(G99GAT), .ZN(n288) );
  XNOR2_X1 U334 ( .A(n289), .B(n288), .ZN(n293) );
  XOR2_X1 U335 ( .A(KEYINPUT87), .B(G71GAT), .Z(n291) );
  XNOR2_X1 U336 ( .A(KEYINPUT20), .B(KEYINPUT88), .ZN(n290) );
  XNOR2_X1 U337 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n293), .B(n292), .ZN(n304) );
  XOR2_X1 U339 ( .A(G43GAT), .B(G134GAT), .Z(n331) );
  XOR2_X1 U340 ( .A(G183GAT), .B(KEYINPUT17), .Z(n295) );
  XNOR2_X1 U341 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n295), .B(n294), .ZN(n395) );
  XOR2_X1 U343 ( .A(n331), .B(n395), .Z(n297) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U345 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U346 ( .A(n298), .B(KEYINPUT86), .Z(n302) );
  XOR2_X1 U347 ( .A(G120GAT), .B(G127GAT), .Z(n300) );
  XNOR2_X1 U348 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n416) );
  XNOR2_X1 U350 ( .A(G15GAT), .B(n416), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U352 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n306) );
  NAND2_X1 U353 ( .A1(G230GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n308) );
  INV_X1 U355 ( .A(KEYINPUT33), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n313) );
  XOR2_X1 U357 ( .A(KEYINPUT74), .B(G64GAT), .Z(n310) );
  XNOR2_X1 U358 ( .A(G176GAT), .B(G204GAT), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n397) );
  XNOR2_X1 U360 ( .A(G71GAT), .B(G57GAT), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n311), .B(KEYINPUT13), .ZN(n355) );
  XNOR2_X1 U362 ( .A(n397), .B(n355), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U364 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n315) );
  XNOR2_X1 U365 ( .A(G120GAT), .B(G92GAT), .ZN(n314) );
  XOR2_X1 U366 ( .A(n315), .B(n314), .Z(n316) );
  XNOR2_X1 U367 ( .A(n317), .B(n316), .ZN(n323) );
  XOR2_X1 U368 ( .A(G78GAT), .B(G148GAT), .Z(n319) );
  XNOR2_X1 U369 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n440) );
  XOR2_X1 U371 ( .A(G85GAT), .B(KEYINPUT72), .Z(n321) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(G106GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n328) );
  XNOR2_X1 U374 ( .A(n440), .B(n328), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n570) );
  XOR2_X1 U376 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n325) );
  NAND2_X1 U377 ( .A1(G232GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n326), .B(KEYINPUT77), .ZN(n330) );
  XNOR2_X1 U380 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n327), .B(KEYINPUT8), .ZN(n367) );
  XNOR2_X1 U382 ( .A(n367), .B(n328), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n336) );
  XOR2_X1 U384 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  XNOR2_X1 U385 ( .A(n331), .B(n428), .ZN(n334) );
  XOR2_X1 U386 ( .A(G92GAT), .B(G218GAT), .Z(n333) );
  XNOR2_X1 U387 ( .A(G36GAT), .B(G190GAT), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n394) );
  XOR2_X1 U389 ( .A(KEYINPUT10), .B(KEYINPUT68), .Z(n338) );
  XNOR2_X1 U390 ( .A(KEYINPUT9), .B(KEYINPUT75), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n553) );
  XNOR2_X1 U393 ( .A(KEYINPUT78), .B(n553), .ZN(n532) );
  XOR2_X1 U394 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n343) );
  XNOR2_X1 U395 ( .A(G8GAT), .B(KEYINPUT79), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n360) );
  XOR2_X1 U397 ( .A(G211GAT), .B(G78GAT), .Z(n345) );
  XNOR2_X1 U398 ( .A(G127GAT), .B(G183GAT), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U400 ( .A(KEYINPUT82), .B(KEYINPUT12), .Z(n347) );
  XNOR2_X1 U401 ( .A(KEYINPUT80), .B(KEYINPUT14), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U403 ( .A(n349), .B(n348), .Z(n354) );
  XOR2_X1 U404 ( .A(KEYINPUT83), .B(G64GAT), .Z(n351) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U407 ( .A(KEYINPUT84), .B(n352), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n356) );
  XOR2_X1 U409 ( .A(n356), .B(n355), .Z(n358) );
  XOR2_X1 U410 ( .A(G15GAT), .B(G1GAT), .Z(n372) );
  XOR2_X1 U411 ( .A(G22GAT), .B(G155GAT), .Z(n436) );
  XNOR2_X1 U412 ( .A(n372), .B(n436), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n575) );
  AND2_X1 U415 ( .A1(n479), .A2(n575), .ZN(n363) );
  XOR2_X1 U416 ( .A(KEYINPUT117), .B(KEYINPUT45), .Z(n361) );
  XNOR2_X1 U417 ( .A(KEYINPUT67), .B(n361), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n364) );
  NOR2_X1 U419 ( .A1(n570), .A2(n364), .ZN(n379) );
  XOR2_X1 U420 ( .A(G113GAT), .B(G36GAT), .Z(n366) );
  XNOR2_X1 U421 ( .A(G50GAT), .B(G43GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n378) );
  XNOR2_X1 U423 ( .A(n367), .B(KEYINPUT29), .ZN(n369) );
  AND2_X1 U424 ( .A1(G229GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n376) );
  XOR2_X1 U426 ( .A(KEYINPUT30), .B(G197GAT), .Z(n371) );
  XNOR2_X1 U427 ( .A(G22GAT), .B(G141GAT), .ZN(n370) );
  XOR2_X1 U428 ( .A(n371), .B(n370), .Z(n374) );
  XOR2_X1 U429 ( .A(G169GAT), .B(G8GAT), .Z(n396) );
  XNOR2_X1 U430 ( .A(n372), .B(n396), .ZN(n373) );
  XOR2_X1 U431 ( .A(n378), .B(n377), .Z(n565) );
  INV_X1 U432 ( .A(n565), .ZN(n539) );
  NAND2_X1 U433 ( .A1(n379), .A2(n539), .ZN(n389) );
  XNOR2_X1 U434 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n380) );
  XNOR2_X1 U435 ( .A(n570), .B(n380), .ZN(n556) );
  NAND2_X1 U436 ( .A1(n556), .A2(n565), .ZN(n382) );
  XOR2_X1 U437 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n383) );
  NOR2_X1 U439 ( .A1(n383), .A2(n575), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n384), .B(KEYINPUT115), .ZN(n385) );
  NOR2_X1 U441 ( .A1(n553), .A2(n385), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n386), .B(KEYINPUT47), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n387), .B(KEYINPUT116), .ZN(n388) );
  NAND2_X1 U444 ( .A1(n389), .A2(n388), .ZN(n392) );
  INV_X1 U445 ( .A(KEYINPUT64), .ZN(n390) );
  XNOR2_X1 U446 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n393), .B(G211GAT), .ZN(n427) );
  XNOR2_X1 U448 ( .A(n395), .B(n394), .ZN(n401) );
  XOR2_X1 U449 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U453 ( .A(n427), .B(n402), .ZN(n510) );
  NOR2_X1 U454 ( .A1(n536), .A2(n510), .ZN(n403) );
  XNOR2_X1 U455 ( .A(n403), .B(KEYINPUT54), .ZN(n425) );
  XOR2_X1 U456 ( .A(KEYINPUT90), .B(KEYINPUT2), .Z(n405) );
  XNOR2_X1 U457 ( .A(KEYINPUT3), .B(KEYINPUT91), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U459 ( .A(G141GAT), .B(n406), .Z(n432) );
  XOR2_X1 U460 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n408) );
  NAND2_X1 U461 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U462 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U463 ( .A(KEYINPUT94), .B(n409), .ZN(n423) );
  XOR2_X1 U464 ( .A(KEYINPUT1), .B(KEYINPUT93), .Z(n411) );
  XNOR2_X1 U465 ( .A(G148GAT), .B(G155GAT), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U467 ( .A(KEYINPUT95), .B(G57GAT), .Z(n413) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U470 ( .A(n415), .B(n414), .Z(n421) );
  XOR2_X1 U471 ( .A(G85GAT), .B(G162GAT), .Z(n418) );
  XNOR2_X1 U472 ( .A(n416), .B(G134GAT), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U477 ( .A(n432), .B(n424), .ZN(n507) );
  NAND2_X1 U478 ( .A1(n425), .A2(n507), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n426), .B(KEYINPUT66), .ZN(n563) );
  XOR2_X1 U480 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U483 ( .A(n432), .B(n431), .ZN(n444) );
  XOR2_X1 U484 ( .A(G204GAT), .B(KEYINPUT92), .Z(n434) );
  XNOR2_X1 U485 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U487 ( .A(n435), .B(G106GAT), .Z(n438) );
  XNOR2_X1 U488 ( .A(n436), .B(G218GAT), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U490 ( .A(n439), .B(KEYINPUT89), .Z(n442) );
  XNOR2_X1 U491 ( .A(n440), .B(KEYINPUT24), .ZN(n441) );
  XNOR2_X1 U492 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U493 ( .A(n444), .B(n443), .ZN(n461) );
  NOR2_X1 U494 ( .A1(n563), .A2(n461), .ZN(n445) );
  XNOR2_X1 U495 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  NOR2_X2 U496 ( .A1(n514), .A2(n446), .ZN(n561) );
  NAND2_X1 U497 ( .A1(n561), .A2(n532), .ZN(n450) );
  XOR2_X1 U498 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n448) );
  NOR2_X1 U499 ( .A1(n570), .A2(n539), .ZN(n482) );
  INV_X1 U500 ( .A(n507), .ZN(n459) );
  NOR2_X1 U501 ( .A1(n514), .A2(n510), .ZN(n451) );
  NOR2_X1 U502 ( .A1(n461), .A2(n451), .ZN(n452) );
  XNOR2_X1 U503 ( .A(n452), .B(KEYINPUT25), .ZN(n453) );
  XNOR2_X1 U504 ( .A(n453), .B(KEYINPUT97), .ZN(n457) );
  NAND2_X1 U505 ( .A1(n461), .A2(n514), .ZN(n454) );
  XNOR2_X1 U506 ( .A(n454), .B(KEYINPUT26), .ZN(n564) );
  XNOR2_X1 U507 ( .A(KEYINPUT27), .B(n510), .ZN(n460) );
  NOR2_X1 U508 ( .A1(n564), .A2(n460), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n455), .B(KEYINPUT96), .ZN(n456) );
  NOR2_X1 U510 ( .A1(n457), .A2(n456), .ZN(n458) );
  NOR2_X1 U511 ( .A1(n459), .A2(n458), .ZN(n463) );
  NOR2_X1 U512 ( .A1(n460), .A2(n507), .ZN(n538) );
  XOR2_X1 U513 ( .A(n461), .B(KEYINPUT28), .Z(n518) );
  NAND2_X1 U514 ( .A1(n538), .A2(n518), .ZN(n522) );
  INV_X1 U515 ( .A(n514), .ZN(n523) );
  NOR2_X1 U516 ( .A1(n522), .A2(n523), .ZN(n462) );
  NOR2_X1 U517 ( .A1(n463), .A2(n462), .ZN(n477) );
  XNOR2_X1 U518 ( .A(KEYINPUT85), .B(KEYINPUT16), .ZN(n465) );
  INV_X1 U519 ( .A(n575), .ZN(n548) );
  NOR2_X1 U520 ( .A1(n532), .A2(n548), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n465), .B(n464), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n477), .A2(n466), .ZN(n495) );
  NAND2_X1 U523 ( .A1(n482), .A2(n495), .ZN(n473) );
  NOR2_X1 U524 ( .A1(n507), .A2(n473), .ZN(n467) );
  XOR2_X1 U525 ( .A(KEYINPUT34), .B(n467), .Z(n468) );
  XNOR2_X1 U526 ( .A(G1GAT), .B(n468), .ZN(G1324GAT) );
  NOR2_X1 U527 ( .A1(n510), .A2(n473), .ZN(n469) );
  XOR2_X1 U528 ( .A(G8GAT), .B(n469), .Z(G1325GAT) );
  NOR2_X1 U529 ( .A1(n514), .A2(n473), .ZN(n471) );
  XNOR2_X1 U530 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U532 ( .A(G15GAT), .B(n472), .ZN(G1326GAT) );
  NOR2_X1 U533 ( .A1(n518), .A2(n473), .ZN(n474) );
  XOR2_X1 U534 ( .A(G22GAT), .B(n474), .Z(G1327GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n476) );
  XNOR2_X1 U536 ( .A(G29GAT), .B(KEYINPUT99), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(n486) );
  XNOR2_X1 U538 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n484) );
  NOR2_X1 U539 ( .A1(n477), .A2(n575), .ZN(n478) );
  XOR2_X1 U540 ( .A(KEYINPUT101), .B(n478), .Z(n480) );
  NAND2_X1 U541 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(KEYINPUT37), .ZN(n506) );
  NAND2_X1 U543 ( .A1(n506), .A2(n482), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n491) );
  NOR2_X1 U545 ( .A1(n507), .A2(n491), .ZN(n485) );
  XOR2_X1 U546 ( .A(n486), .B(n485), .Z(G1328GAT) );
  NOR2_X1 U547 ( .A1(n510), .A2(n491), .ZN(n487) );
  XOR2_X1 U548 ( .A(G36GAT), .B(n487), .Z(G1329GAT) );
  NOR2_X1 U549 ( .A1(n514), .A2(n491), .ZN(n489) );
  XNOR2_X1 U550 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U552 ( .A(G43GAT), .B(n490), .Z(G1330GAT) );
  NOR2_X1 U553 ( .A1(n518), .A2(n491), .ZN(n492) );
  XOR2_X1 U554 ( .A(G50GAT), .B(n492), .Z(G1331GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n494) );
  XNOR2_X1 U556 ( .A(G57GAT), .B(KEYINPUT105), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(n497) );
  INV_X1 U558 ( .A(n556), .ZN(n543) );
  NOR2_X1 U559 ( .A1(n565), .A2(n543), .ZN(n505) );
  NAND2_X1 U560 ( .A1(n505), .A2(n495), .ZN(n501) );
  NOR2_X1 U561 ( .A1(n507), .A2(n501), .ZN(n496) );
  XOR2_X1 U562 ( .A(n497), .B(n496), .Z(G1332GAT) );
  NOR2_X1 U563 ( .A1(n510), .A2(n501), .ZN(n499) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n498) );
  XNOR2_X1 U565 ( .A(n499), .B(n498), .ZN(G1333GAT) );
  NOR2_X1 U566 ( .A1(n514), .A2(n501), .ZN(n500) );
  XOR2_X1 U567 ( .A(G71GAT), .B(n500), .Z(G1334GAT) );
  NOR2_X1 U568 ( .A1(n518), .A2(n501), .ZN(n503) );
  XNOR2_X1 U569 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(n504), .ZN(G1335GAT) );
  NAND2_X1 U572 ( .A1(n506), .A2(n505), .ZN(n517) );
  NOR2_X1 U573 ( .A1(n507), .A2(n517), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1336GAT) );
  NOR2_X1 U576 ( .A1(n510), .A2(n517), .ZN(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G92GAT), .B(n513), .ZN(G1337GAT) );
  NOR2_X1 U580 ( .A1(n514), .A2(n517), .ZN(n515) );
  XOR2_X1 U581 ( .A(KEYINPUT112), .B(n515), .Z(n516) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(n516), .ZN(G1338GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n520) );
  XNOR2_X1 U584 ( .A(KEYINPUT113), .B(KEYINPUT44), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n536), .A2(n522), .ZN(n524) );
  NAND2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n531) );
  NOR2_X1 U589 ( .A1(n539), .A2(n531), .ZN(n525) );
  XOR2_X1 U590 ( .A(G113GAT), .B(n525), .Z(G1340GAT) );
  NOR2_X1 U591 ( .A1(n543), .A2(n531), .ZN(n527) );
  XNOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(G1341GAT) );
  NOR2_X1 U594 ( .A1(n548), .A2(n531), .ZN(n529) );
  XNOR2_X1 U595 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U597 ( .A(G127GAT), .B(n530), .Z(G1342GAT) );
  XOR2_X1 U598 ( .A(G134GAT), .B(KEYINPUT51), .Z(n535) );
  INV_X1 U599 ( .A(n531), .ZN(n533) );
  NAND2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(G1343GAT) );
  NOR2_X1 U602 ( .A1(n536), .A2(n564), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n551) );
  NOR2_X1 U604 ( .A1(n539), .A2(n551), .ZN(n540) );
  XOR2_X1 U605 ( .A(G141GAT), .B(n540), .Z(G1344GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n542) );
  XNOR2_X1 U607 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n547) );
  NOR2_X1 U609 ( .A1(n543), .A2(n551), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(n547), .B(n546), .Z(G1345GAT) );
  NOR2_X1 U613 ( .A1(n548), .A2(n551), .ZN(n549) );
  XOR2_X1 U614 ( .A(KEYINPUT122), .B(n549), .Z(n550) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  INV_X1 U616 ( .A(n551), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U619 ( .A1(n561), .A2(n565), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n558) );
  NAND2_X1 U622 ( .A1(n561), .A2(n556), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n560) );
  XOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT123), .Z(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U626 ( .A1(n575), .A2(n561), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT60), .Z(n567) );
  NOR2_X1 U629 ( .A1(n563), .A2(n564), .ZN(n577) );
  NAND2_X1 U630 ( .A1(n577), .A2(n565), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n568) );
  XNOR2_X1 U633 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n572) );
  NAND2_X1 U635 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n572), .B(n571), .ZN(n574) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT126), .Z(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n577), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n479), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

