//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G101), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n192), .A2(new_n195), .A3(new_n199), .A4(new_n196), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(KEYINPUT4), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT4), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n202), .A3(G101), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G113), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT2), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G113), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT66), .A2(G119), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT66), .A2(G119), .ZN(new_n212));
  INV_X1    g026(.A(G116), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G119), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT67), .B1(new_n215), .B2(G116), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n213), .A3(G119), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n210), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT68), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n215), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT66), .A2(G119), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(G116), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n218), .A3(new_n216), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n210), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n225), .A2(new_n209), .A3(new_n218), .A4(new_n216), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n216), .A2(new_n218), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(KEYINPUT69), .A3(new_n209), .A4(new_n225), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n204), .B1(new_n229), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n191), .A2(G107), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n194), .A2(G104), .ZN(new_n238));
  OAI21_X1  g052(.A(G101), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n200), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT5), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n205), .B1(new_n214), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n241), .B2(new_n226), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n235), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n190), .B1(new_n236), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n235), .A2(new_n240), .A3(new_n243), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n221), .A2(new_n228), .B1(new_n232), .B2(new_n234), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n246), .B(new_n189), .C1(new_n247), .C2(new_n204), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(KEYINPUT6), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT6), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n250), .B(new_n190), .C1(new_n236), .C2(new_n244), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT1), .B1(new_n252), .B2(G146), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(G146), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G143), .ZN(new_n256));
  OAI211_X1 g070(.A(G128), .B(new_n253), .C1(new_n254), .C2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G125), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n252), .A2(G146), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n259), .B(new_n260), .C1(KEYINPUT1), .C2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT0), .A4(G128), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n254), .A2(new_n256), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G128), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n263), .B1(new_n267), .B2(new_n258), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G224), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n268), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n249), .A2(new_n251), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G902), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n189), .B(KEYINPUT8), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n240), .B1(new_n235), .B2(new_n243), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n244), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT82), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT82), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n278), .B(new_n274), .C1(new_n244), .C2(new_n275), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n270), .A2(KEYINPUT7), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(KEYINPUT83), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n268), .A2(new_n282), .ZN(new_n283));
  OAI221_X1 g097(.A(new_n263), .B1(KEYINPUT83), .B2(new_n281), .C1(new_n267), .C2(new_n258), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n283), .A2(new_n284), .B1(KEYINPUT83), .B2(new_n281), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n277), .A2(new_n248), .A3(new_n279), .A4(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n272), .A2(new_n273), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G210), .B1(G237), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n272), .A2(new_n286), .A3(new_n273), .A4(new_n288), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n188), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(KEYINPUT84), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT84), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n294), .B(new_n188), .C1(new_n290), .C2(new_n291), .ZN(new_n295));
  XNOR2_X1  g109(.A(G110), .B(G140), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n269), .A2(G227), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT11), .ZN(new_n299));
  INV_X1    g113(.A(G134), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(G137), .ZN(new_n301));
  INV_X1    g115(.A(G137), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT11), .A3(G134), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(G137), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G131), .ZN(new_n306));
  INV_X1    g120(.A(G131), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n301), .A2(new_n303), .A3(new_n307), .A4(new_n304), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n306), .A2(KEYINPUT70), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT70), .B1(new_n306), .B2(new_n308), .ZN(new_n310));
  AND4_X1   g124(.A1(new_n262), .A2(new_n257), .A3(new_n200), .A4(new_n239), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n262), .A2(new_n257), .B1(new_n200), .B2(new_n239), .ZN(new_n312));
  OAI22_X1  g126(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT12), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n257), .A2(new_n262), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n200), .A2(new_n239), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n315), .B(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n314), .B1(new_n306), .B2(new_n308), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n313), .A2(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n267), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n201), .A2(new_n320), .A3(new_n203), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n257), .A2(new_n262), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n240), .A3(KEYINPUT10), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n315), .B2(new_n316), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n306), .A2(new_n308), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT70), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n306), .A2(KEYINPUT70), .A3(new_n308), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n298), .B1(new_n319), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n326), .A2(new_n331), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n309), .A2(new_n310), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n335), .A2(new_n321), .A3(new_n323), .A4(new_n325), .ZN(new_n336));
  INV_X1    g150(.A(new_n298), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(G469), .B1(new_n340), .B2(G902), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n334), .A2(new_n336), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n298), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n317), .A2(new_n318), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT12), .B1(new_n317), .B2(new_n331), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n336), .B(new_n337), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(G902), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G469), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n342), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n337), .B1(new_n326), .B2(new_n331), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(new_n319), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n337), .B1(new_n334), .B2(new_n336), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n349), .B(new_n273), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(KEYINPUT81), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n341), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G221), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT9), .B(G234), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT79), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n360), .B2(new_n273), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n356), .A2(new_n362), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n293), .A2(new_n295), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT89), .ZN(new_n365));
  INV_X1    g179(.A(G217), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n359), .A2(new_n366), .A3(G953), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n213), .A2(KEYINPUT14), .A3(G122), .ZN(new_n368));
  INV_X1    g182(.A(G122), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G116), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n213), .A2(G122), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(G107), .B(new_n368), .C1(new_n372), .C2(KEYINPUT14), .ZN(new_n373));
  XNOR2_X1  g187(.A(G128), .B(G143), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n374), .A2(G134), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n370), .A2(new_n371), .A3(new_n194), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(G134), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n373), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT86), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n370), .A2(new_n371), .A3(new_n194), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n194), .B1(new_n370), .B2(new_n371), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n372), .A2(G107), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n376), .A3(KEYINPUT86), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT13), .B1(new_n261), .B2(G143), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(new_n300), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(new_n374), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n385), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n386), .B1(new_n385), .B2(new_n389), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n367), .B(new_n378), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT88), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n385), .A2(new_n389), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT87), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n385), .A2(new_n389), .A3(new_n386), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n398), .A2(KEYINPUT88), .A3(new_n367), .A4(new_n378), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n378), .B1(new_n390), .B2(new_n391), .ZN(new_n400));
  INV_X1    g214(.A(new_n367), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n394), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G478), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(KEYINPUT15), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n403), .A2(new_n273), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n406), .B1(new_n403), .B2(new_n273), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n365), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n403), .A2(new_n273), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n405), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n403), .A2(new_n273), .A3(new_n406), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(KEYINPUT89), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G113), .B(G122), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(new_n191), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n258), .A2(KEYINPUT16), .A3(G140), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G140), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G125), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n258), .A2(G140), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT16), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n422), .A3(G146), .ZN(new_n423));
  NOR2_X1   g237(.A1(G237), .A2(G953), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(G143), .A3(G214), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(G143), .B1(new_n424), .B2(G214), .ZN(new_n427));
  OAI21_X1  g241(.A(G131), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G237), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n269), .A3(G214), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n252), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n307), .A3(new_n425), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G125), .B(G140), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n434), .B(KEYINPUT19), .Z(new_n435));
  OAI211_X1 g249(.A(new_n423), .B(new_n433), .C1(new_n435), .C2(G146), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n425), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT18), .A3(G131), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n434), .B(new_n255), .ZN(new_n439));
  NAND2_X1  g253(.A1(KEYINPUT18), .A2(G131), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n431), .A2(new_n425), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n416), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n442), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT17), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n428), .A2(new_n445), .A3(new_n432), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n437), .A2(KEYINPUT17), .A3(G131), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n418), .A2(new_n422), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(KEYINPUT77), .A3(new_n255), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n417), .B1(new_n434), .B2(KEYINPUT16), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n451), .B1(new_n452), .B2(G146), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT76), .B1(new_n452), .B2(G146), .ZN(new_n454));
  AND4_X1   g268(.A1(KEYINPUT76), .A2(new_n418), .A3(new_n422), .A4(G146), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n450), .B(new_n453), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n448), .B1(new_n456), .B2(KEYINPUT85), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT76), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n423), .B(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n450), .A4(new_n453), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n444), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n443), .B1(new_n462), .B2(new_n416), .ZN(new_n463));
  NOR2_X1   g277(.A1(G475), .A2(G902), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT20), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n467));
  INV_X1    g281(.A(new_n416), .ZN(new_n468));
  AOI211_X1 g282(.A(new_n468), .B(new_n444), .C1(new_n457), .C2(new_n461), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n467), .B(new_n464), .C1(new_n469), .C2(new_n443), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n462), .A2(new_n416), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n273), .B1(new_n471), .B2(new_n469), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n466), .A2(new_n470), .B1(new_n472), .B2(G475), .ZN(new_n473));
  INV_X1    g287(.A(G952), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(G953), .ZN(new_n475));
  INV_X1    g289(.A(G234), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n429), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT21), .B(G898), .Z(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT90), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n273), .B(new_n269), .C1(G234), .C2(G237), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n473), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT91), .B1(new_n414), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n466), .A2(new_n470), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n472), .A2(G475), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n487), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n489), .A2(new_n490), .A3(new_n413), .A4(new_n409), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n364), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT22), .B(G137), .ZN(new_n494));
  NOR3_X1   g308(.A1(new_n357), .A2(new_n476), .A3(G953), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n494), .B(new_n495), .Z(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n434), .A2(new_n255), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n423), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G128), .B1(new_n211), .B2(new_n212), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n215), .A2(new_n261), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT24), .B(G110), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(KEYINPUT75), .ZN(new_n503));
  INV_X1    g317(.A(G110), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n504), .A2(KEYINPUT24), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(KEYINPUT24), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT75), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n500), .B(new_n501), .C1(new_n503), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n500), .A2(KEYINPUT23), .A3(new_n501), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n261), .B1(new_n211), .B2(new_n212), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT23), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n504), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT78), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT78), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n509), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n499), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n504), .B1(new_n510), .B2(new_n513), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n503), .A2(new_n508), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n500), .A2(new_n501), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n456), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n497), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n509), .A2(new_n517), .A3(new_n514), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n517), .B1(new_n509), .B2(new_n514), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n423), .B(new_n498), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n524), .A3(new_n496), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n366), .B1(G234), .B2(new_n273), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n532), .A2(G902), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n526), .A2(new_n530), .A3(new_n273), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT25), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n526), .A2(new_n530), .A3(KEYINPUT25), .A4(new_n273), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n535), .B1(new_n540), .B2(new_n532), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n424), .A2(G210), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT27), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT26), .B(G101), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n300), .A2(G137), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n302), .A2(G134), .ZN(new_n550));
  OAI21_X1  g364(.A(G131), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n257), .A2(new_n308), .A3(new_n551), .A4(new_n262), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT71), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n320), .B1(new_n309), .B2(new_n310), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n247), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n267), .A2(KEYINPUT64), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT64), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n264), .B(new_n558), .C1(new_n265), .C2(new_n266), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n327), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n308), .A2(new_n551), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT65), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n308), .A2(new_n551), .A3(KEYINPUT65), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n322), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n229), .A2(new_n235), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n548), .B1(new_n556), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n247), .A2(new_n552), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT28), .B1(new_n570), .B2(new_n555), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n547), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT30), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n554), .B2(new_n555), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n560), .A2(new_n565), .A3(new_n573), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n567), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n578));
  NAND4_X1  g392(.A1(new_n577), .A2(new_n556), .A3(new_n546), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n267), .B1(new_n329), .B2(new_n330), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n308), .A2(new_n551), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n322), .A2(new_n581), .A3(new_n553), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n552), .A2(KEYINPUT71), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT30), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n247), .B1(new_n585), .B2(new_n575), .ZN(new_n586));
  INV_X1    g400(.A(new_n556), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n586), .A2(new_n587), .A3(new_n547), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT31), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n572), .B(new_n579), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(G472), .A2(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT32), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT32), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n594), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n556), .A2(KEYINPUT73), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT73), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n554), .A2(new_n555), .A3(new_n598), .A4(new_n247), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n567), .B1(new_n580), .B2(new_n584), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT28), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n571), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT29), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n547), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT74), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n547), .B1(new_n586), .B2(new_n587), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n569), .A2(new_n571), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n604), .B(new_n609), .C1(new_n610), .C2(new_n547), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n556), .A2(KEYINPUT73), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n600), .A3(new_n599), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n571), .B1(new_n613), .B2(KEYINPUT28), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(KEYINPUT74), .A3(new_n605), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n608), .A2(new_n611), .A3(new_n615), .A4(new_n273), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(G472), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n542), .B1(new_n596), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n493), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(new_n199), .ZN(G3));
  INV_X1    g435(.A(KEYINPUT92), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n590), .A2(new_n273), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n592), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n356), .A2(new_n541), .A3(new_n362), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n622), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n623), .A2(G472), .B1(new_n591), .B2(new_n590), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n354), .A2(KEYINPUT81), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n344), .A2(new_n347), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n630), .A2(new_n342), .A3(new_n349), .A4(new_n273), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n361), .B1(new_n632), .B2(new_n341), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n628), .A2(KEYINPUT92), .A3(new_n541), .A4(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n627), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n410), .A2(new_n404), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n403), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n402), .A2(KEYINPUT33), .A3(new_n392), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n404), .A2(G902), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n636), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n487), .A2(new_n488), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n292), .A2(KEYINPUT93), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT93), .ZN(new_n648));
  AOI211_X1 g462(.A(new_n648), .B(new_n188), .C1(new_n290), .C2(new_n291), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n484), .B(new_n646), .C1(new_n647), .C2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n635), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  AOI21_X1  g468(.A(new_n644), .B1(new_n413), .B2(new_n409), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n484), .B(new_n655), .C1(new_n647), .C2(new_n649), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT94), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n248), .A2(new_n285), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(KEYINPUT82), .B2(new_n276), .ZN(new_n659));
  AOI21_X1  g473(.A(G902), .B1(new_n659), .B2(new_n279), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n288), .B1(new_n660), .B2(new_n272), .ZN(new_n661));
  INV_X1    g475(.A(new_n291), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n187), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n648), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n292), .A2(KEYINPUT93), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT94), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n484), .A4(new_n655), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n657), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n635), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NAND2_X1  g486(.A1(new_n529), .A2(new_n524), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n497), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  AOI22_X1  g489(.A1(new_n540), .A2(new_n532), .B1(new_n533), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n625), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n364), .A2(new_n492), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  AOI21_X1  g494(.A(new_n676), .B1(new_n596), .B2(new_n617), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n478), .B1(new_n482), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n414), .A2(new_n473), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n681), .A2(new_n666), .A3(new_n633), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  NAND2_X1  g501(.A1(new_n290), .A2(new_n291), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT38), .Z(new_n689));
  NAND2_X1  g503(.A1(new_n540), .A2(new_n532), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n675), .A2(new_n533), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n414), .A2(new_n644), .ZN(new_n693));
  NOR4_X1   g507(.A1(new_n689), .A2(new_n188), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n683), .B(KEYINPUT39), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n633), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n696), .B(KEYINPUT40), .Z(new_n697));
  NOR2_X1   g511(.A1(new_n586), .A2(new_n587), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n547), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n273), .B1(new_n613), .B2(new_n546), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n596), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n694), .A2(new_n697), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  NAND3_X1  g518(.A1(new_n643), .A2(new_n644), .A3(new_n684), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n681), .A2(new_n666), .A3(new_n633), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT95), .ZN(new_n708));
  AOI211_X1 g522(.A(new_n676), .B(new_n363), .C1(new_n596), .C2(new_n617), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT95), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n710), .A3(new_n666), .A4(new_n706), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  INV_X1    g527(.A(KEYINPUT96), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n349), .B1(new_n348), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n714), .B2(new_n348), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n632), .A3(new_n362), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n542), .B(new_n717), .C1(new_n596), .C2(new_n617), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT97), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n651), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n717), .ZN(new_n721));
  INV_X1    g535(.A(new_n617), .ZN(new_n722));
  INV_X1    g536(.A(new_n595), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n594), .B1(new_n590), .B2(new_n591), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n721), .B(new_n541), .C1(new_n722), .C2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT97), .B1(new_n726), .B2(new_n650), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n720), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT98), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n728), .B(new_n730), .ZN(G15));
  NAND2_X1  g545(.A1(new_n669), .A2(new_n718), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  AOI21_X1  g547(.A(new_n717), .B1(new_n664), .B2(new_n665), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n492), .A3(new_n681), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT99), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n734), .A2(new_n492), .A3(new_n681), .A4(KEYINPUT99), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  INV_X1    g554(.A(new_n693), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n666), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n591), .ZN(new_n743));
  INV_X1    g557(.A(new_n579), .ZN(new_n744));
  INV_X1    g558(.A(new_n588), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n744), .B1(new_n745), .B2(KEYINPUT31), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n614), .A2(new_n546), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(G472), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n749), .B1(new_n590), .B2(new_n273), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n721), .A3(new_n541), .A4(new_n484), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n742), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n369), .ZN(G24));
  NOR4_X1   g568(.A1(new_n705), .A2(new_n748), .A3(new_n750), .A4(new_n676), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n734), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  NAND2_X1  g571(.A1(G469), .A2(G902), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT100), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n340), .B2(G469), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n350), .B2(new_n355), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(KEYINPUT101), .A3(new_n362), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT101), .ZN(new_n763));
  INV_X1    g577(.A(new_n759), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n339), .B2(new_n349), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n629), .B2(new_n631), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n763), .B1(new_n766), .B2(new_n361), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n290), .A2(new_n187), .A3(new_n291), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n762), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n618), .A3(new_n706), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n770), .A2(new_n618), .A3(KEYINPUT42), .A4(new_n706), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  NAND3_X1  g590(.A1(new_n770), .A2(new_n618), .A3(new_n685), .ZN(new_n777));
  XOR2_X1   g591(.A(KEYINPUT102), .B(G134), .Z(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(G36));
  NAND2_X1  g593(.A1(new_n643), .A2(new_n473), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT103), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT43), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n625), .A3(new_n692), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT44), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n340), .A2(KEYINPUT45), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n340), .A2(KEYINPUT45), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(G469), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT46), .B1(new_n790), .B2(new_n764), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(new_n631), .B2(new_n629), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(KEYINPUT46), .A3(new_n764), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n361), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n695), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n768), .B(KEYINPUT104), .Z(new_n796));
  NOR4_X1   g610(.A1(new_n786), .A2(new_n787), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n302), .ZN(G39));
  XNOR2_X1  g612(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n794), .B(new_n799), .Z(new_n800));
  NAND3_X1  g614(.A1(new_n706), .A2(new_n542), .A3(new_n769), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n801), .A2(new_n725), .A3(new_n722), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  NAND2_X1  g618(.A1(new_n686), .A2(new_n756), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n692), .A2(new_n683), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n766), .A2(new_n361), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n807), .A2(KEYINPUT109), .A3(new_n808), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(new_n666), .A3(new_n702), .A4(new_n741), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n712), .A2(new_n806), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT52), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n805), .B1(new_n711), .B2(new_n708), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n818), .A3(new_n814), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n753), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n728), .A2(new_n739), .A3(new_n732), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n755), .A2(new_n770), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n407), .A2(new_n408), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n473), .A2(new_n825), .A3(new_n684), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n768), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n681), .A2(new_n633), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n777), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n775), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n293), .A2(new_n295), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT107), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n644), .A2(new_n825), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n831), .A2(new_n832), .A3(new_n484), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n663), .A2(new_n294), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n292), .A2(KEYINPUT84), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n484), .A3(new_n836), .A4(new_n833), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT107), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n635), .A2(new_n834), .A3(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n293), .A2(new_n295), .A3(new_n483), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n645), .B(KEYINPUT106), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n841), .A3(new_n627), .A4(new_n634), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n364), .B(new_n492), .C1(new_n618), .C2(new_n677), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n830), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT108), .B1(new_n823), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n739), .A2(new_n728), .A3(new_n732), .A4(new_n822), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n843), .A2(new_n842), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n775), .A3(new_n839), .A4(new_n829), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT108), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n821), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(KEYINPUT110), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT110), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n823), .A2(new_n845), .A3(KEYINPUT108), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n850), .B1(new_n847), .B2(new_n849), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n820), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n855), .B1(new_n858), .B2(KEYINPUT53), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n847), .A2(new_n849), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n853), .B1(new_n805), .B2(KEYINPUT52), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n821), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n854), .A2(new_n859), .A3(new_n860), .A4(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n858), .A2(KEYINPUT53), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT53), .B1(new_n805), .B2(KEYINPUT52), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n866), .B(new_n820), .C1(new_n857), .C2(new_n856), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT54), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT111), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT111), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n864), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n783), .A2(new_n478), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n717), .A2(new_n768), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n619), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT48), .ZN(new_n877));
  INV_X1    g691(.A(new_n702), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n541), .A3(new_n478), .A4(new_n874), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n783), .A2(new_n541), .A3(new_n478), .A4(new_n751), .ZN(new_n880));
  INV_X1    g694(.A(new_n734), .ZN(new_n881));
  OAI221_X1 g695(.A(new_n475), .B1(new_n645), .B2(new_n879), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT112), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n689), .A2(new_n188), .A3(new_n721), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n884), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT50), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n880), .A2(new_n796), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n716), .A2(new_n632), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n362), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n800), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n879), .A2(new_n644), .A3(new_n643), .ZN(new_n895));
  INV_X1    g709(.A(new_n875), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n748), .A2(new_n676), .A3(new_n750), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n894), .A2(KEYINPUT51), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n883), .B1(new_n890), .B2(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n888), .A2(KEYINPUT113), .A3(new_n889), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT113), .B1(new_n888), .B2(new_n889), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT114), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT114), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n905), .B(new_n898), .C1(new_n901), .C2(new_n902), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n906), .A3(new_n894), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT51), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n900), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n870), .A2(new_n872), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT115), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT115), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n870), .A2(new_n912), .A3(new_n872), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n474), .A2(new_n269), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n892), .B(KEYINPUT49), .Z(new_n916));
  NOR4_X1   g730(.A1(new_n542), .A2(new_n780), .A3(new_n361), .A4(new_n188), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n878), .A3(new_n689), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(G75));
  NOR2_X1   g733(.A1(new_n269), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n863), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n852), .A2(new_n853), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n855), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n273), .B1(new_n923), .B2(new_n854), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(G210), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT56), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n249), .A2(new_n251), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT116), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT117), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT55), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n271), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n920), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n925), .A2(KEYINPUT118), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT118), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n924), .A2(new_n935), .A3(G210), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n932), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n934), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n933), .A2(new_n939), .ZN(G51));
  XNOR2_X1  g754(.A(new_n759), .B(KEYINPUT57), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n860), .B1(new_n923), .B2(new_n854), .ZN(new_n942));
  INV_X1    g756(.A(new_n864), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n630), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n924), .A2(G469), .A3(new_n789), .A4(new_n788), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n920), .B1(new_n945), .B2(new_n946), .ZN(G54));
  NAND3_X1  g761(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n948), .A2(new_n463), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n463), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n920), .ZN(G60));
  INV_X1    g765(.A(new_n640), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT59), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n952), .B(new_n954), .C1(new_n942), .C2(new_n943), .ZN(new_n955));
  INV_X1    g769(.A(new_n920), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n870), .A2(new_n872), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n954), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n957), .B1(new_n640), .B2(new_n959), .ZN(G63));
  NAND2_X1  g774(.A1(new_n923), .A2(new_n854), .ZN(new_n961));
  XNOR2_X1  g775(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n366), .A2(new_n273), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n531), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n961), .A2(new_n675), .A3(new_n964), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n956), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(G66));
  INV_X1    g784(.A(G224), .ZN(new_n971));
  OAI21_X1  g785(.A(G953), .B1(new_n481), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n847), .A2(new_n844), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n973), .B2(G953), .ZN(new_n974));
  INV_X1    g788(.A(new_n929), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(G898), .B2(new_n269), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n974), .B(new_n976), .ZN(G69));
  NOR2_X1   g791(.A1(new_n696), .A2(new_n768), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n618), .B(new_n978), .C1(new_n841), .C2(new_n833), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT122), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n797), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n982), .A2(KEYINPUT123), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(KEYINPUT123), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n817), .A2(new_n703), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n986), .A2(KEYINPUT62), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT121), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(KEYINPUT62), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n985), .A2(new_n803), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n269), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n585), .A2(new_n575), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(new_n435), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n803), .A2(new_n777), .ZN(new_n994));
  INV_X1    g808(.A(new_n775), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n795), .A2(new_n619), .A3(new_n742), .ZN(new_n996));
  NOR4_X1   g810(.A1(new_n994), .A2(new_n797), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n997), .A2(new_n269), .A3(new_n817), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n993), .B1(G900), .B2(G953), .ZN(new_n999));
  AOI22_X1  g813(.A1(new_n991), .A2(new_n993), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n998), .A2(new_n999), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(KEYINPUT124), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1000), .B(new_n1003), .ZN(G72));
  INV_X1    g818(.A(new_n699), .ZN(new_n1005));
  OR3_X1    g819(.A1(new_n990), .A2(new_n847), .A3(new_n844), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT125), .Z(new_n1009));
  AOI21_X1  g823(.A(new_n1005), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n997), .A2(new_n817), .A3(new_n973), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n1009), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n547), .B(new_n698), .C1(new_n1012), .C2(KEYINPUT126), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n1012), .A2(KEYINPUT126), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n956), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n865), .A2(new_n867), .ZN(new_n1017));
  AOI211_X1 g831(.A(new_n1016), .B(new_n1017), .C1(new_n547), .C2(new_n698), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n1010), .A2(new_n1015), .A3(new_n1018), .ZN(G57));
endmodule


