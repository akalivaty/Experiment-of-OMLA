//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n187));
  INV_X1    g001(.A(G107), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G104), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G107), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G101), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n192), .A2(KEYINPUT85), .A3(new_n193), .A4(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n194), .A2(new_n189), .A3(new_n193), .A4(new_n191), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT85), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT4), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n189), .A3(new_n191), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G101), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G143), .B(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n209), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n201), .A2(new_n200), .A3(G101), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n190), .A2(G107), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n188), .A2(G104), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n218), .B(G101), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G104), .B(G107), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT86), .B1(new_n222), .B2(new_n193), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n195), .A2(new_n198), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT10), .ZN(new_n225));
  AOI21_X1  g039(.A(G128), .B1(new_n205), .B2(new_n207), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n205), .A2(new_n207), .A3(G128), .ZN(new_n227));
  AND2_X1   g041(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g042(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n226), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n206), .B(G146), .C1(new_n228), .C2(new_n229), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n225), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n203), .A2(new_n217), .B1(new_n224), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n235));
  INV_X1    g049(.A(G134), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G137), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT11), .A3(G134), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(G137), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G131), .ZN(new_n242));
  INV_X1    g056(.A(G131), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n237), .A2(new_n239), .A3(new_n243), .A4(new_n240), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n230), .A2(new_n213), .A3(G128), .ZN(new_n247));
  INV_X1    g061(.A(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n208), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n206), .A2(KEYINPUT1), .A3(G146), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n223), .A2(new_n221), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n196), .A2(new_n197), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n196), .A2(new_n197), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n255), .A2(KEYINPUT87), .A3(new_n225), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT87), .B1(new_n255), .B2(new_n225), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n234), .B(new_n246), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n247), .A2(new_n232), .A3(new_n249), .ZN(new_n259));
  OR2_X1    g073(.A1(new_n224), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n246), .B1(new_n260), .B2(new_n255), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n261), .A2(KEYINPUT12), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(KEYINPUT12), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(G110), .B(G140), .ZN(new_n265));
  INV_X1    g079(.A(G953), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n266), .A2(G227), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n265), .B(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n258), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(new_n268), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n234), .B1(new_n256), .B2(new_n257), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n245), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n264), .A2(new_n268), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G469), .B1(new_n273), .B2(G902), .ZN(new_n274));
  INV_X1    g088(.A(G469), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n255), .A2(new_n225), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT87), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n255), .A2(KEYINPUT87), .A3(new_n225), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n246), .B1(new_n281), .B2(new_n234), .ZN(new_n282));
  OAI211_X1 g096(.A(KEYINPUT88), .B(new_n268), .C1(new_n282), .C2(new_n269), .ZN(new_n283));
  INV_X1    g097(.A(new_n268), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n284), .B(new_n258), .C1(new_n262), .C2(new_n263), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n272), .A2(new_n258), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT88), .B1(new_n287), .B2(new_n268), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n275), .B(new_n276), .C1(new_n286), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n274), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT9), .B(G234), .ZN(new_n291));
  OAI21_X1  g105(.A(G221), .B1(new_n291), .B2(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT17), .ZN(new_n294));
  OR2_X1    g108(.A1(KEYINPUT69), .A2(G237), .ZN(new_n295));
  NAND2_X1  g109(.A1(KEYINPUT69), .A2(G237), .ZN(new_n296));
  AOI21_X1  g110(.A(G953), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(G143), .A3(G214), .ZN(new_n298));
  AND2_X1   g112(.A1(KEYINPUT69), .A2(G237), .ZN(new_n299));
  NOR2_X1   g113(.A1(KEYINPUT69), .A2(G237), .ZN(new_n300));
  OAI211_X1 g114(.A(G214), .B(new_n266), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n206), .ZN(new_n302));
  AOI211_X1 g116(.A(new_n294), .B(new_n243), .C1(new_n298), .C2(new_n302), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n298), .A2(new_n243), .A3(new_n302), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n243), .B1(new_n298), .B2(new_n302), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n303), .B1(new_n306), .B2(new_n294), .ZN(new_n307));
  OR2_X1    g121(.A1(KEYINPUT76), .A2(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(KEYINPUT76), .A2(G140), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(G125), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT77), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT77), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G125), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n314), .A3(G140), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(new_n315), .A3(KEYINPUT16), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT78), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n310), .A2(new_n315), .A3(new_n318), .A4(KEYINPUT16), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n312), .A2(new_n314), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(G146), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT79), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n320), .A2(new_n324), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n204), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n320), .A2(new_n329), .A3(G146), .A4(new_n324), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n307), .A2(new_n326), .A3(new_n328), .A4(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G113), .B(G122), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(new_n190), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n301), .B(G143), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT18), .A2(G131), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT94), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n298), .A2(new_n302), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT18), .A4(G131), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n335), .B(KEYINPUT95), .Z(new_n340));
  NAND2_X1  g154(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n310), .A2(new_n315), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G146), .ZN(new_n343));
  INV_X1    g157(.A(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G125), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n311), .A2(G140), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n345), .B2(new_n346), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n204), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n336), .A2(new_n339), .A3(new_n341), .A4(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n331), .A2(new_n333), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT19), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n348), .B2(new_n349), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT96), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n342), .A2(KEYINPUT19), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT96), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n358), .B(new_n354), .C1(new_n348), .C2(new_n349), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n356), .A2(new_n204), .A3(new_n357), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n337), .A2(G131), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n298), .A2(new_n302), .A3(new_n243), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n325), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n352), .ZN(new_n365));
  INV_X1    g179(.A(new_n333), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT97), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT97), .ZN(new_n368));
  AOI211_X1 g182(.A(new_n368), .B(new_n333), .C1(new_n364), .C2(new_n352), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n353), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G475), .A2(G902), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT98), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(KEYINPUT98), .A3(new_n371), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(KEYINPUT20), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT98), .B1(new_n370), .B2(new_n371), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n378));
  INV_X1    g192(.A(new_n353), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n333), .B1(new_n331), .B2(new_n352), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n276), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n377), .A2(new_n378), .B1(G475), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G210), .B1(G237), .B2(G902), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(G110), .B(G122), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT90), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT2), .B(G113), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G116), .B(G119), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n389), .A2(KEYINPUT67), .A3(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(G116), .B(G119), .Z(new_n392));
  INV_X1    g206(.A(KEYINPUT67), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n216), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n199), .B2(new_n202), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n390), .A2(KEYINPUT5), .ZN(new_n397));
  INV_X1    g211(.A(G116), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n398), .A2(KEYINPUT5), .A3(G119), .ZN(new_n399));
  INV_X1    g213(.A(G113), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n397), .A2(new_n401), .B1(new_n389), .B2(new_n390), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n402), .B(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n387), .B1(new_n396), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n387), .ZN(new_n406));
  INV_X1    g220(.A(new_n202), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(new_n198), .B2(new_n195), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n403), .B(new_n406), .C1(new_n408), .C2(new_n395), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(KEYINPUT6), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n411), .B(new_n387), .C1(new_n396), .C2(new_n404), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n212), .A2(new_n214), .A3(new_n321), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT91), .B(new_n413), .C1(new_n259), .C2(new_n321), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT91), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n231), .A2(new_n415), .A3(new_n232), .A4(new_n322), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G224), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(G953), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n417), .B(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n410), .A2(new_n412), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT93), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n414), .B(new_n416), .C1(new_n424), .C2(new_n419), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n409), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT92), .B(KEYINPUT8), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n387), .B(new_n429), .Z(new_n430));
  NOR2_X1   g244(.A1(new_n224), .A2(new_n402), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n432), .B2(new_n403), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n423), .B(new_n276), .C1(new_n428), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n422), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n387), .B(new_n429), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n431), .B2(new_n404), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n437), .A2(new_n409), .A3(new_n426), .A4(new_n427), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n423), .B1(new_n438), .B2(new_n276), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n385), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n276), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT93), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n442), .A2(new_n384), .A3(new_n422), .A4(new_n434), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G214), .B1(G237), .B2(G902), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n445), .B(KEYINPUT89), .Z(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(G234), .A2(G237), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(G952), .A3(new_n266), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT100), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n448), .A2(G902), .A3(G953), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(G898), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n444), .A2(new_n447), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT15), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n457), .A2(KEYINPUT99), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(KEYINPUT99), .ZN(new_n459));
  OAI21_X1  g273(.A(G478), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n206), .A2(G128), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n248), .A2(G143), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n236), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n398), .A2(KEYINPUT14), .A3(G122), .ZN(new_n465));
  XNOR2_X1  g279(.A(G116), .B(G122), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(G107), .B(new_n465), .C1(new_n467), .C2(KEYINPUT14), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n464), .B(new_n468), .C1(G107), .C2(new_n467), .ZN(new_n469));
  INV_X1    g283(.A(new_n461), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n470), .A2(KEYINPUT13), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n462), .B1(new_n470), .B2(KEYINPUT13), .ZN(new_n472));
  OAI21_X1  g286(.A(G134), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n463), .A2(new_n236), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n466), .B(new_n188), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G217), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n291), .A2(new_n477), .A3(G953), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n469), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n478), .B1(new_n469), .B2(new_n476), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n460), .B1(new_n481), .B2(new_n276), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n276), .B(new_n460), .C1(new_n479), .C2(new_n480), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NOR4_X1   g300(.A1(new_n293), .A2(new_n383), .A3(new_n456), .A4(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT26), .B(G101), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n297), .A2(G210), .ZN(new_n490));
  XOR2_X1   g304(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n490), .A2(new_n491), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n494), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n488), .A3(new_n492), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n238), .A2(KEYINPUT65), .A3(G134), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n236), .B2(G137), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n238), .A2(G134), .ZN(new_n504));
  OAI211_X1 g318(.A(G131), .B(new_n501), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n259), .A2(new_n244), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n245), .A2(new_n215), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n391), .A2(new_n394), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n500), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n512), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n514), .A2(KEYINPUT28), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n499), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  XOR2_X1   g330(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n505), .A2(new_n244), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n231), .B2(new_n232), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n242), .A2(new_n244), .B1(new_n212), .B2(new_n214), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT30), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n510), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT68), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT68), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n522), .A2(new_n523), .A3(new_n526), .A4(new_n510), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n498), .A2(new_n512), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n516), .B1(new_n531), .B2(KEYINPUT31), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT71), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n528), .B2(new_n530), .ZN(new_n534));
  AOI211_X1 g348(.A(KEYINPUT71), .B(new_n529), .C1(new_n525), .C2(new_n527), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n532), .B1(new_n536), .B2(KEYINPUT31), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT72), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT31), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n534), .A2(new_n535), .A3(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n542), .B(new_n538), .C1(new_n544), .C2(new_n532), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n513), .A2(new_n515), .A3(new_n499), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(KEYINPUT29), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n514), .B1(new_n525), .B2(new_n527), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n548), .B(KEYINPUT73), .C1(new_n549), .C2(new_n498), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT73), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n549), .A2(new_n498), .ZN(new_n552));
  INV_X1    g366(.A(new_n515), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n511), .A2(new_n512), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT28), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n555), .A3(new_n498), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT29), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n551), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(G902), .B1(new_n547), .B2(KEYINPUT29), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n550), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n529), .B1(new_n525), .B2(new_n527), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n533), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(KEYINPUT31), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n516), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n543), .B2(new_n563), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n539), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g382(.A1(G472), .A2(new_n561), .B1(new_n568), .B2(KEYINPUT32), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n546), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n477), .B1(G234), .B2(new_n276), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G902), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G119), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G128), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n575), .A2(KEYINPUT74), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(KEYINPUT74), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n576), .B(new_n577), .C1(new_n574), .C2(G128), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT24), .B(G110), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n248), .A2(KEYINPUT23), .A3(G119), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n574), .A2(G128), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n575), .B(new_n581), .C1(new_n582), .C2(KEYINPUT23), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n583), .A2(KEYINPUT75), .ZN(new_n584));
  INV_X1    g398(.A(G110), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n583), .B2(KEYINPUT75), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n580), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n323), .B1(new_n317), .B2(new_n319), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n330), .B1(G146), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n329), .B1(new_n588), .B2(G146), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n578), .A2(new_n579), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(G110), .B2(new_n583), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n325), .A2(new_n350), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT81), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT22), .B(G137), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT82), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n595), .A2(KEYINPUT83), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT83), .ZN(new_n602));
  INV_X1    g416(.A(new_n594), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n326), .A2(new_n328), .A3(new_n330), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n603), .B1(new_n604), .B2(new_n587), .ZN(new_n605));
  INV_X1    g419(.A(new_n600), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n599), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n601), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT84), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n606), .B1(new_n591), .B2(new_n594), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n612), .A2(KEYINPUT83), .B1(new_n605), .B2(new_n599), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n607), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT84), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n573), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n571), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n601), .A2(new_n607), .A3(new_n276), .A4(new_n608), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT25), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n613), .A2(KEYINPUT25), .A3(new_n276), .A4(new_n607), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n487), .A2(new_n570), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  OAI21_X1  g439(.A(G472), .B1(new_n537), .B2(G902), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT101), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n628), .B(G472), .C1(new_n537), .C2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n540), .A2(new_n545), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(G478), .A2(G902), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n481), .A2(new_n276), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n633), .B1(new_n634), .B2(G478), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT102), .B1(new_n469), .B2(new_n476), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n481), .B(new_n638), .Z(new_n639));
  AOI21_X1  g453(.A(new_n635), .B1(new_n639), .B2(G478), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n383), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n445), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n444), .A2(new_n455), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n609), .A2(new_n610), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n614), .A2(KEYINPUT84), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n572), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n292), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n274), .B2(new_n289), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n620), .A2(new_n621), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n571), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n647), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n632), .A2(new_n644), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT103), .Z(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  NOR4_X1   g470(.A1(new_n383), .A2(new_n643), .A3(new_n642), .A4(new_n485), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n632), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NOR2_X1   g474(.A1(new_n600), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n595), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n572), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n651), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n632), .A2(new_n487), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT104), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n665), .B(new_n667), .ZN(G12));
  INV_X1    g482(.A(new_n663), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n650), .B2(new_n571), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n546), .B2(new_n569), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n642), .B1(new_n440), .B2(new_n443), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n649), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(G900), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n451), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n450), .A2(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n383), .A2(new_n485), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  INV_X1    g494(.A(new_n536), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n498), .B1(new_n511), .B2(new_n512), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n276), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n683), .A2(G472), .B1(new_n568), .B2(KEYINPUT32), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n664), .B1(new_n546), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n444), .B(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n376), .A2(new_n382), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n689), .A2(new_n642), .A3(new_n485), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n685), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n677), .B(KEYINPUT39), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n649), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT40), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G143), .ZN(G45));
  INV_X1    g512(.A(new_n677), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n383), .A2(new_n640), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n674), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  OAI21_X1  g517(.A(new_n276), .B1(new_n286), .B2(new_n288), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n705), .A2(new_n292), .A3(new_n289), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n644), .A2(new_n570), .A3(new_n623), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND4_X1  g523(.A1(new_n657), .A2(new_n570), .A3(new_n623), .A4(new_n706), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NOR3_X1   g525(.A1(new_n383), .A2(new_n454), .A3(new_n486), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n705), .A2(new_n292), .A3(new_n289), .A4(new_n672), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n713), .A2(KEYINPUT107), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(KEYINPUT107), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n671), .B(new_n712), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  AOI211_X1 g531(.A(new_n642), .B(new_n485), .C1(new_n440), .C2(new_n443), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n383), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT108), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n383), .A2(new_n721), .A3(new_n718), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n568), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n626), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n616), .A3(new_n622), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n292), .A2(new_n705), .A3(new_n289), .A4(new_n455), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  OAI211_X1 g543(.A(new_n626), .B(new_n724), .C1(new_n622), .C2(new_n669), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n700), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n714), .B2(new_n715), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  OAI211_X1 g547(.A(KEYINPUT32), .B(new_n538), .C1(new_n544), .C2(new_n532), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT110), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n568), .A2(KEYINPUT32), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n568), .A2(KEYINPUT110), .A3(KEYINPUT32), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT111), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n568), .B2(KEYINPUT32), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(KEYINPUT32), .B2(new_n568), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n743));
  INV_X1    g557(.A(new_n738), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n561), .A2(G472), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n739), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  OR3_X1    g561(.A1(new_n444), .A2(KEYINPUT109), .A3(new_n642), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT109), .B1(new_n444), .B2(new_n642), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  NOR4_X1   g565(.A1(new_n750), .A2(new_n700), .A3(new_n293), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n747), .A2(new_n752), .A3(new_n623), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n748), .A2(new_n649), .A3(new_n749), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n570), .A3(new_n623), .A4(new_n701), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n751), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT112), .B(G131), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G33));
  NAND4_X1  g573(.A1(new_n754), .A2(new_n570), .A3(new_n623), .A4(new_n678), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  NAND2_X1  g575(.A1(new_n689), .A2(new_n640), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT43), .Z(new_n763));
  NOR2_X1   g577(.A1(new_n632), .A2(new_n670), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n764), .A3(KEYINPUT44), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n273), .A2(KEYINPUT45), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n273), .A2(KEYINPUT45), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(G469), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(G469), .A2(G902), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT46), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n289), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n772), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n648), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(new_n692), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n750), .B(KEYINPUT113), .Z(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n767), .A2(new_n768), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  XNOR2_X1  g596(.A(new_n777), .B(KEYINPUT47), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n570), .A2(new_n750), .A3(new_n623), .A4(new_n700), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  NOR4_X1   g600(.A1(new_n688), .A2(new_n762), .A3(new_n648), .A4(new_n446), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n546), .A2(new_n684), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n705), .A2(new_n289), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT49), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n787), .A2(new_n623), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n450), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n706), .A2(new_n748), .A3(new_n749), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n763), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n730), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n616), .A2(new_n622), .A3(new_n450), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n795), .A2(new_n789), .A3(new_n799), .ZN(new_n800));
  OR3_X1    g614(.A1(new_n800), .A2(new_n383), .A3(new_n640), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(KEYINPUT117), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n763), .A2(new_n793), .A3(new_n726), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n445), .B1(KEYINPUT117), .B2(new_n803), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n706), .A2(new_n687), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(new_n805), .A3(new_n808), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n802), .A2(KEYINPUT118), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n798), .A3(new_n801), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n813), .B1(new_n814), .B2(new_n809), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n790), .A2(new_n648), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n780), .B(new_n806), .C1(new_n783), .C2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n812), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n817), .A2(KEYINPUT51), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n823), .A2(new_n809), .A3(new_n814), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n747), .A2(new_n623), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n796), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT48), .Z(new_n827));
  NOR2_X1   g641(.A1(new_n714), .A2(new_n715), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n806), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(G952), .B(new_n266), .C1(new_n800), .C2(new_n641), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n824), .A2(new_n827), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n822), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n485), .B(KEYINPUT114), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n677), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n689), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT115), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n689), .A2(new_n839), .A3(new_n836), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n838), .A2(new_n671), .A3(new_n754), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n731), .A2(new_n754), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n842), .A3(new_n760), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n756), .B2(new_n753), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n376), .A2(new_n835), .A3(new_n382), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n456), .B1(new_n641), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n652), .A3(new_n631), .A4(new_n630), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n716), .A2(new_n728), .A3(new_n847), .A4(new_n710), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n665), .A2(new_n624), .A3(new_n707), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  AOI211_X1 g666(.A(new_n648), .B(new_n677), .C1(new_n274), .C2(new_n289), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n788), .A2(new_n670), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n383), .A2(new_n721), .A3(new_n718), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n721), .B1(new_n383), .B2(new_n718), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n852), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n723), .A2(new_n685), .A3(KEYINPUT116), .A4(new_n853), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n671), .B(new_n673), .C1(new_n678), .C2(new_n701), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n861), .A2(new_n732), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n860), .B2(new_n862), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT53), .B1(new_n851), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n848), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n665), .A2(new_n624), .A3(new_n707), .ZN(new_n869));
  INV_X1    g683(.A(new_n843), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n868), .A2(new_n757), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  NOR4_X1   g686(.A1(new_n871), .A2(new_n864), .A3(new_n865), .A4(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n834), .B1(new_n867), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n865), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n872), .B1(new_n877), .B2(new_n871), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n851), .A2(new_n866), .A3(KEYINPUT53), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT54), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n820), .A2(new_n821), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n833), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n792), .B1(new_n883), .B2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n266), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n276), .B1(new_n878), .B2(new_n879), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT56), .B1(new_n888), .B2(G210), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n410), .A2(new_n412), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n421), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT55), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n887), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n888), .B(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n385), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n893), .B1(new_n896), .B2(new_n898), .ZN(G51));
  XNOR2_X1  g713(.A(new_n888), .B(KEYINPUT120), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(new_n771), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n772), .B(KEYINPUT57), .Z(new_n902));
  NAND2_X1  g716(.A1(new_n881), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n286), .A2(new_n288), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT121), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n886), .B1(new_n901), .B2(new_n906), .ZN(G54));
  INV_X1    g721(.A(new_n370), .ZN(new_n908));
  NAND2_X1  g722(.A1(KEYINPUT58), .A2(G475), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n908), .B1(new_n900), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .A4(new_n370), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n910), .A2(new_n911), .A3(new_n887), .ZN(G60));
  XOR2_X1   g726(.A(new_n633), .B(KEYINPUT59), .Z(new_n913));
  NOR2_X1   g727(.A1(new_n639), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n874), .A2(new_n880), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT122), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n874), .A2(new_n880), .A3(new_n917), .A4(new_n914), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n913), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n874), .A2(new_n880), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n886), .B1(new_n921), .B2(new_n639), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n919), .A2(KEYINPUT123), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(G63));
  NOR2_X1   g741(.A1(new_n867), .A2(new_n873), .ZN(new_n928));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n662), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n611), .A2(new_n615), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n932), .B(new_n887), .C1(new_n933), .C2(new_n931), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT61), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n934), .B(new_n936), .ZN(G66));
  OAI21_X1  g751(.A(G953), .B1(new_n452), .B2(new_n418), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n850), .B2(G953), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n890), .B1(G898), .B2(new_n266), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G69));
  AOI21_X1  g755(.A(new_n266), .B1(G227), .B2(G900), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n781), .A2(new_n862), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT125), .B1(new_n781), .B2(new_n862), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n778), .A2(new_n723), .A3(new_n825), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n785), .A2(new_n757), .A3(new_n760), .A4(new_n948), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n266), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n522), .A2(new_n523), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(G900), .B2(G953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n697), .A2(new_n862), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n570), .A2(new_n623), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n641), .A2(new_n845), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n960), .A2(new_n962), .A3(new_n692), .A4(new_n754), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n781), .A2(new_n785), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n958), .A2(new_n959), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n266), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n954), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n943), .B1(new_n956), .B2(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(G72));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n681), .B2(new_n552), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n887), .B1(new_n928), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n549), .A2(new_n499), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT127), .Z(new_n976));
  NAND2_X1  g790(.A1(new_n950), .A2(new_n850), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n976), .B1(new_n977), .B2(new_n972), .ZN(new_n978));
  INV_X1    g792(.A(new_n850), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n972), .B1(new_n965), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n549), .A2(new_n499), .ZN(new_n981));
  AOI211_X1 g795(.A(new_n974), .B(new_n978), .C1(new_n980), .C2(new_n981), .ZN(G57));
endmodule


