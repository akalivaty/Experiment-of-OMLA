//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT27), .B(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT67), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(KEYINPUT28), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT28), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT26), .ZN(new_n209));
  INV_X1    g008(.A(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT26), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G169gat), .B2(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  OAI221_X1 g013(.A(new_n209), .B1(new_n210), .B2(new_n204), .C1(new_n212), .C2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n206), .A2(new_n207), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT25), .ZN(new_n218));
  INV_X1    g017(.A(G169gat), .ZN(new_n219));
  INV_X1    g018(.A(G176gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(KEYINPUT23), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n204), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(new_n213), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n210), .ZN(new_n226));
  NAND2_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(G190gat), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n229), .B(new_n230), .C1(G169gat), .C2(G176gat), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT66), .B1(new_n208), .B2(KEYINPUT23), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n224), .A2(new_n228), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n218), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n228), .A2(new_n232), .A3(new_n231), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n234), .B(new_n218), .C1(new_n236), .C2(new_n223), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n217), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(G127gat), .A2(G134gat), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT68), .B(G134gat), .Z(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(G127gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(G113gat), .B2(G120gat), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n244), .B1(G113gat), .B2(G120gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n248));
  OAI21_X1  g047(.A(G120gat), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n240), .ZN(new_n250));
  NAND2_X1  g049(.A1(G127gat), .A2(G134gat), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n244), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n242), .A2(new_n246), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n239), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n234), .B1(new_n236), .B2(new_n223), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT25), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n215), .B1(KEYINPUT28), .B2(new_n205), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n256), .A2(new_n237), .B1(new_n257), .B2(new_n206), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n249), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT68), .B(G134gat), .ZN(new_n260));
  INV_X1    g059(.A(G127gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n250), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n259), .B1(new_n262), .B2(new_n245), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n254), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G227gat), .A2(G233gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n267), .B(KEYINPUT64), .Z(new_n268));
  AOI21_X1  g067(.A(new_n202), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G71gat), .B(G99gat), .Z(new_n270));
  XNOR2_X1  g069(.A(G15gat), .B(G43gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT33), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n254), .A2(new_n264), .A3(new_n268), .A4(new_n272), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT70), .B1(new_n276), .B2(new_n273), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n275), .B1(new_n269), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n268), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n265), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n280), .A2(KEYINPUT34), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(KEYINPUT34), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n278), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n281), .A2(new_n282), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n285), .B(new_n275), .C1(new_n269), .C2(new_n277), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G78gat), .B(G106gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT31), .B(G50gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(KEYINPUT79), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G22gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT72), .B(G211gat), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT22), .B1(new_n296), .B2(G218gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n295), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n302));
  OAI21_X1  g101(.A(G218gat), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(new_n294), .A3(new_n298), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT3), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT83), .ZN(new_n310));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT2), .ZN(new_n312));
  INV_X1    g111(.A(G148gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(G141gat), .ZN(new_n314));
  INV_X1    g113(.A(G141gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(G148gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n312), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n315), .A2(G148gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n313), .A2(G141gat), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n323), .A2(new_n324), .B1(KEYINPUT2), .B2(new_n311), .ZN(new_n325));
  OR2_X1    g124(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n326));
  INV_X1    g125(.A(G155gat), .ZN(new_n327));
  INV_X1    g126(.A(G162gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n329), .A3(new_n311), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n322), .A2(new_n331), .ZN(new_n332));
  OR3_X1    g131(.A1(new_n309), .A2(new_n310), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G228gat), .ZN(new_n334));
  INV_X1    g133(.A(G233gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n318), .A2(new_n320), .ZN(new_n337));
  XNOR2_X1  g136(.A(G141gat), .B(G148gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(G155gat), .B2(G162gat), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n337), .B(new_n329), .C1(new_n338), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n330), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n308), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT84), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n307), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n346), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n310), .B1(new_n309), .B2(new_n332), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n333), .A2(new_n336), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n345), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT82), .B1(new_n351), .B2(new_n307), .ZN(new_n352));
  INV_X1    g151(.A(new_n307), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT82), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n345), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n294), .B1(new_n305), .B2(new_n298), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n357), .B2(KEYINPUT80), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n300), .A2(new_n359), .A3(new_n306), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n360), .A3(KEYINPUT81), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n343), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(new_n322), .B2(new_n331), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT76), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n356), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n293), .B(new_n350), .C1(new_n371), .C2(new_n336), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT3), .B1(new_n361), .B2(new_n362), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n369), .B1(new_n374), .B2(new_n364), .ZN(new_n375));
  OAI22_X1  g174(.A1(new_n375), .A2(new_n356), .B1(new_n334), .B2(new_n335), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n293), .B1(new_n376), .B2(new_n350), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n292), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n350), .B1(new_n371), .B2(new_n336), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G22gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n290), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n372), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n287), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n253), .A2(new_n332), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n341), .A2(new_n342), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n263), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n385), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n387), .A2(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n395), .A2(new_n263), .A3(new_n344), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n390), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n263), .B1(new_n367), .B2(new_n368), .ZN(new_n398));
  AND2_X1   g197(.A1(new_n398), .A2(KEYINPUT4), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n392), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n396), .A2(new_n385), .A3(new_n390), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT4), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT76), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT76), .B1(new_n341), .B2(new_n342), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n393), .B(new_n253), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n402), .B1(new_n405), .B2(KEYINPUT77), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(new_n398), .B2(new_n393), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT78), .B(new_n401), .C1(new_n406), .C2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(KEYINPUT77), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n369), .A2(new_n407), .A3(new_n393), .A4(new_n253), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(new_n402), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT78), .B1(new_n413), .B2(new_n401), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n400), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(G1gat), .B(G29gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT0), .ZN(new_n417));
  XNOR2_X1  g216(.A(G57gat), .B(G85gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421));
  INV_X1    g220(.A(new_n419), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n400), .B(new_n422), .C1(new_n410), .C2(new_n414), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n415), .A2(KEYINPUT6), .A3(new_n419), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT74), .ZN(new_n428));
  XNOR2_X1  g227(.A(G64gat), .B(G92gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n428), .B(new_n429), .Z(new_n430));
  INV_X1    g229(.A(G226gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(new_n335), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n239), .B2(new_n308), .ZN(new_n433));
  INV_X1    g232(.A(new_n432), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n258), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT73), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT73), .B1(new_n239), .B2(new_n432), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n307), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n434), .B1(new_n258), .B2(KEYINPUT29), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n239), .A2(new_n432), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n353), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n430), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n433), .A2(new_n435), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n307), .ZN(new_n446));
  INV_X1    g245(.A(new_n430), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n437), .B1(new_n442), .B2(KEYINPUT73), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n446), .B(new_n447), .C1(new_n448), .C2(new_n307), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n444), .A2(KEYINPUT30), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n439), .A2(new_n443), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT30), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n447), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n426), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT35), .ZN(new_n456));
  OR3_X1    g255(.A1(new_n384), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n456), .B1(new_n384), .B2(new_n455), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n378), .A2(new_n460), .A3(new_n382), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n378), .B2(new_n382), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n455), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OR2_X1    g262(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n287), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n284), .A2(new_n286), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n463), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n469), .B1(new_n463), .B2(new_n468), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n450), .A2(new_n453), .ZN(new_n474));
  INV_X1    g273(.A(new_n420), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n396), .B1(new_n406), .B2(new_n408), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n391), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n477), .B(KEYINPUT39), .C1(new_n391), .C2(new_n389), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT39), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n479), .A3(new_n391), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n480), .A2(new_n481), .A3(new_n422), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n481), .B1(new_n480), .B2(new_n422), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n478), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT40), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n475), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(KEYINPUT40), .B(new_n478), .C1(new_n482), .C2(new_n483), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n480), .A2(new_n422), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT87), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n480), .A2(new_n481), .A3(new_n422), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(KEYINPUT88), .A3(KEYINPUT40), .A4(new_n478), .ZN(new_n494));
  AND4_X1   g293(.A1(new_n474), .A2(new_n486), .A3(new_n489), .A4(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT37), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n446), .B(new_n496), .C1(new_n448), .C2(new_n307), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n496), .B1(new_n445), .B2(new_n353), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(new_n448), .B2(new_n353), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT38), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .A4(new_n430), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n424), .A2(new_n501), .A3(new_n425), .A4(new_n449), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n497), .A2(new_n430), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT37), .B1(new_n439), .B2(new_n443), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n383), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n473), .B1(new_n495), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n502), .A2(new_n505), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n474), .A2(new_n486), .A3(new_n489), .A4(new_n494), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(KEYINPUT89), .A4(new_n383), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n459), .B1(new_n472), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT93), .ZN(new_n514));
  INV_X1    g313(.A(G1gat), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n515), .A2(KEYINPUT16), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  OR3_X1    g317(.A1(new_n516), .A2(new_n518), .A3(G8gat), .ZN(new_n519));
  OAI21_X1  g318(.A(G8gat), .B1(new_n516), .B2(new_n518), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT91), .B(G29gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G36gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT14), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  OR3_X1    g325(.A1(new_n525), .A2(G29gat), .A3(G36gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n524), .A2(KEYINPUT15), .A3(new_n526), .A4(new_n527), .ZN(new_n531));
  XNOR2_X1  g330(.A(G43gat), .B(G50gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n522), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n519), .B2(new_n520), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(KEYINPUT13), .Z(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n535), .A2(KEYINPUT92), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n533), .A2(new_n534), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n543), .A2(KEYINPUT92), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(KEYINPUT92), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n537), .B1(new_n549), .B2(new_n522), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(KEYINPUT18), .A3(new_n540), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n542), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT18), .B1(new_n550), .B2(new_n540), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G113gat), .B(G141gat), .Z(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT90), .B(G197gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT11), .B(G169gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(KEYINPUT12), .Z(new_n560));
  NOR2_X1   g359(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n549), .A2(new_n522), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n538), .ZN(new_n564));
  INV_X1    g363(.A(new_n540), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n566), .A2(new_n542), .A3(new_n551), .A4(new_n560), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT94), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n569), .A3(new_n560), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n561), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  OR2_X1    g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT9), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G64gat), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n576), .A2(G57gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT96), .Z(new_n578));
  NOR2_X1   g377(.A1(new_n576), .A2(G57gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT95), .Z(new_n580));
  OAI21_X1  g379(.A(new_n575), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT9), .B1(new_n577), .B2(new_n579), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n572), .A3(new_n573), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(new_n261), .ZN(new_n589));
  INV_X1    g388(.A(new_n584), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n521), .B1(KEYINPUT21), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n589), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT97), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(new_n327), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n594), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n592), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT103), .ZN(new_n600));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  INV_X1    g402(.A(G92gat), .ZN(new_n604));
  AOI211_X1 g403(.A(new_n603), .B(new_n604), .C1(KEYINPUT99), .C2(KEYINPUT7), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(KEYINPUT99), .B2(KEYINPUT7), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT100), .B(G92gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(G99gat), .A2(G106gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n607), .A2(new_n603), .B1(KEYINPUT8), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n603), .A2(new_n604), .ZN(new_n610));
  OR3_X1    g409(.A1(new_n610), .A2(KEYINPUT99), .A3(KEYINPUT7), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n606), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G99gat), .B(G106gat), .Z(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(KEYINPUT101), .A3(new_n615), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n545), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(KEYINPUT98), .Z(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n619), .A2(new_n618), .B1(new_n544), .B2(new_n548), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n602), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n618), .A2(new_n619), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n549), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n629), .A2(new_n620), .A3(new_n624), .A4(new_n601), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n600), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  AOI211_X1 g435(.A(KEYINPUT103), .B(new_n634), .C1(new_n627), .C2(new_n630), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n627), .A2(new_n630), .A3(new_n634), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT102), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n616), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n614), .A2(KEYINPUT104), .A3(new_n615), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n590), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n614), .A2(new_n584), .A3(KEYINPUT104), .A4(new_n615), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT10), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n618), .A2(KEYINPUT10), .A3(new_n590), .A4(new_n619), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n642), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n642), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n646), .A2(new_n652), .A3(new_n647), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n651), .A2(new_n653), .A3(new_n657), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n599), .A2(new_n641), .A3(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n512), .A2(new_n571), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n426), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g466(.A(KEYINPUT16), .B(G8gat), .Z(new_n668));
  NAND3_X1  g467(.A1(new_n664), .A2(new_n474), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n664), .A2(new_n474), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(G8gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n669), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n671), .B1(new_n674), .B2(KEYINPUT42), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT105), .ZN(G1325gat));
  INV_X1    g475(.A(new_n664), .ZN(new_n677));
  INV_X1    g476(.A(new_n287), .ZN(new_n678));
  OR3_X1    g477(.A1(new_n677), .A2(G15gat), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n677), .B2(new_n468), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(G1326gat));
  NAND2_X1  g480(.A1(new_n383), .A2(KEYINPUT85), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n378), .A2(new_n460), .A3(new_n382), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n664), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT106), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  NOR2_X1   g487(.A1(new_n512), .A2(new_n641), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n599), .A2(new_n571), .A3(new_n661), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n691), .A2(new_n426), .A3(new_n523), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT45), .Z(new_n693));
  INV_X1    g492(.A(new_n690), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT44), .B1(new_n512), .B2(new_n641), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n455), .B(new_n696), .C1(new_n461), .C2(new_n462), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n468), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n684), .B2(new_n455), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n511), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n459), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT108), .B1(new_n638), .B2(new_n640), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n639), .B(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n707), .B(new_n708), .C1(new_n636), .C2(new_n637), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n703), .A2(new_n704), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n694), .B1(new_n695), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n523), .B1(new_n714), .B2(new_n426), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n693), .A2(new_n715), .ZN(G1328gat));
  NOR3_X1   g515(.A1(new_n691), .A2(G36gat), .A3(new_n454), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT46), .ZN(new_n718));
  OAI21_X1  g517(.A(G36gat), .B1(new_n714), .B2(new_n454), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(G1329gat));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721));
  INV_X1    g520(.A(G43gat), .ZN(new_n722));
  INV_X1    g521(.A(new_n468), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n713), .B2(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n691), .A2(G43gat), .A3(new_n678), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g526(.A(G50gat), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n713), .B2(new_n684), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n689), .A2(new_n728), .A3(new_n684), .A4(new_n690), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n729), .B1(KEYINPUT110), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n730), .B1(new_n733), .B2(KEYINPUT48), .ZN(new_n734));
  NAND2_X1  g533(.A1(KEYINPUT48), .A2(G50gat), .ZN(new_n735));
  INV_X1    g534(.A(new_n383), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n713), .B2(new_n736), .ZN(new_n737));
  OAI22_X1  g536(.A1(new_n732), .A2(KEYINPUT48), .B1(new_n734), .B2(new_n737), .ZN(G1331gat));
  AOI21_X1  g537(.A(new_n459), .B1(new_n511), .B2(new_n700), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n599), .A2(new_n641), .A3(new_n571), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n661), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n426), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g543(.A1(new_n742), .A2(new_n454), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT111), .ZN(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n742), .B2(new_n468), .ZN(new_n751));
  INV_X1    g550(.A(G71gat), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n662), .A2(new_n678), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n741), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT50), .Z(G1334gat));
  INV_X1    g555(.A(new_n684), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(G78gat), .Z(G1335gat));
  INV_X1    g558(.A(KEYINPUT112), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n567), .A2(KEYINPUT94), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n567), .A2(KEYINPUT94), .ZN(new_n762));
  OAI22_X1  g561(.A1(new_n761), .A2(new_n762), .B1(new_n554), .B2(new_n560), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n599), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n661), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n472), .A2(new_n511), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n702), .ZN(new_n768));
  INV_X1    g567(.A(new_n641), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n704), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n739), .A2(KEYINPUT44), .A3(new_n710), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n766), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n760), .B1(new_n772), .B2(new_n426), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n765), .B1(new_n695), .B2(new_n712), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(KEYINPUT112), .A3(new_n665), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(G85gat), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n764), .A2(new_n769), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n739), .B2(new_n777), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n665), .A2(new_n603), .A3(new_n661), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n776), .B1(new_n782), .B2(new_n783), .ZN(G1336gat));
  AOI21_X1  g583(.A(new_n607), .B1(new_n774), .B2(new_n474), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n474), .A2(new_n661), .A3(new_n604), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n782), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT52), .Z(G1337gat));
  NAND2_X1  g589(.A1(new_n779), .A2(new_n781), .ZN(new_n791));
  XNOR2_X1  g590(.A(KEYINPUT114), .B(G99gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n753), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n772), .A2(new_n468), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(new_n792), .ZN(G1338gat));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n662), .A2(G106gat), .A3(new_n383), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT115), .B1(new_n791), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  INV_X1    g598(.A(new_n797), .ZN(new_n800));
  AOI211_X1 g599(.A(new_n799), .B(new_n800), .C1(new_n779), .C2(new_n781), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G106gat), .B1(new_n772), .B2(new_n757), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n796), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(G106gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n805), .B1(new_n774), .B2(new_n736), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n797), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n796), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT116), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n806), .A2(new_n808), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n805), .B1(new_n774), .B2(new_n684), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n813), .A2(new_n798), .A3(new_n801), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n811), .B(new_n812), .C1(new_n814), .C2(new_n796), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n810), .A2(new_n815), .ZN(G1339gat));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  INV_X1    g616(.A(new_n648), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n652), .A3(new_n649), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n651), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n821), .B(new_n642), .C1(new_n648), .C2(new_n650), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n658), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n817), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n823), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n651), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(KEYINPUT55), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n763), .A2(new_n660), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n541), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n536), .A2(new_n538), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT117), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n540), .B2(new_n550), .ZN(new_n832));
  INV_X1    g631(.A(new_n559), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n834), .B(new_n661), .C1(new_n761), .C2(new_n762), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n828), .A2(new_n835), .B1(new_n705), .B2(new_n709), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n827), .A2(new_n660), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT55), .B1(new_n825), .B2(new_n826), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n570), .A2(new_n568), .B1(new_n832), .B2(new_n833), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n839), .A2(new_n705), .A3(new_n709), .A4(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n598), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n663), .A2(new_n763), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n660), .A3(new_n827), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n835), .B1(new_n848), .B2(new_n571), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n710), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n599), .B1(new_n850), .B2(new_n841), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT118), .B1(new_n851), .B2(new_n845), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n847), .A2(new_n852), .A3(new_n757), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n474), .A2(new_n426), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(KEYINPUT119), .A3(new_n287), .A4(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n847), .A2(new_n852), .A3(new_n287), .A4(new_n757), .ZN(new_n857));
  INV_X1    g656(.A(new_n854), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n855), .A2(new_n763), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(G113gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n847), .A2(new_n852), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n858), .A2(new_n384), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n571), .A2(new_n248), .A3(new_n247), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT120), .Z(new_n867));
  OAI22_X1  g666(.A1(new_n860), .A2(new_n861), .B1(new_n865), .B2(new_n867), .ZN(G1340gat));
  NAND4_X1  g667(.A1(new_n855), .A2(new_n859), .A3(G120gat), .A4(new_n661), .ZN(new_n869));
  INV_X1    g668(.A(G120gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n865), .B2(new_n662), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n869), .A2(new_n871), .ZN(G1341gat));
  AND3_X1   g671(.A1(new_n855), .A2(new_n599), .A3(new_n859), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n599), .A2(new_n261), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n873), .A2(new_n261), .B1(new_n865), .B2(new_n874), .ZN(G1342gat));
  NAND4_X1  g674(.A1(new_n863), .A2(new_n260), .A3(new_n769), .A4(new_n864), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT56), .Z(new_n877));
  NAND3_X1  g676(.A1(new_n855), .A2(new_n769), .A3(new_n859), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n878), .A2(KEYINPUT121), .A3(G134gat), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT121), .B1(new_n878), .B2(G134gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(G1343gat));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n847), .A2(new_n852), .A3(new_n882), .A4(new_n736), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n723), .A2(new_n858), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n849), .A2(new_n641), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n599), .B1(new_n886), .B2(new_n841), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n684), .B1(new_n887), .B2(new_n845), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n885), .B1(new_n888), .B2(KEYINPUT57), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G141gat), .B1(new_n890), .B2(new_n571), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n862), .A2(new_n383), .A3(new_n885), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n315), .A3(new_n763), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n313), .A3(new_n661), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n883), .A2(new_n889), .A3(new_n661), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n313), .A2(KEYINPUT59), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n769), .B1(new_n828), .B2(new_n835), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n839), .A2(new_n840), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n641), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n598), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n757), .B1(new_n908), .B2(new_n846), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n904), .B1(new_n909), .B2(KEYINPUT57), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n847), .A2(new_n852), .A3(KEYINPUT57), .A4(new_n736), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n886), .B1(new_n641), .B2(new_n906), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n845), .B1(new_n912), .B2(new_n598), .ZN(new_n913));
  OAI211_X1 g712(.A(KEYINPUT123), .B(new_n882), .C1(new_n913), .C2(new_n757), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n661), .A3(new_n884), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n903), .B1(new_n916), .B2(G148gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n896), .B1(new_n902), .B2(new_n917), .ZN(G1345gat));
  OAI21_X1  g717(.A(G155gat), .B1(new_n890), .B2(new_n598), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n892), .A2(new_n327), .A3(new_n599), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  NAND3_X1  g720(.A1(new_n892), .A2(new_n328), .A3(new_n769), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(new_n890), .B2(new_n710), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G162gat), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n890), .A2(new_n923), .A3(new_n710), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n384), .A2(new_n454), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n847), .A2(new_n852), .A3(new_n426), .A4(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n763), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n474), .A2(new_n426), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n857), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n571), .A2(new_n219), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1348gat));
  OAI21_X1  g734(.A(new_n220), .B1(new_n929), .B2(new_n662), .ZN(new_n936));
  NOR4_X1   g735(.A1(new_n932), .A2(new_n662), .A3(new_n678), .A4(new_n220), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n853), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT125), .Z(G1349gat));
  NAND3_X1  g739(.A1(new_n930), .A2(new_n203), .A3(new_n599), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n857), .A2(new_n598), .A3(new_n932), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n210), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n930), .A2(new_n204), .A3(new_n711), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n857), .A2(new_n641), .A3(new_n932), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n946), .A2(new_n204), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n204), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(G1351gat));
  INV_X1    g750(.A(G197gat), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n723), .A2(new_n454), .A3(new_n383), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n863), .A2(new_n426), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n954), .B2(new_n571), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n723), .A2(new_n932), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT126), .Z(new_n957));
  NAND4_X1  g756(.A1(new_n915), .A2(G197gat), .A3(new_n763), .A4(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n955), .A2(new_n958), .ZN(G1352gat));
  NAND3_X1  g758(.A1(new_n915), .A2(new_n661), .A3(new_n957), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G204gat), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n662), .A2(G204gat), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  OR3_X1    g762(.A1(new_n954), .A2(KEYINPUT62), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(KEYINPUT62), .B1(new_n954), .B2(new_n963), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n961), .A2(new_n964), .A3(new_n965), .ZN(G1353gat));
  OR3_X1    g765(.A1(new_n954), .A2(new_n296), .A3(new_n598), .ZN(new_n967));
  INV_X1    g766(.A(G211gat), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n723), .A2(new_n598), .A3(new_n932), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n915), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g769(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n974), .B1(new_n970), .B2(new_n972), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n967), .B1(new_n973), .B2(new_n975), .ZN(G1354gat));
  INV_X1    g775(.A(G218gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n977), .B1(new_n954), .B2(new_n710), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n915), .A2(G218gat), .A3(new_n769), .A4(new_n957), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(G1355gat));
endmodule


