//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n205), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(G197gat), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(G197gat), .B1(new_n206), .B2(new_n207), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT12), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(new_n207), .ZN(new_n212));
  INV_X1    g011(.A(G197gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT12), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n208), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(KEYINPUT87), .ZN(new_n221));
  INV_X1    g020(.A(G1gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G8gat), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n218), .B(KEYINPUT87), .C1(new_n219), .C2(G1gat), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n224), .B1(new_n223), .B2(new_n225), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(G43gat), .A2(G50gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(G43gat), .A2(G50gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT85), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G43gat), .ZN(new_n232));
  INV_X1    g031(.A(G50gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT85), .ZN(new_n235));
  NAND2_X1  g034(.A1(G43gat), .A2(G50gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT15), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT14), .ZN(new_n240));
  INV_X1    g039(.A(G29gat), .ZN(new_n241));
  INV_X1    g040(.A(G36gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT15), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n234), .A2(new_n246), .A3(new_n236), .ZN(new_n247));
  NAND2_X1  g046(.A1(G29gat), .A2(G36gat), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n239), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n246), .B1(new_n231), .B2(new_n237), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT86), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n243), .A2(new_n252), .A3(new_n244), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n248), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n243), .B2(new_n244), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT17), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n250), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n257), .B1(new_n250), .B2(new_n256), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n228), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G229gat), .A2(G233gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT88), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n223), .A2(new_n225), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G8gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n256), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n260), .A2(KEYINPUT18), .A3(new_n263), .A4(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n262), .B(KEYINPUT13), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n267), .A2(new_n268), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n265), .A2(new_n266), .B1(new_n256), .B2(new_n250), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n263), .A3(new_n269), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT18), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n217), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n278), .A2(new_n217), .A3(new_n270), .A4(new_n274), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT89), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT89), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n275), .A2(new_n282), .A3(new_n278), .A4(new_n217), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n279), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT21), .ZN(new_n286));
  AND2_X1   g085(.A1(G71gat), .A2(G78gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(G71gat), .A2(G78gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G57gat), .B(G64gat), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(G57gat), .A2(G64gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G57gat), .A2(G64gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G71gat), .B(G78gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n291), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n228), .B1(new_n286), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(new_n300), .B(KEYINPUT91), .Z(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n303));
  NAND2_X1  g102(.A1(new_n299), .A2(new_n286), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT90), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(G231gat), .A2(G233gat), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n307), .ZN(new_n309));
  XNOR2_X1  g108(.A(G127gat), .B(G155gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n310), .B1(new_n308), .B2(new_n309), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n303), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n306), .B(new_n307), .ZN(new_n315));
  INV_X1    g114(.A(new_n310), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n303), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n311), .A3(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(G183gat), .B(G211gat), .Z(new_n320));
  AND3_X1   g119(.A1(new_n314), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n314), .B2(new_n319), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n302), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n320), .ZN(new_n324));
  INV_X1    g123(.A(new_n319), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n318), .B1(new_n317), .B2(new_n311), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n314), .A2(new_n319), .A3(new_n320), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n301), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G232gat), .A2(G233gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT92), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT41), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G99gat), .A2(G106gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT8), .ZN(new_n335));
  NAND2_X1  g134(.A1(G85gat), .A2(G92gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT7), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G85gat), .ZN(new_n339));
  INV_X1    g138(.A(G92gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n335), .A2(new_n338), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G99gat), .B(G106gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  AND3_X1   g145(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI22_X1  g148(.A1(KEYINPUT8), .A2(new_n334), .B1(new_n339), .B2(new_n340), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n344), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n333), .B1(new_n268), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n258), .A2(new_n259), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n353), .B1(new_n354), .B2(new_n352), .ZN(new_n355));
  XNOR2_X1  g154(.A(G190gat), .B(G218gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n356), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n353), .B(new_n358), .C1(new_n354), .C2(new_n352), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n331), .A2(new_n332), .ZN(new_n361));
  XNOR2_X1  g160(.A(G134gat), .B(G162gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT93), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n365), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n323), .A2(new_n329), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT96), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n343), .A2(new_n345), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n349), .A2(new_n344), .A3(new_n350), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n371), .A2(new_n292), .A3(new_n372), .A4(new_n298), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n371), .A2(new_n372), .B1(new_n292), .B2(new_n298), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT94), .B(KEYINPUT10), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT95), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT95), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n292), .A2(new_n298), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n352), .A2(new_n380), .A3(KEYINPUT10), .A4(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n376), .A2(new_n377), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G230gat), .A2(G233gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n370), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(new_n382), .ZN(new_n387));
  INV_X1    g186(.A(new_n375), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(new_n373), .A3(new_n377), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(KEYINPUT96), .A3(new_n384), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n376), .B2(new_n384), .ZN(new_n393));
  XNOR2_X1  g192(.A(G120gat), .B(G148gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G176gat), .B(G204gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n383), .A2(new_n385), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n396), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n399), .B(new_n400), .C1(new_n376), .C2(new_n384), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n369), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT97), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n403), .A2(KEYINPUT97), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n285), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(KEYINPUT31), .B(G50gat), .Z(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(G197gat), .B(G204gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT22), .ZN(new_n411));
  XNOR2_X1  g210(.A(G211gat), .B(G218gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G211gat), .ZN(new_n415));
  INV_X1    g214(.A(G218gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n412), .B(new_n410), .C1(KEYINPUT22), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G155gat), .ZN(new_n420));
  INV_X1    g219(.A(G162gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(G155gat), .A2(G162gat), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT2), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(G141gat), .B(G148gat), .Z(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(KEYINPUT75), .ZN(new_n429));
  XNOR2_X1  g228(.A(G141gat), .B(G148gat), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n427), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT3), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT74), .B(KEYINPUT2), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n422), .A2(new_n424), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n433), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n419), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT80), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n414), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n411), .A2(KEYINPUT79), .A3(new_n413), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n418), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT3), .B1(new_n446), .B2(new_n440), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n428), .A2(KEYINPUT75), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n431), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n448), .A2(new_n449), .B1(new_n423), .B2(new_n426), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n422), .B(new_n424), .C1(new_n428), .C2(new_n435), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI22_X1  g251(.A1(new_n441), .A2(new_n442), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n441), .A2(new_n442), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n409), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT3), .B1(new_n419), .B2(new_n440), .ZN(new_n456));
  OAI211_X1 g255(.A(G228gat), .B(G233gat), .C1(new_n456), .C2(new_n452), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n457), .A2(new_n441), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(G22gat), .ZN(new_n460));
  INV_X1    g259(.A(G22gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n455), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G78gat), .B(G106gat), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n460), .B2(new_n462), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n408), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n460), .A2(new_n462), .ZN(new_n467));
  INV_X1    g266(.A(new_n463), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n470));
  INV_X1    g269(.A(new_n408), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT25), .ZN(new_n474));
  XOR2_X1   g273(.A(KEYINPUT65), .B(G169gat), .Z(new_n475));
  INV_X1    g274(.A(G176gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(KEYINPUT23), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G169gat), .A2(G176gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n205), .A2(new_n476), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT23), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT66), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(G169gat), .A2(G176gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT66), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT23), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n477), .B(new_n478), .C1(new_n481), .C2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT64), .ZN(new_n487));
  NAND2_X1  g286(.A1(G183gat), .A2(G190gat), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n474), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n478), .A2(KEYINPUT25), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(KEYINPUT23), .B2(new_n482), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n489), .A2(new_n488), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n486), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n493), .B(new_n495), .C1(new_n481), .C2(new_n484), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT67), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT26), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n482), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(KEYINPUT26), .B2(new_n479), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n479), .A2(KEYINPUT67), .A3(KEYINPUT26), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n478), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n488), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT68), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(KEYINPUT68), .B(new_n488), .C1(new_n501), .C2(new_n503), .ZN(new_n507));
  XNOR2_X1  g306(.A(KEYINPUT27), .B(G183gat), .ZN(new_n508));
  INV_X1    g307(.A(G190gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n510), .B(KEYINPUT28), .Z(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G120gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G113gat), .ZN(new_n515));
  INV_X1    g314(.A(G113gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G120gat), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT1), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G127gat), .B(G134gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT69), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G127gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G134gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n520), .B1(new_n525), .B2(new_n518), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n513), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G227gat), .ZN(new_n529));
  INV_X1    g328(.A(G233gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n497), .A2(new_n512), .A3(new_n526), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(G15gat), .B(G43gat), .Z(new_n534));
  XNOR2_X1  g333(.A(G71gat), .B(G99gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT33), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(KEYINPUT32), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n533), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n537), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n536), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(new_n533), .B2(KEYINPUT32), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT33), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n533), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n531), .B1(new_n528), .B2(new_n532), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n528), .ZN(new_n553));
  INV_X1    g352(.A(new_n532), .ZN(new_n554));
  OAI221_X1 g353(.A(new_n551), .B1(new_n529), .B2(new_n530), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n548), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n540), .A2(new_n541), .B1(new_n546), .B2(new_n544), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT84), .B1(new_n473), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n542), .A2(new_n556), .A3(new_n547), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n556), .B1(new_n542), .B2(new_n547), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT84), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n472), .A4(new_n466), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT73), .ZN(new_n568));
  INV_X1    g367(.A(new_n419), .ZN(new_n569));
  INV_X1    g368(.A(G226gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(new_n530), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n497), .A2(new_n512), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n440), .B1(new_n570), .B2(new_n530), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(new_n497), .B2(new_n512), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n569), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n497), .A2(new_n512), .A3(new_n571), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n511), .A2(new_n507), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n577), .A2(new_n506), .B1(new_n491), .B2(new_n496), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n576), .B(new_n419), .C1(new_n578), .C2(new_n573), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G8gat), .B(G36gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(G64gat), .B(G92gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT30), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n568), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n580), .A2(KEYINPUT73), .A3(KEYINPUT30), .A4(new_n584), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT30), .B1(new_n580), .B2(new_n584), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n587), .A2(new_n588), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT6), .ZN(new_n592));
  XNOR2_X1  g391(.A(G1gat), .B(G29gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT0), .ZN(new_n594));
  XNOR2_X1  g393(.A(G57gat), .B(G85gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  INV_X1    g395(.A(KEYINPUT76), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n526), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT3), .B1(new_n450), .B2(new_n451), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n515), .A2(new_n517), .ZN(new_n600));
  OAI221_X1 g399(.A(new_n522), .B1(new_n521), .B2(new_n524), .C1(KEYINPUT1), .C2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(KEYINPUT76), .A3(new_n520), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n598), .A2(new_n599), .A3(new_n439), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G225gat), .A2(G233gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n527), .A2(KEYINPUT4), .A3(new_n452), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n433), .A2(new_n601), .A3(new_n520), .A4(new_n438), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT4), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n603), .A2(new_n604), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT78), .ZN(new_n610));
  OR3_X1    g409(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT5), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n610), .B1(new_n609), .B2(KEYINPUT5), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n608), .A2(new_n605), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT77), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n614), .A2(new_n615), .A3(new_n604), .A4(new_n603), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT5), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n602), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n606), .B1(new_n618), .B2(new_n452), .ZN(new_n619));
  INV_X1    g418(.A(new_n604), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n609), .A2(KEYINPUT77), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n616), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI211_X1 g422(.A(new_n592), .B(new_n596), .C1(new_n613), .C2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n613), .A2(new_n623), .A3(new_n596), .ZN(new_n625));
  INV_X1    g424(.A(new_n612), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT5), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n596), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT6), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n624), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n591), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n562), .A2(new_n567), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT35), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT72), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n564), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT72), .B1(new_n559), .B2(new_n556), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n560), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n628), .A2(new_n629), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n639), .A2(new_n592), .A3(new_n625), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n628), .A2(KEYINPUT6), .A3(new_n629), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT35), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n643), .A3(new_n590), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n638), .A2(new_n644), .A3(new_n473), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n634), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT36), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n638), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n565), .A2(KEYINPUT36), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT83), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n575), .A2(new_n579), .A3(KEYINPUT37), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n653), .A2(new_n583), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT37), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT82), .B1(new_n580), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT82), .ZN(new_n657));
  AOI211_X1 g456(.A(new_n657), .B(KEYINPUT37), .C1(new_n575), .C2(new_n579), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n654), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT38), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n654), .B(new_n661), .C1(new_n656), .C2(new_n658), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n640), .A2(new_n641), .A3(new_n585), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n604), .B(new_n606), .C1(new_n618), .C2(new_n452), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT81), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(KEYINPUT81), .ZN(new_n668));
  INV_X1    g467(.A(new_n603), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n608), .A2(new_n605), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n620), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT39), .A4(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(KEYINPUT39), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(new_n596), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n672), .A2(KEYINPUT40), .A3(new_n673), .A4(new_n596), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n639), .A3(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n466), .B(new_n472), .C1(new_n590), .C2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n652), .B1(new_n665), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n631), .A2(new_n585), .A3(new_n660), .A4(new_n662), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n590), .A2(new_n678), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n466), .A2(new_n472), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n681), .A2(KEYINPUT83), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n473), .B1(new_n631), .B2(new_n591), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n651), .A2(new_n680), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n407), .B1(new_n647), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n631), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  NAND3_X1  g489(.A1(new_n687), .A2(new_n591), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(KEYINPUT42), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n687), .A2(new_n591), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(G8gat), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n692), .B1(new_n691), .B2(new_n695), .ZN(G1325gat));
  INV_X1    g495(.A(new_n651), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n687), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n638), .A2(G15gat), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n698), .A2(G15gat), .B1(new_n687), .B2(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT98), .Z(G1326gat));
  NAND2_X1  g500(.A1(new_n687), .A2(new_n473), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT43), .B(G22gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  AOI21_X1  g503(.A(new_n368), .B1(new_n647), .B2(new_n686), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n323), .A2(new_n329), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n707), .A2(new_n284), .A3(new_n402), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(G29gat), .A3(new_n642), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT45), .Z(new_n711));
  AND4_X1   g510(.A1(new_n651), .A2(new_n680), .A3(new_n684), .A4(new_n685), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n645), .B1(new_n633), .B2(KEYINPUT35), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT99), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT99), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n647), .A2(new_n715), .A3(new_n686), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n368), .A2(KEYINPUT44), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n366), .A2(new_n367), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n712), .B2(new_n713), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT44), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n708), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n642), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n711), .A2(new_n724), .ZN(G1328gat));
  NOR3_X1   g524(.A1(new_n709), .A2(G36gat), .A3(new_n590), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT46), .ZN(new_n727));
  OAI21_X1  g526(.A(G36gat), .B1(new_n723), .B2(new_n590), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1329gat));
  OAI21_X1  g528(.A(new_n232), .B1(new_n709), .B2(new_n638), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n697), .A2(G43gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n723), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT100), .B(KEYINPUT47), .Z(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1330gat));
  INV_X1    g533(.A(new_n708), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n683), .B(new_n735), .C1(new_n718), .C2(new_n721), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n473), .A2(new_n233), .ZN(new_n737));
  OAI22_X1  g536(.A1(new_n736), .A2(new_n233), .B1(new_n709), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT48), .B1(new_n738), .B2(KEYINPUT101), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n709), .A2(new_n737), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n722), .A2(new_n473), .A3(new_n708), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(G50gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT101), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n739), .A2(new_n745), .ZN(G1331gat));
  INV_X1    g545(.A(new_n402), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n369), .A2(new_n285), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n714), .A2(new_n716), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT102), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT102), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n714), .A2(new_n716), .A3(new_n751), .A4(new_n748), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n631), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G57gat), .ZN(G1332gat));
  INV_X1    g553(.A(KEYINPUT49), .ZN(new_n755));
  INV_X1    g554(.A(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n591), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT103), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n750), .A2(new_n752), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n756), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1333gat));
  NAND4_X1  g560(.A1(new_n750), .A2(G71gat), .A3(new_n697), .A4(new_n752), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n638), .B(KEYINPUT104), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n750), .A2(new_n752), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n765), .B2(G71gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n473), .A3(new_n752), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT105), .B(G78gat), .Z(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n707), .A2(new_n285), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n747), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n718), .B2(new_n721), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n642), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n720), .B2(new_n772), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n705), .A2(KEYINPUT51), .A3(new_n771), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n779), .A2(new_n780), .A3(KEYINPUT106), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT106), .B1(new_n779), .B2(new_n780), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n402), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n631), .A2(new_n339), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n777), .B1(new_n783), .B2(new_n784), .ZN(G1336gat));
  NAND2_X1  g584(.A1(new_n779), .A2(new_n780), .ZN(new_n786));
  AND4_X1   g585(.A1(new_n340), .A2(new_n786), .A3(new_n591), .A4(new_n402), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n340), .B1(new_n775), .B2(new_n591), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT52), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT107), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n776), .B2(new_n590), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n775), .A2(KEYINPUT107), .A3(new_n591), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n340), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n787), .A2(KEYINPUT52), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(G1337gat));
  XOR2_X1   g594(.A(KEYINPUT108), .B(G99gat), .Z(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n776), .B2(new_n651), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n638), .A2(new_n796), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n783), .B2(new_n798), .ZN(G1338gat));
  NOR2_X1   g598(.A1(new_n683), .A2(G106gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n786), .A2(new_n402), .A3(new_n800), .ZN(new_n801));
  AOI211_X1 g600(.A(new_n683), .B(new_n774), .C1(new_n718), .C2(new_n721), .ZN(new_n802));
  XOR2_X1   g601(.A(KEYINPUT109), .B(G106gat), .Z(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT110), .B1(new_n802), .B2(new_n803), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  OAI221_X1 g606(.A(new_n801), .B1(KEYINPUT110), .B2(KEYINPUT53), .C1(new_n802), .C2(new_n803), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(G1339gat));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n811));
  OR3_X1    g610(.A1(new_n272), .A2(new_n273), .A3(new_n271), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n260), .A2(new_n269), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n262), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n812), .A2(new_n814), .B1(new_n208), .B2(new_n214), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n281), .B2(new_n283), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n399), .A2(KEYINPUT54), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n390), .A2(new_n384), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n386), .A2(new_n820), .A3(new_n391), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n396), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT111), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n824), .A3(new_n396), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n819), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n719), .B(new_n816), .C1(new_n826), .C2(KEYINPUT55), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n821), .A2(new_n824), .A3(new_n396), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n824), .B1(new_n821), .B2(new_n396), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n828), .A2(new_n829), .B1(new_n818), .B2(new_n817), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n401), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n811), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n401), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n834), .B1(new_n826), .B2(KEYINPUT55), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n368), .B1(new_n830), .B2(new_n831), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT112), .A4(new_n816), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n816), .A2(new_n402), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n284), .B1(new_n830), .B2(new_n831), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n833), .B(new_n837), .C1(new_n840), .C2(new_n719), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n706), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n369), .A2(new_n285), .A3(new_n402), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n810), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  AOI211_X1 g644(.A(KEYINPUT113), .B(new_n843), .C1(new_n841), .C2(new_n706), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n562), .A2(new_n567), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n591), .A2(new_n642), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n516), .A3(new_n285), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n850), .A2(new_n638), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n683), .B1(new_n845), .B2(new_n846), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT114), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n858), .B(new_n683), .C1(new_n845), .C2(new_n846), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n855), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n516), .B1(new_n860), .B2(new_n285), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n853), .B1(new_n863), .B2(new_n864), .ZN(G1340gat));
  AOI21_X1  g664(.A(G120gat), .B1(new_n852), .B2(new_n402), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n747), .A2(new_n514), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n860), .B2(new_n867), .ZN(G1341gat));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n707), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n523), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n857), .A2(new_n859), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n706), .A2(new_n523), .ZN(new_n873));
  AND4_X1   g672(.A1(new_n871), .A2(new_n872), .A3(new_n854), .A4(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n871), .B1(new_n860), .B2(new_n873), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT117), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n878), .B(new_n870), .C1(new_n874), .C2(new_n875), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(G1342gat));
  NOR4_X1   g679(.A1(new_n848), .A2(G134gat), .A3(new_n591), .A4(new_n368), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n847), .A2(new_n631), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT56), .ZN(new_n883));
  INV_X1    g682(.A(G134gat), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n860), .B2(new_n719), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886));
  OR3_X1    g685(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n883), .B2(new_n885), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1343gat));
  NOR2_X1   g688(.A1(new_n697), .A2(new_n683), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n847), .A2(new_n631), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT119), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n847), .A2(new_n893), .A3(new_n631), .A4(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n284), .A2(G141gat), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n895), .A2(new_n591), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n842), .A2(new_n844), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n473), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n697), .B(new_n850), .C1(new_n899), .C2(KEYINPUT57), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n847), .A2(new_n473), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n900), .B(new_n285), .C1(new_n901), .C2(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G141gat), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n891), .A2(new_n591), .A3(new_n896), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n902), .B2(G141gat), .ZN(new_n907));
  OAI22_X1  g706(.A1(new_n897), .A2(new_n905), .B1(new_n907), .B2(new_n904), .ZN(G1344gat));
  NOR2_X1   g707(.A1(new_n895), .A2(new_n591), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n402), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(G148gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n900), .B1(new_n901), .B2(KEYINPUT57), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n911), .B1(new_n913), .B2(new_n747), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n284), .B1(new_n405), .B2(new_n406), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n840), .A2(new_n719), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n827), .A2(new_n832), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n706), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n915), .A2(KEYINPUT120), .A3(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n473), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT120), .B1(new_n915), .B2(new_n918), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n901), .A2(KEYINPUT57), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n651), .A2(KEYINPUT59), .A3(new_n402), .A4(new_n849), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n914), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n910), .A2(new_n912), .B1(new_n927), .B2(G148gat), .ZN(G1345gat));
  NAND3_X1  g727(.A1(new_n909), .A2(new_n420), .A3(new_n707), .ZN(new_n929));
  OAI21_X1  g728(.A(G155gat), .B1(new_n913), .B2(new_n706), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1346gat));
  NOR3_X1   g730(.A1(new_n591), .A2(G162gat), .A3(new_n368), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n892), .A2(new_n894), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n913), .A2(new_n368), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n421), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g736(.A(KEYINPUT121), .B(new_n933), .C1(new_n934), .C2(new_n421), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1347gat));
  NAND3_X1  g738(.A1(new_n562), .A2(new_n567), .A3(new_n591), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n642), .B1(new_n845), .B2(new_n846), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT122), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT122), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n943), .B(new_n642), .C1(new_n845), .C2(new_n846), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n940), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n475), .A3(new_n285), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n591), .A2(new_n642), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n763), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n872), .A2(new_n285), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n949), .B2(new_n205), .ZN(G1348gat));
  NOR2_X1   g749(.A1(new_n747), .A2(new_n476), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n872), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT124), .ZN(new_n953));
  AOI21_X1  g752(.A(G176gat), .B1(new_n945), .B2(new_n402), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n954), .A2(KEYINPUT123), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(KEYINPUT123), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(G1349gat));
  NAND3_X1  g756(.A1(new_n872), .A2(new_n707), .A3(new_n948), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G183gat), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n707), .A2(new_n508), .ZN(new_n960));
  AOI22_X1  g759(.A1(new_n945), .A2(new_n960), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n961));
  OR2_X1    g760(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n959), .B2(new_n961), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(G1350gat));
  AND3_X1   g764(.A1(new_n872), .A2(new_n719), .A3(new_n948), .ZN(new_n966));
  XNOR2_X1  g765(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n967));
  OR3_X1    g766(.A1(new_n966), .A2(new_n509), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n966), .B2(new_n509), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n945), .A2(new_n509), .A3(new_n719), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(G1351gat));
  NAND2_X1  g770(.A1(new_n942), .A2(new_n944), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n890), .A2(new_n591), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n972), .A2(new_n213), .A3(new_n285), .A4(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n697), .A2(new_n947), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n925), .A2(new_n284), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n975), .B1(new_n978), .B2(new_n213), .ZN(G1352gat));
  NAND4_X1  g778(.A1(new_n923), .A2(new_n924), .A3(new_n402), .A4(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(G204gat), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n747), .A2(G204gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n972), .A2(new_n974), .A3(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  OAI22_X1  g787(.A1(new_n982), .A2(new_n983), .B1(new_n987), .B2(new_n988), .ZN(G1353gat));
  NAND4_X1  g788(.A1(new_n972), .A2(new_n415), .A3(new_n707), .A4(new_n974), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n923), .A2(new_n924), .A3(new_n707), .A4(new_n976), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(G1354gat));
  NAND4_X1  g793(.A1(new_n972), .A2(new_n416), .A3(new_n719), .A4(new_n974), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n925), .A2(new_n368), .A3(new_n977), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n996), .B2(new_n416), .ZN(G1355gat));
endmodule


