//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1187, new_n1188,
    new_n1189, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n206), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n215), .A2(new_n216), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n222), .B1(new_n215), .B2(new_n216), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G87), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n206), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  INV_X1    g0029(.A(G77), .ZN(new_n230));
  INV_X1    g0030(.A(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G107), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n229), .B1(new_n230), .B2(new_n231), .C1(new_n232), .C2(new_n214), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n210), .B1(new_n228), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT1), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n223), .A2(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  NAND2_X1  g0051(.A1(KEYINPUT66), .A2(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT8), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(new_n208), .A3(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n217), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n207), .B2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G50), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n260), .B(new_n262), .C1(G50), .C2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT9), .ZN(new_n265));
  INV_X1    g0065(.A(G200), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n271), .A2(new_n267), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n272), .A2(G226), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n280), .A2(G223), .B1(G77), .B2(new_n278), .ZN(new_n281));
  INV_X1    g0081(.A(G222), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n281), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  AOI211_X1 g0088(.A(new_n269), .B(new_n273), .C1(new_n288), .C2(new_n270), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n265), .B1(new_n266), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n289), .A2(G190), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n290), .A2(new_n291), .B1(KEYINPUT69), .B2(KEYINPUT10), .ZN(new_n292));
  NAND2_X1  g0092(.A1(KEYINPUT69), .A2(KEYINPUT10), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n264), .B1(new_n289), .B2(G169), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G97), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n286), .A2(G232), .ZN(new_n302));
  INV_X1    g0102(.A(G226), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n301), .B1(new_n302), .B2(new_n279), .C1(new_n303), .C2(new_n287), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n270), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n269), .B1(new_n272), .B2(G238), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g0107(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n305), .A2(new_n308), .A3(new_n306), .ZN(new_n310));
  OAI21_X1  g0110(.A(G169), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT14), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT14), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n313), .B(G169), .C1(new_n309), .C2(new_n310), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n305), .A2(new_n306), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n310), .B1(KEYINPUT13), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G179), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n261), .A2(G68), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT12), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n263), .B2(G68), .ZN(new_n321));
  INV_X1    g0121(.A(new_n263), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(KEYINPUT12), .A3(new_n225), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT71), .ZN(new_n325));
  INV_X1    g0125(.A(new_n255), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n202), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n208), .A2(G33), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n328), .A2(new_n230), .B1(new_n208), .B2(G68), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n259), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT11), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n318), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n316), .A2(G190), .ZN(new_n334));
  INV_X1    g0134(.A(new_n332), .ZN(new_n335));
  OAI21_X1  g0135(.A(G200), .B1(new_n309), .B2(new_n310), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n272), .A2(G244), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n280), .A2(G238), .B1(G107), .B2(new_n278), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT65), .B(G1698), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n302), .ZN(new_n342));
  AOI211_X1 g0142(.A(new_n269), .B(new_n339), .C1(new_n342), .C2(new_n270), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G190), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n266), .B2(new_n343), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT15), .B(G87), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n346), .A2(new_n328), .B1(new_n208), .B2(new_n230), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT8), .B(G58), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT67), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n349), .B2(new_n255), .ZN(new_n350));
  INV_X1    g0150(.A(new_n259), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n261), .A2(G77), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G77), .B2(new_n263), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT68), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n345), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n343), .A2(G169), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n295), .B2(new_n343), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n356), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NOR4_X1   g0161(.A1(new_n300), .A2(new_n338), .A3(new_n357), .A4(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT75), .ZN(new_n363));
  OR2_X1    g0163(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n364));
  NAND2_X1  g0164(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(G223), .A3(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n303), .A2(new_n279), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n278), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G87), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n363), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n367), .B1(new_n285), .B2(G223), .ZN(new_n373));
  OAI211_X1 g0173(.A(KEYINPUT75), .B(new_n370), .C1(new_n373), .C2(new_n278), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n374), .A3(new_n270), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n269), .B1(new_n272), .B2(G232), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n375), .A2(G190), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n266), .B1(new_n375), .B2(new_n376), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G58), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n225), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(new_n201), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(G20), .B1(G159), .B2(new_n255), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n286), .B2(G20), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n386));
  AOI211_X1 g0186(.A(KEYINPUT72), .B(new_n225), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT72), .ZN(new_n388));
  AOI21_X1  g0188(.A(G20), .B1(new_n275), .B2(new_n277), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n208), .A2(KEYINPUT7), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n389), .A2(KEYINPUT7), .B1(new_n286), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n388), .B1(new_n391), .B2(G68), .ZN(new_n392));
  OAI211_X1 g0192(.A(KEYINPUT16), .B(new_n383), .C1(new_n387), .C2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n383), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n286), .A2(KEYINPUT73), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT73), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n390), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT74), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n395), .A2(KEYINPUT74), .A3(new_n398), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n402), .A3(new_n385), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n394), .B1(new_n403), .B2(G68), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n393), .B(new_n259), .C1(new_n404), .C2(KEYINPUT16), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n253), .A2(new_n263), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n253), .B2(new_n261), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n379), .A2(new_n405), .A3(KEYINPUT77), .A4(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n391), .A2(G68), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT72), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n391), .A2(new_n388), .A3(G68), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n394), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n351), .B1(new_n415), .B2(KEYINPUT16), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n402), .A2(new_n385), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT74), .B1(new_n395), .B2(new_n398), .ZN(new_n418));
  OAI21_X1  g0218(.A(G68), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT16), .B1(new_n419), .B2(new_n383), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n411), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n422), .A2(KEYINPUT77), .A3(KEYINPUT17), .A4(new_n379), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n410), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n393), .A2(new_n259), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n407), .B1(new_n425), .B2(new_n420), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n375), .A2(G179), .A3(new_n376), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n375), .A2(new_n376), .ZN(new_n428));
  INV_X1    g0228(.A(G169), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT18), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(KEYINPUT18), .A3(new_n430), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n431), .B1(KEYINPUT76), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT76), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n426), .A2(new_n434), .A3(KEYINPUT18), .A4(new_n430), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n424), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n362), .A2(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n280), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n278), .A2(new_n341), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(KEYINPUT4), .A3(G244), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT4), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n287), .B2(new_n231), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n271), .B1(new_n443), .B2(KEYINPUT78), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT78), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n438), .A2(new_n440), .A3(new_n442), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT5), .B(G41), .ZN(new_n448));
  INV_X1    g0248(.A(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(G1), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n451), .A2(new_n268), .A3(new_n270), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n270), .B1(new_n450), .B2(new_n448), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n452), .B1(G257), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n447), .A2(new_n295), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n263), .A2(G97), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n207), .A2(G33), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n351), .A2(new_n263), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n456), .B1(new_n459), .B2(G97), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT6), .ZN(new_n461));
  INV_X1    g0261(.A(G97), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n461), .A2(new_n462), .A3(G107), .ZN(new_n463));
  XNOR2_X1  g0263(.A(G97), .B(G107), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n465), .A2(new_n208), .B1(new_n230), .B2(new_n326), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n403), .B2(G107), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n460), .B1(new_n467), .B2(new_n351), .ZN(new_n468));
  INV_X1    g0268(.A(new_n454), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n444), .B2(new_n446), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n455), .B(new_n468), .C1(G169), .C2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n447), .A2(G190), .A3(new_n454), .ZN(new_n472));
  INV_X1    g0272(.A(new_n460), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n403), .A2(G107), .ZN(new_n474));
  INV_X1    g0274(.A(new_n466), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n473), .B1(new_n476), .B2(new_n259), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n472), .B(new_n477), .C1(new_n266), .C2(new_n470), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n286), .A2(G244), .A3(G1698), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G116), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n479), .B(new_n480), .C1(new_n287), .C2(new_n226), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT79), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n439), .A2(G238), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n479), .A4(new_n480), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n270), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n450), .A2(new_n206), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n271), .A2(new_n488), .B1(G274), .B2(new_n450), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n295), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n286), .A2(new_n208), .A3(G68), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT19), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n328), .B2(new_n462), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n227), .A2(new_n462), .A3(new_n232), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n494), .B(KEYINPUT80), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n301), .A2(new_n492), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(G20), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n491), .B(new_n493), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n259), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n346), .A2(new_n322), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(new_n500), .C1(new_n346), .C2(new_n458), .ZN(new_n501));
  INV_X1    g0301(.A(new_n489), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n502), .B1(new_n486), .B2(new_n270), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n490), .B(new_n501), .C1(G169), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n487), .A2(G190), .A3(new_n489), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n459), .A2(G87), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n499), .A2(new_n500), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n505), .B(new_n507), .C1(new_n266), .C2(new_n503), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n471), .A2(new_n478), .A3(new_n504), .A4(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT81), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n451), .A2(new_n271), .ZN(new_n511));
  INV_X1    g0311(.A(G270), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n453), .A2(KEYINPUT81), .A3(G270), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n286), .A2(G264), .A3(G1698), .ZN(new_n516));
  INV_X1    g0316(.A(G303), .ZN(new_n517));
  OAI221_X1 g0317(.A(new_n516), .B1(new_n517), .B2(new_n286), .C1(new_n287), .C2(new_n213), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n270), .ZN(new_n519));
  INV_X1    g0319(.A(new_n452), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n515), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G200), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT83), .ZN(new_n523));
  AOI21_X1  g0323(.A(G20), .B1(G33), .B2(G283), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(G33), .B2(new_n462), .ZN(new_n525));
  INV_X1    g0325(.A(G116), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G20), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n259), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT20), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n263), .A2(G116), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n459), .B2(G116), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n522), .A2(new_n523), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n452), .B1(new_n518), .B2(new_n270), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n266), .B1(new_n536), .B2(new_n515), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT83), .B1(new_n537), .B2(new_n533), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(G190), .A3(new_n515), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT82), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n429), .B1(new_n530), .B2(new_n532), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n521), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n533), .A2(new_n536), .A3(G179), .A4(new_n515), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n542), .B1(new_n521), .B2(new_n543), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n232), .B1(KEYINPUT84), .B2(KEYINPUT25), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n263), .ZN(new_n550));
  NAND2_X1  g0350(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n458), .A2(new_n232), .ZN(new_n553));
  OR3_X1    g0353(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT85), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT85), .B1(new_n552), .B2(new_n553), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n480), .A2(G20), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT23), .B1(new_n232), .B2(G20), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n232), .A2(KEYINPUT23), .A3(G20), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n286), .A2(new_n208), .A3(G87), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n563), .A2(KEYINPUT22), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(KEYINPUT22), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT24), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n259), .B1(new_n566), .B2(KEYINPUT24), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n556), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XOR2_X1   g0370(.A(KEYINPUT86), .B(G294), .Z(new_n571));
  AOI22_X1  g0371(.A1(new_n280), .A2(G257), .B1(G33), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n439), .A2(G250), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n270), .B1(G264), .B2(new_n453), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n520), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n429), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n295), .A3(new_n520), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n570), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n576), .A2(G200), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n564), .A2(new_n565), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n582), .B2(new_n562), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(new_n259), .A3(new_n567), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n575), .A2(G190), .A3(new_n520), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n580), .A2(new_n584), .A3(new_n556), .A4(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n540), .A2(new_n548), .A3(new_n579), .A4(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n509), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n437), .A2(new_n588), .ZN(G372));
  NAND2_X1  g0389(.A1(new_n426), .A2(new_n430), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT18), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n592), .A2(new_n432), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n333), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n337), .B1(new_n595), .B2(new_n361), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n594), .B1(new_n596), .B2(new_n424), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n298), .B1(new_n597), .B2(new_n294), .ZN(new_n598));
  INV_X1    g0398(.A(new_n437), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n504), .A2(new_n508), .ZN(new_n600));
  INV_X1    g0400(.A(new_n471), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT26), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n504), .A2(new_n508), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT26), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n603), .A2(new_n471), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n504), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n471), .A2(new_n478), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n607), .A2(KEYINPUT87), .A3(new_n600), .A4(new_n586), .ZN(new_n608));
  INV_X1    g0408(.A(new_n548), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n579), .A2(KEYINPUT88), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT88), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n570), .A2(new_n577), .A3(new_n611), .A4(new_n578), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n609), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n600), .A2(new_n471), .A3(new_n478), .A4(new_n586), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT87), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n606), .B1(new_n608), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n598), .B1(new_n599), .B2(new_n617), .ZN(G369));
  AND2_X1   g0418(.A1(new_n208), .A2(G13), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n207), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT89), .ZN(new_n621));
  OR2_X1    g0421(.A1(new_n621), .A2(KEYINPUT27), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(KEYINPUT27), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(G213), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(G343), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(new_n534), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n609), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n540), .A2(new_n548), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n630), .B2(new_n628), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G330), .ZN(new_n632));
  INV_X1    g0432(.A(new_n579), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n626), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n570), .A2(new_n626), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n579), .A2(new_n586), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n548), .A2(new_n626), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n579), .A3(new_n586), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n610), .A2(new_n612), .A3(new_n627), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n639), .A2(new_n643), .ZN(G399));
  NOR2_X1   g0444(.A1(new_n212), .A2(G41), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n495), .A2(new_n526), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(G1), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n220), .B2(new_n646), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT28), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT92), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n617), .B2(new_n626), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT29), .ZN(new_n654));
  INV_X1    g0454(.A(new_n586), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n615), .B1(new_n509), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n613), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n608), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n504), .ZN(new_n659));
  INV_X1    g0459(.A(new_n605), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n604), .B1(new_n603), .B2(new_n471), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(KEYINPUT92), .A3(new_n627), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n653), .A2(new_n654), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT93), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT93), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n653), .A2(new_n667), .A3(new_n654), .A4(new_n664), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n609), .A2(new_n633), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n614), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n626), .B1(new_n662), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT29), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n666), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT91), .B1(new_n588), .B2(new_n627), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT91), .ZN(new_n675));
  NOR4_X1   g0475(.A1(new_n509), .A2(new_n587), .A3(new_n675), .A4(new_n626), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT30), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n503), .A2(KEYINPUT90), .A3(new_n575), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n521), .A2(new_n295), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n470), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT90), .B1(new_n503), .B2(new_n575), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n681), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n470), .A2(new_n679), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(KEYINPUT30), .A4(new_n678), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n576), .A2(new_n295), .A3(new_n521), .ZN(new_n686));
  OR3_X1    g0486(.A1(new_n686), .A2(new_n470), .A3(new_n503), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n682), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT31), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n688), .A2(new_n689), .A3(new_n626), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n688), .B2(new_n626), .ZN(new_n691));
  OAI22_X1  g0491(.A1(new_n674), .A2(new_n676), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G330), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n673), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n651), .B1(new_n698), .B2(G1), .ZN(G364));
  AOI21_X1  g0499(.A(new_n207), .B1(new_n619), .B2(G45), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n645), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n631), .B2(G330), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(G330), .B2(new_n631), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n211), .A2(new_n286), .ZN(new_n705));
  INV_X1    g0505(.A(G355), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n705), .A2(new_n706), .B1(G116), .B2(new_n211), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n212), .A2(new_n286), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n449), .B2(new_n221), .ZN(new_n710));
  OR2_X1    g0510(.A1(new_n247), .A2(new_n449), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G13), .A2(G33), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n217), .B1(G20), .B2(new_n429), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n702), .B1(new_n712), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(G20), .A2(G179), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n720), .B(KEYINPUT94), .Z(new_n721));
  INV_X1    g0521(.A(G190), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n266), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(G190), .A3(new_n266), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n725), .A2(new_n225), .B1(new_n380), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n721), .A2(G190), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n266), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n727), .B1(G50), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G179), .A2(G200), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(G20), .A3(new_n722), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G159), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT32), .ZN(new_n735));
  NOR4_X1   g0535(.A1(new_n208), .A2(new_n722), .A3(new_n266), .A4(G179), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n286), .B1(new_n737), .B2(new_n227), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n731), .A2(G190), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G97), .ZN(new_n741));
  NOR4_X1   g0541(.A1(new_n208), .A2(new_n266), .A3(G179), .A4(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n741), .B1(new_n743), .B2(new_n232), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n735), .A2(new_n738), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n723), .A2(G200), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n747), .A2(KEYINPUT95), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(KEYINPUT95), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n730), .B(new_n745), .C1(new_n751), .C2(new_n230), .ZN(new_n752));
  XNOR2_X1  g0552(.A(KEYINPUT33), .B(G317), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G326), .A2(new_n729), .B1(new_n724), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n746), .A2(G311), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n286), .B1(new_n733), .B2(G329), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n517), .B2(new_n737), .ZN(new_n757));
  INV_X1    g0557(.A(new_n571), .ZN(new_n758));
  INV_X1    g0558(.A(new_n740), .ZN(new_n759));
  INV_X1    g0559(.A(G283), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n758), .A2(new_n759), .B1(new_n743), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n726), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G322), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n754), .A2(new_n755), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n752), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n719), .B1(new_n766), .B2(new_n716), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n715), .B(KEYINPUT96), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n631), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n704), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(G396));
  NAND2_X1  g0571(.A1(new_n361), .A2(new_n627), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n356), .A2(new_n626), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n360), .B1(new_n773), .B2(new_n357), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n653), .A2(new_n664), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n775), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n663), .A2(new_n627), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n702), .B1(new_n779), .B2(new_n696), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n776), .A2(new_n695), .A3(new_n778), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n716), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G137), .A2(new_n729), .B1(new_n763), .B2(G143), .ZN(new_n784));
  INV_X1    g0584(.A(G150), .ZN(new_n785));
  INV_X1    g0585(.A(G159), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n784), .B1(new_n785), .B2(new_n725), .C1(new_n751), .C2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT97), .B(KEYINPUT34), .Z(new_n788));
  XNOR2_X1  g0588(.A(new_n787), .B(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G132), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n286), .B1(new_n732), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(G58), .B2(new_n740), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n736), .A2(G50), .B1(new_n742), .B2(G68), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n789), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n741), .B(new_n278), .C1(new_n795), .C2(new_n732), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n736), .A2(G107), .B1(new_n742), .B2(G87), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(G303), .C2(new_n729), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G283), .A2(new_n724), .B1(new_n763), .B2(G294), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(new_n751), .C2(new_n526), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n783), .B1(new_n794), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n716), .A2(new_n713), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n702), .B1(G77), .B2(new_n804), .ZN(new_n805));
  OR3_X1    g0605(.A1(new_n802), .A2(KEYINPUT98), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(KEYINPUT98), .B1(new_n802), .B2(new_n805), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n775), .A2(new_n713), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n782), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G384));
  INV_X1    g0611(.A(new_n465), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT35), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(KEYINPUT35), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n813), .A2(G116), .A3(new_n218), .A4(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT36), .Z(new_n816));
  OR3_X1    g0616(.A1(new_n220), .A2(new_n230), .A3(new_n381), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n202), .A2(G68), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n207), .B(G13), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n422), .A2(new_n379), .ZN(new_n821));
  INV_X1    g0621(.A(new_n624), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n426), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n821), .A2(new_n590), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(KEYINPUT37), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n415), .A2(KEYINPUT16), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n407), .B1(new_n826), .B2(new_n425), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n430), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n822), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n821), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n825), .B1(KEYINPUT37), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n410), .A2(new_n423), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n432), .A2(KEYINPUT76), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n834), .A2(new_n435), .A3(new_n592), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n829), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT99), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT99), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n839), .B(new_n829), .C1(new_n833), .C2(new_n835), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n832), .B(KEYINPUT38), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT100), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n839), .B1(new_n436), .B2(new_n829), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n836), .A2(KEYINPUT99), .A3(new_n837), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n831), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(KEYINPUT100), .A3(KEYINPUT38), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n846), .A2(KEYINPUT101), .A3(KEYINPUT38), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT101), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n832), .B1(new_n838), .B2(new_n840), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n843), .B(new_n847), .C1(new_n848), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n778), .A2(new_n772), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n627), .A2(new_n335), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n318), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n338), .B2(new_n856), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n853), .A2(new_n860), .B1(new_n593), .B2(new_n624), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n593), .B1(new_n862), .B2(new_n424), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n833), .A2(KEYINPUT103), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n823), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT102), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n824), .A2(new_n866), .A3(KEYINPUT37), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n866), .B1(new_n824), .B2(KEYINPUT37), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n867), .A2(new_n868), .A3(new_n825), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n851), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n870), .A2(new_n841), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n853), .B2(KEYINPUT39), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n333), .A2(new_n626), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n861), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n666), .A2(new_n437), .A3(new_n668), .A4(new_n672), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n877), .A2(new_n598), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n876), .B(new_n878), .Z(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n870), .A2(new_n841), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n692), .A2(new_n777), .A3(new_n858), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n880), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n853), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n437), .A2(new_n692), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(G330), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n879), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n207), .B2(new_n619), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n879), .A2(new_n890), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n820), .B1(new_n892), .B2(new_n893), .ZN(G367));
  OR2_X1    g0694(.A1(new_n627), .A2(new_n507), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n600), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n504), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n471), .A2(new_n627), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT105), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n607), .B1(new_n477), .B2(new_n627), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OR3_X1    g0702(.A1(new_n902), .A2(KEYINPUT42), .A3(new_n641), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n471), .B1(new_n902), .B2(new_n579), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n627), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT42), .B1(new_n902), .B2(new_n641), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n905), .A2(KEYINPUT106), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT106), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n898), .B(new_n903), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT107), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n909), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n897), .B(KEYINPUT43), .Z(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n639), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n915), .B1(new_n916), .B2(new_n902), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n902), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n911), .A2(new_n918), .A3(new_n914), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n902), .A2(new_n643), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT44), .Z(new_n921));
  NOR2_X1   g0721(.A1(new_n902), .A2(new_n643), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT45), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n916), .A2(KEYINPUT108), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n641), .B1(new_n637), .B2(new_n640), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n632), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n698), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n645), .B(KEYINPUT41), .Z(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n917), .B(new_n919), .C1(new_n701), .C2(new_n932), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n717), .B1(new_n211), .B2(new_n346), .C1(new_n709), .C2(new_n243), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n934), .A2(new_n702), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n737), .A2(new_n380), .B1(new_n759), .B2(new_n225), .ZN(new_n936));
  INV_X1    g0736(.A(G137), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n286), .B1(new_n937), .B2(new_n732), .C1(new_n743), .C2(new_n230), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n936), .B(new_n938), .C1(new_n724), .C2(G159), .ZN(new_n939));
  AOI22_X1  g0739(.A1(G143), .A2(new_n729), .B1(new_n763), .B2(G150), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n939), .B(new_n940), .C1(new_n751), .C2(new_n202), .ZN(new_n941));
  AOI22_X1  g0741(.A1(G311), .A2(new_n729), .B1(new_n724), .B2(new_n571), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n517), .B2(new_n726), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n286), .B1(new_n733), .B2(G317), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n944), .B1(new_n759), .B2(new_n232), .C1(new_n462), .C2(new_n743), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n736), .A2(G116), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT46), .Z(new_n947));
  NOR3_X1   g0747(.A1(new_n943), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n751), .B2(new_n760), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT47), .Z(new_n951));
  OAI221_X1 g0751(.A(new_n935), .B1(new_n768), .B2(new_n897), .C1(new_n951), .C2(new_n783), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n933), .A2(new_n952), .ZN(G387));
  INV_X1    g0753(.A(new_n928), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n698), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n697), .A2(new_n928), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(new_n645), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n637), .A2(new_n768), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n349), .A2(new_n202), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT50), .Z(new_n960));
  OAI21_X1  g0760(.A(new_n449), .B1(new_n225), .B2(new_n230), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n648), .B2(KEYINPUT109), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n960), .B(new_n962), .C1(KEYINPUT109), .C2(new_n648), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n963), .B(new_n708), .C1(new_n449), .C2(new_n240), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(G107), .B2(new_n211), .C1(new_n648), .C2(new_n705), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n717), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n702), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n737), .A2(new_n230), .B1(new_n759), .B2(new_n346), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n286), .B1(new_n785), .B2(new_n732), .C1(new_n743), .C2(new_n462), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(new_n746), .C2(G68), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G159), .A2(new_n729), .B1(new_n724), .B2(new_n253), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n970), .B(new_n971), .C1(new_n202), .C2(new_n726), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n286), .B1(new_n733), .B2(G326), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n737), .A2(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G322), .A2(new_n729), .B1(new_n763), .B2(G317), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n795), .B2(new_n725), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(new_n750), .B2(G303), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n974), .B1(new_n977), .B2(KEYINPUT48), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(KEYINPUT48), .B2(new_n977), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT49), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n973), .B1(new_n526), .B2(new_n743), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n972), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n958), .B(new_n967), .C1(new_n983), .C2(new_n716), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n954), .B2(new_n701), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n957), .A2(new_n985), .ZN(G393));
  XNOR2_X1  g0786(.A(new_n924), .B(new_n639), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n955), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n988), .B(new_n645), .C1(new_n955), .C2(new_n926), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n708), .A2(new_n250), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n990), .B(new_n717), .C1(new_n462), .C2(new_n211), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n702), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT110), .Z(new_n993));
  AOI22_X1  g0793(.A1(new_n746), .A2(G294), .B1(G116), .B2(new_n740), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n517), .B2(new_n725), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT111), .Z(new_n996));
  AOI22_X1  g0796(.A1(G317), .A2(new_n729), .B1(new_n763), .B2(G311), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT52), .Z(new_n998));
  INV_X1    g0798(.A(G322), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n278), .B1(new_n732), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n743), .A2(new_n232), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G283), .C2(new_n736), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n996), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT112), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n750), .A2(new_n349), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n737), .A2(new_n225), .B1(new_n759), .B2(new_n230), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n278), .B1(new_n733), .B2(G143), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n227), .B2(new_n743), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1006), .B(new_n1008), .C1(new_n724), .C2(G50), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G150), .A2(new_n729), .B1(new_n763), .B2(G159), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT51), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1005), .B(new_n1009), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1004), .A2(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT113), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n716), .B1(new_n1016), .B2(KEYINPUT113), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n993), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n715), .B2(new_n902), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n987), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n701), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n989), .A2(new_n1022), .ZN(G390));
  AOI22_X1  g0823(.A1(new_n671), .A2(new_n774), .B1(new_n361), .B2(new_n627), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n875), .B1(new_n1024), .B2(new_n859), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n881), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n874), .B1(new_n854), .B2(new_n858), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1027), .B1(new_n873), .B2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n692), .A2(G330), .A3(new_n777), .A4(new_n858), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(KEYINPUT114), .ZN(new_n1032));
  AND4_X1   g0832(.A1(new_n540), .A2(new_n548), .A3(new_n579), .A4(new_n586), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1033), .A2(new_n607), .A3(new_n600), .A4(new_n627), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n675), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n588), .A2(KEYINPUT91), .A3(new_n627), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n688), .A2(new_n626), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT31), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n688), .A2(new_n689), .A3(new_n626), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n775), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT114), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1042), .A2(new_n1043), .A3(G330), .A4(new_n858), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1032), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(KEYINPUT115), .B1(new_n1030), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT115), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1045), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n872), .B(new_n1028), .C1(new_n853), .C2(KEYINPUT39), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1047), .B(new_n1048), .C1(new_n1049), .C2(new_n1027), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n872), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n1052), .A3(new_n1029), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1027), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n1054), .A3(new_n1031), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1046), .A2(new_n701), .A3(new_n1050), .A4(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n702), .B1(new_n253), .B2(new_n804), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n729), .A2(G128), .B1(G159), .B2(new_n740), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n278), .B1(new_n733), .B2(G125), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n202), .B2(new_n743), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT116), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n736), .A2(G150), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT53), .Z(new_n1064));
  AND3_X1   g0864(.A1(new_n1058), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n725), .A2(new_n937), .B1(new_n790), .B2(new_n726), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1061), .B2(new_n1060), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(KEYINPUT54), .B(G143), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1065), .B(new_n1067), .C1(new_n751), .C2(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n751), .A2(new_n462), .B1(new_n232), .B2(new_n725), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(KEYINPUT117), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n286), .B1(new_n736), .B2(G87), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT118), .Z(new_n1073));
  INV_X1    g0873(.A(G294), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n743), .A2(new_n225), .B1(new_n1074), .B2(new_n732), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G77), .B2(new_n740), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n526), .B2(new_n726), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1073), .B(new_n1077), .C1(G283), .C2(new_n729), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1071), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1070), .A2(KEYINPUT117), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1069), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1057), .B1(new_n1081), .B2(new_n716), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n873), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1082), .B1(new_n1083), .B2(new_n714), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1056), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1046), .A2(new_n1050), .A3(new_n1055), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n437), .A2(new_n695), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n877), .A2(new_n598), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1024), .A2(new_n1031), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n858), .B1(new_n1042), .B2(G330), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1090), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1045), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1091), .B1(new_n1093), .B2(new_n854), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1088), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n646), .B1(new_n1086), .B2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1046), .A2(new_n1050), .A3(new_n1055), .A4(new_n1095), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1085), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(G378));
  INV_X1    g0900(.A(new_n1088), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT57), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n822), .A2(new_n264), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n300), .B(new_n1104), .Z(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n886), .B2(new_n694), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1106), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1105), .B(new_n1109), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n843), .A2(new_n847), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT101), .B1(new_n846), .B2(KEYINPUT38), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n850), .A2(new_n849), .A3(new_n851), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n884), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1110), .B(G330), .C1(new_n1115), .C2(new_n883), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1108), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n876), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1083), .A2(new_n874), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1119), .A2(new_n1108), .A3(new_n861), .A4(new_n1116), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1103), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1102), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n876), .A2(KEYINPUT122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1117), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n876), .A2(new_n1108), .A3(KEYINPUT122), .A4(new_n1116), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1101), .B2(new_n1098), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1122), .B(new_n645), .C1(new_n1127), .C2(KEYINPUT57), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n702), .B1(G50), .B2(new_n804), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT121), .Z(new_n1130));
  NAND2_X1  g0930(.A1(new_n729), .A2(G116), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n747), .B2(new_n346), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n740), .A2(G68), .ZN(new_n1133));
  AOI211_X1 g0933(.A(G41), .B(new_n286), .C1(new_n733), .C2(G283), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n736), .A2(G77), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n742), .A2(G58), .ZN(new_n1136));
  AND4_X1   g0936(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n232), .B2(new_n726), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1132), .B(new_n1138), .C1(G97), .C2(new_n724), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1139), .A2(KEYINPUT58), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(KEYINPUT58), .ZN(new_n1141));
  AOI21_X1  g0941(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1140), .B(new_n1141), .C1(G50), .C2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G125), .A2(new_n729), .B1(new_n724), .B2(G132), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n937), .B2(new_n747), .C1(new_n785), .C2(new_n759), .ZN(new_n1145));
  INV_X1    g0945(.A(G128), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n726), .A2(new_n1146), .B1(new_n737), .B2(new_n1068), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT119), .Z(new_n1148));
  NOR2_X1   g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI211_X1 g0951(.A(G33), .B(G41), .C1(new_n733), .C2(G124), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n786), .B2(new_n743), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1143), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1130), .B1(new_n1155), .B2(new_n783), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n1107), .B2(new_n713), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1126), .B2(new_n700), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1128), .A2(new_n1160), .ZN(G375));
  NAND2_X1  g0961(.A1(new_n859), .A2(new_n713), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n702), .B1(G68), .B2(new_n804), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n278), .B1(new_n743), .B2(new_n230), .C1(new_n346), .C2(new_n759), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n725), .A2(new_n526), .B1(new_n760), .B2(new_n726), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(G294), .C2(new_n729), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n736), .A2(G97), .B1(new_n733), .B2(G303), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT123), .Z(new_n1168));
  OAI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(new_n232), .C2(new_n751), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT124), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G132), .A2(new_n729), .B1(new_n763), .B2(G137), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n725), .B2(new_n1068), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1172), .A2(KEYINPUT125), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(KEYINPUT125), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1136), .B(new_n286), .C1(new_n1146), .C2(new_n732), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n737), .A2(new_n786), .B1(new_n759), .B2(new_n202), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(G150), .C2(new_n746), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1173), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1170), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1163), .B1(new_n1179), .B2(new_n716), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1162), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1094), .B2(new_n700), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1095), .A2(new_n930), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1088), .A2(new_n1094), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(G381));
  NOR2_X1   g0986(.A1(G375), .A2(G378), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n957), .A2(new_n770), .A3(new_n985), .ZN(new_n1188));
  NOR4_X1   g0988(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1187), .A2(new_n933), .A3(new_n952), .A4(new_n1189), .ZN(G407));
  NAND3_X1  g0990(.A1(new_n1187), .A2(G213), .A3(new_n625), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(G407), .A2(G213), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT126), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT126), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(G407), .A2(new_n1191), .A3(new_n1194), .A4(G213), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(G409));
  AOI21_X1  g0996(.A(G390), .B1(new_n933), .B2(new_n952), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1188), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n770), .B1(new_n957), .B2(new_n985), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n933), .A2(new_n952), .A3(G390), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1198), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1201), .B1(new_n1198), .B2(new_n1202), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT61), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT127), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1088), .A2(new_n1094), .A3(KEYINPUT60), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1209), .A2(new_n645), .ZN(new_n1210));
  OAI21_X1  g1010(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1094), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1184), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1182), .ZN(new_n1214));
  AOI21_X1  g1014(.A(G384), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n810), .B(new_n1182), .C1(new_n1210), .C2(new_n1212), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1208), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1209), .A2(new_n645), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1184), .B2(new_n1211), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n810), .B1(new_n1219), .B2(new_n1182), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1213), .A2(G384), .A3(new_n1214), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(KEYINPUT127), .A3(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n625), .A2(G213), .A3(G2897), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1217), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1223), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1220), .A2(KEYINPUT127), .A3(new_n1221), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1099), .B1(new_n1128), .B2(new_n1160), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n625), .A2(G213), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1050), .A2(new_n1055), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1047), .B1(new_n1231), .B2(new_n1048), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1096), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n645), .A3(new_n1098), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1056), .A2(new_n1084), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1157), .B1(new_n1236), .B2(new_n701), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1102), .A2(new_n931), .A3(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1229), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1227), .B1(new_n1228), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1228), .A2(new_n1243), .A3(new_n1241), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT62), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1207), .B(new_n1242), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1102), .A2(new_n1239), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1103), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n646), .B1(new_n1102), .B2(new_n1121), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1159), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1247), .B(new_n1229), .C1(new_n1251), .C2(new_n1099), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1252), .A2(KEYINPUT62), .A3(new_n1243), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1206), .B1(new_n1246), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT63), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1252), .B2(new_n1243), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1252), .B2(new_n1227), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1244), .A2(KEYINPUT63), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1205), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1254), .A2(new_n1259), .ZN(G405));
  OAI211_X1 g1060(.A(new_n1220), .B(new_n1221), .C1(new_n1187), .C2(new_n1228), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1228), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1251), .A2(new_n1099), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1243), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1261), .A2(new_n1205), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1205), .B1(new_n1261), .B2(new_n1264), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(G402));
endmodule


