//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n590, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT65), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  AND2_X1   g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G101), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n463), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n469), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n477), .A2(KEYINPUT66), .A3(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n469), .A2(new_n472), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n480), .A2(new_n481), .B1(G124), .B2(new_n482), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT67), .Z(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n465), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G102), .ZN(new_n491));
  NAND2_X1  g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n460), .B2(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n491), .B1(new_n494), .B2(new_n472), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n472), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n460), .A2(KEYINPUT4), .A3(G138), .A4(new_n472), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n489), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n491), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n466), .A2(new_n468), .A3(G126), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(new_n492), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n502), .B1(new_n504), .B2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n505), .A2(KEYINPUT68), .A3(new_n498), .A4(new_n499), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n508), .A2(KEYINPUT6), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT69), .B(G651), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  INV_X1    g087(.A(new_n510), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n513), .A2(G75), .ZN(new_n514));
  OAI21_X1  g089(.A(G543), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT69), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT69), .A2(G651), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT6), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n509), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n510), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n515), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NOR2_X1   g106(.A1(new_n520), .A2(new_n524), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(KEYINPUT70), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(KEYINPUT70), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n525), .A2(new_n527), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n520), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n537), .A2(new_n540), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G64), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n538), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT71), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(new_n513), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(KEYINPUT72), .A3(new_n513), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n539), .A2(G90), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n532), .A2(G52), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n538), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n532), .A2(G43), .B1(new_n513), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n539), .A2(G81), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g146(.A(new_n571), .B(KEYINPUT73), .Z(G188));
  NAND2_X1  g147(.A1(new_n511), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  NAND2_X1  g149(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n573), .A2(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n532), .A2(G53), .A3(new_n575), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n528), .A2(G65), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n508), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n528), .A2(new_n518), .A3(G91), .A4(new_n519), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT75), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT75), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n511), .A2(new_n586), .A3(G91), .A4(new_n528), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n583), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n580), .A2(new_n588), .ZN(G299));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n544), .B(new_n590), .ZN(G286));
  NAND2_X1  g166(.A1(new_n532), .A2(G49), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n539), .A2(G87), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G288));
  NAND3_X1  g170(.A1(new_n511), .A2(G86), .A3(new_n528), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT78), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n538), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(new_n513), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT77), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n603), .A3(new_n513), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n532), .A2(G48), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n597), .A2(new_n605), .A3(new_n606), .ZN(G305));
  NAND2_X1  g182(.A1(new_n539), .A2(G85), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n532), .A2(G47), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n608), .B(new_n609), .C1(new_n510), .C2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(new_n528), .A2(G66), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n508), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n511), .A2(new_n528), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n539), .A2(KEYINPUT10), .A3(G92), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n614), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G54), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n573), .ZN(new_n622));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G171), .B2(new_n623), .ZN(G284));
  OAI21_X1  g200(.A(new_n624), .B1(G171), .B2(new_n623), .ZN(G321));
  INV_X1    g201(.A(G286), .ZN(new_n627));
  OR3_X1    g202(.A1(new_n627), .A2(KEYINPUT79), .A3(new_n623), .ZN(new_n628));
  OAI21_X1  g203(.A(KEYINPUT79), .B1(new_n627), .B2(new_n623), .ZN(new_n629));
  INV_X1    g204(.A(G299), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n628), .B(new_n629), .C1(G868), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT80), .Z(G297));
  XOR2_X1   g207(.A(new_n631), .B(KEYINPUT81), .Z(G280));
  OR2_X1    g208(.A1(new_n622), .A2(G559), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n573), .A2(new_n621), .ZN(new_n636));
  AOI211_X1 g211(.A(new_n614), .B(new_n636), .C1(new_n618), .C2(new_n619), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n635), .B1(G860), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g214(.A1(new_n564), .A2(new_n623), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n635), .B2(new_n623), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g217(.A1(new_n460), .A2(new_n490), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n482), .A2(G123), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n477), .A2(G135), .ZN(new_n649));
  NOR2_X1   g224(.A1(G99), .A2(G2105), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(new_n472), .B2(G111), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n646), .A2(G2100), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n647), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT83), .Z(G156));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XOR2_X1   g233(.A(G2443), .B(G2446), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT15), .B(G2435), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2438), .ZN(new_n664));
  XOR2_X1   g239(.A(G2427), .B(G2430), .Z(new_n665));
  INV_X1    g240(.A(KEYINPUT14), .ZN(new_n666));
  AOI22_X1  g241(.A1(new_n664), .A2(new_n665), .B1(KEYINPUT84), .B2(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(KEYINPUT84), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n667), .B(new_n668), .C1(new_n664), .C2(new_n665), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n662), .B(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(G14), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2067), .B(G2678), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(new_n677), .A3(KEYINPUT17), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT18), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2072), .B(G2078), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n680), .B(new_n681), .C1(new_n679), .C2(new_n675), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n681), .B2(new_n680), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n687), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n691), .A2(KEYINPUT20), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n693), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n695), .A2(new_n687), .A3(new_n690), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n694), .B(new_n696), .C1(KEYINPUT20), .C2(new_n691), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n697), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT85), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G19), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n565), .B2(new_n705), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G1341), .ZN(new_n708));
  NOR2_X1   g283(.A1(G27), .A2(G29), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G164), .B2(G29), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G2078), .ZN(new_n711));
  NAND2_X1  g286(.A1(G168), .A2(G16), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G16), .B2(G21), .ZN(new_n713));
  INV_X1    g288(.A(G1966), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT97), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n713), .A2(new_n714), .B1(G1341), .B2(new_n707), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G1961), .ZN(new_n719));
  NAND2_X1  g294(.A1(G171), .A2(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G5), .B2(G16), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n711), .B(new_n718), .C1(new_n719), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n705), .A2(G20), .ZN(new_n723));
  OAI211_X1 g298(.A(KEYINPUT23), .B(new_n723), .C1(new_n630), .C2(new_n705), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(KEYINPUT23), .B2(new_n723), .ZN(new_n725));
  INV_X1    g300(.A(G1956), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(KEYINPUT24), .A2(G34), .ZN(new_n729));
  NOR2_X1   g304(.A1(KEYINPUT24), .A2(G34), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n729), .A2(new_n730), .A3(G29), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n474), .B2(G29), .ZN(new_n732));
  INV_X1    g307(.A(G2084), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n652), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT30), .B(G28), .ZN(new_n738));
  OR2_X1    g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  NAND2_X1  g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n738), .A2(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n734), .A2(new_n735), .A3(new_n737), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n490), .A2(G103), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT94), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT25), .ZN(new_n746));
  NAND2_X1  g321(.A1(G115), .A2(G2104), .ZN(new_n747));
  INV_X1    g322(.A(G127), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n469), .B2(new_n748), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n749), .A2(G2105), .B1(new_n477), .B2(G139), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(KEYINPUT95), .B1(new_n746), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT25), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n745), .B(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT95), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n754), .A2(new_n755), .A3(new_n750), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n752), .A2(G29), .A3(new_n756), .ZN(new_n757));
  OR2_X1    g332(.A1(G29), .A2(G33), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n742), .B1(new_n760), .B2(G2072), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n736), .A2(G35), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n736), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G2090), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n761), .B(new_n766), .C1(G2072), .C2(new_n760), .ZN(new_n767));
  NOR2_X1   g342(.A1(G29), .A2(G32), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n477), .A2(G141), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT26), .Z(new_n773));
  AOI22_X1  g348(.A1(new_n482), .A2(G129), .B1(G105), .B2(new_n490), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n768), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT27), .B(G1996), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n765), .A2(G2090), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n767), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n721), .A2(new_n719), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT90), .B1(G4), .B2(G16), .ZN(new_n783));
  OR3_X1    g358(.A1(KEYINPUT90), .A2(G4), .A3(G16), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n783), .B(new_n784), .C1(new_n622), .C2(new_n705), .ZN(new_n785));
  INV_X1    g360(.A(G1348), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n736), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n482), .A2(KEYINPUT91), .A3(G128), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT91), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n460), .A2(G2105), .ZN(new_n792));
  INV_X1    g367(.A(G128), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n790), .A2(new_n794), .B1(G140), .B2(new_n477), .ZN(new_n795));
  OR2_X1    g370(.A1(G104), .A2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n796), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT92), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G29), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n800), .A2(KEYINPUT93), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(KEYINPUT93), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n789), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2067), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n782), .A2(new_n787), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n722), .A2(new_n728), .A3(new_n781), .A4(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G24), .B(G290), .S(G16), .Z(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT86), .Z(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(G1986), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(G1986), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n482), .A2(G119), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n477), .A2(G131), .ZN(new_n812));
  OR2_X1    g387(.A1(G95), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n813), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  MUX2_X1   g390(.A(G25), .B(new_n815), .S(G29), .Z(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT35), .B(G1991), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n810), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G305), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(new_n705), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G6), .B2(new_n705), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT32), .B(G1981), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT87), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n705), .A2(G22), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G166), .B2(new_n705), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n822), .A2(new_n824), .B1(G1971), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(G16), .A2(G23), .ZN(new_n829));
  OR2_X1    g404(.A1(G288), .A2(KEYINPUT88), .ZN(new_n830));
  NAND2_X1  g405(.A1(G288), .A2(KEYINPUT88), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n829), .B1(new_n832), .B2(G16), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT33), .B(G1976), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT89), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n827), .A2(G1971), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n825), .A2(new_n828), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AOI211_X1 g413(.A(new_n809), .B(new_n819), .C1(new_n838), .C2(KEYINPUT34), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n816), .A2(new_n817), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(KEYINPUT34), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT36), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n839), .A2(new_n844), .A3(new_n840), .A4(new_n841), .ZN(new_n845));
  AOI211_X1 g420(.A(new_n708), .B(new_n806), .C1(new_n843), .C2(new_n845), .ZN(G311));
  AOI21_X1  g421(.A(new_n806), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G1341), .B2(new_n707), .ZN(G150));
  NAND2_X1  g423(.A1(new_n532), .A2(G55), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT99), .B(G93), .ZN(new_n851));
  OAI221_X1 g426(.A(new_n849), .B1(new_n510), .B2(new_n850), .C1(new_n616), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n852), .B(new_n564), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT39), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n637), .A2(G559), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT38), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n856), .B(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n854), .B1(new_n859), .B2(G860), .ZN(G145));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n474), .B(new_n652), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n487), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n795), .A2(new_n798), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n775), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n799), .A2(new_n773), .A3(new_n771), .A4(new_n774), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n495), .A2(new_n500), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n865), .A2(new_n868), .A3(new_n866), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n746), .A2(KEYINPUT95), .A3(new_n751), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n755), .B1(new_n754), .B2(new_n750), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT100), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n752), .A2(new_n877), .A3(new_n756), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n871), .A3(new_n870), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n482), .A2(G130), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n477), .A2(G142), .ZN(new_n882));
  NOR2_X1   g457(.A1(G106), .A2(G2105), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(new_n472), .B2(G118), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(new_n644), .Z(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(new_n815), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n815), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(KEYINPUT101), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n876), .A2(new_n880), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT101), .B1(new_n887), .B2(new_n888), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n893), .A2(new_n876), .A3(new_n889), .A4(new_n880), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n863), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n861), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI211_X1 g472(.A(KEYINPUT102), .B(new_n863), .C1(new_n892), .C2(new_n894), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n892), .A2(new_n863), .A3(new_n894), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g477(.A1(new_n852), .A2(G868), .ZN(new_n903));
  XNOR2_X1  g478(.A(G303), .B(G290), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(new_n832), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n832), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(G305), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n820), .A3(new_n906), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n912), .A2(KEYINPUT103), .ZN(new_n913));
  INV_X1    g488(.A(new_n855), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n634), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n622), .A2(new_n630), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n637), .A2(G299), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n918), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(new_n915), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n912), .A2(KEYINPUT103), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n913), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n912), .A2(KEYINPUT103), .A3(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n903), .B1(new_n928), .B2(G868), .ZN(G295));
  AOI21_X1  g504(.A(new_n903), .B1(new_n928), .B2(G868), .ZN(G331));
  AND2_X1   g505(.A1(new_n910), .A2(KEYINPUT107), .ZN(new_n931));
  NAND2_X1  g506(.A1(G301), .A2(G168), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n552), .A2(new_n553), .B1(G52), .B2(new_n532), .ZN(new_n933));
  NAND3_X1  g508(.A1(G286), .A2(new_n933), .A3(new_n555), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n934), .A3(new_n855), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n855), .B1(new_n932), .B2(new_n934), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n920), .B(KEYINPUT105), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n932), .A2(new_n934), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n914), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n932), .A2(new_n934), .A3(KEYINPUT106), .A4(new_n855), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n940), .A2(new_n942), .A3(new_n918), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n935), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT105), .B1(new_n946), .B2(new_n920), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n931), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n920), .B1(new_n936), .B2(new_n937), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n910), .A2(KEYINPUT107), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n944), .A4(new_n938), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n948), .A2(new_n861), .A3(new_n953), .ZN(new_n954));
  XOR2_X1   g529(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n920), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n942), .A2(new_n960), .A3(new_n918), .A4(new_n935), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n942), .A2(new_n918), .A3(new_n935), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT108), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n910), .ZN(new_n965));
  INV_X1    g540(.A(new_n910), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n951), .A2(new_n966), .A3(new_n944), .A4(new_n938), .ZN(new_n967));
  INV_X1    g542(.A(new_n955), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n965), .A2(new_n861), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n956), .A2(new_n957), .A3(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n964), .A2(new_n910), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n967), .A2(new_n861), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT43), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n948), .A2(new_n953), .A3(new_n861), .A4(new_n968), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n957), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n970), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n495), .B2(new_n500), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n463), .A2(new_n473), .A3(G40), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  OR3_X1    g558(.A1(new_n983), .A2(G1986), .A3(G290), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(G1986), .A3(G290), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT109), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n775), .B(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n864), .B(G2067), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n983), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT110), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n815), .B(new_n817), .Z(new_n993));
  NOR2_X1   g568(.A1(new_n983), .A2(new_n993), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n987), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n981), .B1(new_n978), .B2(new_n979), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n501), .A2(new_n506), .A3(new_n977), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n997), .B2(new_n979), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G2078), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT121), .B(G1961), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n981), .B1(new_n997), .B2(KEYINPUT50), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n978), .A2(KEYINPUT50), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n997), .A2(new_n979), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT111), .ZN(new_n1009));
  INV_X1    g584(.A(G2078), .ZN(new_n1010));
  INV_X1    g585(.A(new_n981), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT45), .B(new_n977), .C1(new_n495), .C2(new_n500), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n997), .A2(new_n1015), .A3(new_n979), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1009), .A2(new_n1010), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  AOI211_X1 g592(.A(new_n1002), .B(new_n1007), .C1(new_n1017), .C2(new_n999), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1018), .A2(G301), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1005), .A2(new_n733), .A3(new_n1006), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n998), .A2(new_n714), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(G168), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n1023), .B2(G8), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT51), .B1(new_n1025), .B2(G168), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1023), .A2(G8), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT62), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1019), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  INV_X1    g606(.A(G1981), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n597), .A2(new_n605), .A3(new_n1032), .A4(new_n606), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n606), .A2(new_n602), .A3(new_n604), .ZN(new_n1034));
  INV_X1    g609(.A(new_n596), .ZN(new_n1035));
  OAI21_X1  g610(.A(G1981), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT49), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n978), .A2(new_n981), .ZN(new_n1040));
  INV_X1    g615(.A(G8), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1033), .A2(new_n1036), .A3(KEYINPUT49), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n832), .A2(G1976), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1042), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1046), .B1(new_n830), .B2(new_n831), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1042), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT52), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1009), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT112), .B(G1971), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1056), .A2(new_n1011), .A3(new_n1006), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT113), .B(G2090), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1053), .A2(new_n1055), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(new_n1041), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G303), .A2(G8), .ZN(new_n1062));
  XOR2_X1   g637(.A(new_n1062), .B(KEYINPUT55), .Z(new_n1063));
  AOI21_X1  g638(.A(new_n1052), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1063), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n978), .A2(KEYINPUT50), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1011), .B(new_n1066), .C1(new_n997), .C2(KEYINPUT50), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(new_n1058), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1065), .B1(new_n1069), .B2(new_n1041), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT123), .B1(new_n1064), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1005), .A2(new_n1059), .A3(new_n1006), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n997), .A2(new_n1015), .A3(new_n979), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1015), .B1(new_n997), .B2(new_n979), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1073), .A2(new_n1074), .A3(new_n1013), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1072), .B1(new_n1075), .B2(new_n1054), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(G8), .A3(new_n1063), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1044), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1070), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1030), .B(new_n1031), .C1(new_n1071), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G288), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1044), .A2(new_n1046), .A3(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1084), .A2(new_n1033), .ZN(new_n1085));
  OAI22_X1  g660(.A1(new_n1085), .A2(new_n1050), .B1(new_n1077), .B2(new_n1052), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1079), .A2(KEYINPUT63), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1025), .A2(new_n1041), .A3(G286), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1067), .A2(new_n726), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1091), .B(KEYINPUT118), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1090), .B1(new_n1053), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n630), .A2(KEYINPUT57), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n585), .A2(new_n587), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT116), .B1(new_n1096), .B2(new_n583), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n588), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n580), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(KEYINPUT117), .A3(new_n1101), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1094), .A2(new_n1095), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(new_n1095), .A3(new_n1105), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1075), .A2(new_n1092), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(new_n1090), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n637), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1040), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(G2067), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1056), .A2(new_n1011), .A3(new_n1006), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(new_n786), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT119), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n1116));
  AOI21_X1  g691(.A(G1348), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(new_n1112), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1106), .B1(new_n1110), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT120), .B(G1996), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT58), .B(G1341), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n1053), .A2(new_n1121), .B1(new_n1040), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n565), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT59), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1126), .A3(new_n565), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1114), .A2(KEYINPUT119), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1117), .A2(new_n1116), .A3(new_n1112), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT60), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1115), .A2(new_n1132), .A3(new_n1118), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(new_n637), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1119), .A2(KEYINPUT60), .A3(new_n622), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1128), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1106), .A2(new_n1109), .A3(KEYINPUT61), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT61), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1120), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1017), .A2(new_n999), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1007), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n996), .A2(new_n1012), .A3(new_n1000), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1143), .B(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(G171), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1018), .A2(G301), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1149), .A2(KEYINPUT54), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1141), .A2(G301), .A3(new_n1145), .A4(new_n1142), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1018), .B2(G301), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1028), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1152), .B(new_n1156), .C1(new_n1071), .C2(new_n1081), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1082), .B(new_n1089), .C1(new_n1140), .C2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT114), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1060), .B2(new_n1041), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1076), .A2(KEYINPUT114), .A3(G8), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1161), .A2(new_n1162), .A3(new_n1065), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT115), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n1078), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1163), .B2(new_n1078), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1077), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1159), .B1(new_n1168), .B2(new_n1088), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n995), .B1(new_n1158), .B2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n984), .B(KEYINPUT48), .Z(new_n1171));
  NOR3_X1   g746(.A1(new_n1171), .A2(new_n992), .A3(new_n994), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n983), .B1(new_n990), .B2(new_n776), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT126), .ZN(new_n1174));
  XOR2_X1   g749(.A(KEYINPUT125), .B(KEYINPUT46), .Z(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n983), .B2(G1996), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n982), .B(new_n988), .C1(new_n1177), .C2(KEYINPUT46), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1174), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1180));
  XNOR2_X1  g755(.A(new_n1179), .B(new_n1180), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n815), .A2(new_n817), .ZN(new_n1182));
  OAI22_X1  g757(.A1(new_n992), .A2(new_n1182), .B1(G2067), .B2(new_n799), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1172), .B(new_n1181), .C1(new_n1183), .C2(new_n982), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1170), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g760(.A1(G229), .A2(G401), .ZN(new_n1187));
  INV_X1    g761(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g762(.A(new_n1188), .B1(new_n899), .B2(new_n900), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n956), .A2(new_n969), .ZN(new_n1190));
  NOR2_X1   g764(.A1(G227), .A2(new_n458), .ZN(new_n1191));
  AND3_X1   g765(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(G308));
  NAND3_X1  g766(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(G225));
endmodule


