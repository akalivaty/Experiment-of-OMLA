//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT65), .Z(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n462), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(new_n466), .B2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n463), .A2(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n468), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(new_n462), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n462), .A2(G112), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n469), .A2(KEYINPUT67), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n469), .A2(KEYINPUT67), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n478), .B1(new_n481), .B2(G136), .ZN(G162));
  OAI211_X1 g057(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT68), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n462), .B2(G114), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n486), .A2(new_n488), .A3(new_n489), .A4(G2104), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT70), .ZN(new_n491));
  INV_X1    g066(.A(new_n469), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n460), .A2(G138), .A3(new_n462), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n492), .A2(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n484), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  AND2_X1   g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  OAI211_X1 g075(.A(G50), .B(G543), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n504), .A2(KEYINPUT71), .A3(G50), .A4(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(G75), .A2(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(new_n511), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(G88), .A3(new_n504), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n506), .A2(new_n514), .A3(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  OAI21_X1  g093(.A(G543), .B1(new_n499), .B2(new_n500), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n521), .B(G543), .C1(new_n499), .C2(new_n500), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n523), .A2(G51), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  AND3_X1   g103(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(G543), .B1(KEYINPUT72), .B2(KEYINPUT5), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n529), .A2(new_n530), .B1(new_n499), .B2(new_n500), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n525), .B(new_n527), .C1(new_n528), .C2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n524), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n523), .A2(G52), .ZN(new_n537));
  INV_X1    g112(.A(new_n531), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G90), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n529), .A2(new_n530), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n535), .B1(new_n545), .B2(KEYINPUT74), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n546), .B1(KEYINPUT74), .B2(new_n545), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n523), .A2(G43), .B1(G81), .B2(new_n538), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G860), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n543), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(new_n538), .B2(G91), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OR3_X1    g137(.A1(new_n519), .A2(KEYINPUT9), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n519), .B2(new_n562), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n567));
  NOR3_X1   g142(.A1(new_n524), .A2(new_n567), .A3(new_n532), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n532), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n523), .A2(G51), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT77), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G286));
  INV_X1    g150(.A(new_n519), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n515), .A2(G87), .A3(new_n504), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n538), .A2(G86), .B1(new_n576), .B2(G48), .ZN(new_n581));
  OAI21_X1  g156(.A(G61), .B1(new_n529), .B2(new_n530), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(KEYINPUT78), .B1(new_n584), .B2(G651), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  AOI211_X1 g161(.A(new_n586), .B(new_n535), .C1(new_n582), .C2(new_n583), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n581), .B1(new_n585), .B2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n543), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(new_n538), .B2(G85), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n523), .A2(G47), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n531), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n543), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n523), .A2(G54), .B1(new_n601), .B2(G651), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n595), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n595), .B1(new_n604), .B2(G868), .ZN(G321));
  AND2_X1   g181(.A1(new_n561), .A2(new_n565), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT79), .B1(new_n607), .B2(G868), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n574), .A2(new_n609), .ZN(new_n610));
  MUX2_X1   g185(.A(new_n608), .B(KEYINPUT79), .S(new_n610), .Z(G297));
  MUX2_X1   g186(.A(new_n608), .B(KEYINPUT79), .S(new_n610), .Z(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n604), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n549), .A2(new_n609), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n603), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n481), .A2(G135), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n474), .A2(G123), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n462), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT80), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(G2096), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(G2096), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n638), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G14), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n642), .A2(new_n645), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(G401));
  NOR2_X1   g224(.A1(G2072), .A2(G2078), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n442), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT17), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT83), .Z(new_n654));
  NOR2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n651), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2084), .B(G2090), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n655), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n651), .A2(new_n653), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n652), .A2(new_n654), .A3(new_n660), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n661), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2100), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT84), .B(G2096), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT85), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n673), .A2(KEYINPUT86), .A3(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT19), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n673), .A2(new_n674), .ZN(new_n683));
  INV_X1    g258(.A(new_n680), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(new_n675), .A3(new_n684), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n682), .B(new_n685), .C1(new_n684), .C2(new_n683), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1991), .B(G1996), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n686), .B(new_n687), .ZN(new_n692));
  INV_X1    g267(.A(new_n690), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n691), .A2(new_n694), .A3(new_n696), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  XOR2_X1   g276(.A(KEYINPUT93), .B(G28), .Z(new_n702));
  AOI21_X1  g277(.A(G29), .B1(new_n702), .B2(KEYINPUT30), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(KEYINPUT30), .B2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT31), .B(G11), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NOR2_X1   g282(.A1(G171), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G5), .B2(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(G1961), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(G21), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G168), .B2(new_n707), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n706), .B(new_n711), .C1(G1966), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(G1966), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT94), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n714), .B(new_n716), .C1(new_n717), .C2(new_n625), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT95), .Z(new_n719));
  NOR2_X1   g294(.A1(G29), .A2(G32), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n481), .A2(G141), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n474), .A2(G129), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT26), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n725), .A2(new_n726), .B1(G105), .B2(new_n464), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT92), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n720), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT27), .B(G1996), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n547), .A2(new_n548), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G16), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G16), .B2(G19), .ZN(new_n736));
  INV_X1    g311(.A(G1341), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n717), .B1(KEYINPUT24), .B2(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(KEYINPUT24), .B2(G34), .ZN(new_n740));
  INV_X1    g315(.A(G160), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT91), .B(G2084), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n717), .A2(G26), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT28), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n481), .A2(G140), .ZN(new_n747));
  OAI21_X1  g322(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n748));
  INV_X1    g323(.A(G116), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G2105), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n474), .B2(G128), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n746), .B1(new_n753), .B2(new_n717), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n738), .B(new_n744), .C1(G2067), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n707), .A2(G20), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT23), .Z(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1956), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n736), .B2(new_n737), .ZN(new_n760));
  OR3_X1    g335(.A1(new_n733), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(G164), .A2(G29), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G27), .B2(G29), .ZN(new_n763));
  INV_X1    g338(.A(G2078), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n710), .A2(new_n709), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n754), .A2(G2067), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n604), .A2(new_n707), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G4), .B2(new_n707), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT90), .B(G1348), .Z(new_n769));
  OAI211_X1 g344(.A(new_n765), .B(new_n766), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n717), .A2(G33), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT25), .Z(new_n773));
  AOI22_X1  g348(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n462), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n481), .B2(G139), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n771), .B1(new_n776), .B2(new_n717), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n768), .A2(new_n769), .B1(G2072), .B2(new_n777), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n778), .B1(G2072), .B2(new_n777), .C1(new_n764), .C2(new_n763), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n717), .A2(G35), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G162), .B2(new_n717), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT29), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2090), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n761), .A2(new_n770), .A3(new_n779), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n785));
  INV_X1    g360(.A(G305), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n786), .A2(new_n707), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G6), .B2(new_n707), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT32), .B(G1981), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G16), .A2(G23), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT88), .Z(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G288), .B2(new_n707), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT33), .ZN(new_n795));
  INV_X1    g370(.A(G1976), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n707), .A2(G22), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G166), .B2(new_n707), .ZN(new_n799));
  INV_X1    g374(.A(G1971), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n788), .A2(new_n790), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n791), .A2(new_n797), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(KEYINPUT34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n481), .A2(G131), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  INV_X1    g382(.A(G107), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G2105), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT87), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n811), .A2(new_n812), .B1(new_n474), .B2(G119), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G25), .B(new_n814), .S(G29), .Z(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n815), .B(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G24), .B(G290), .S(G16), .Z(new_n819));
  AOI22_X1  g394(.A1(new_n819), .A2(G1986), .B1(KEYINPUT89), .B2(KEYINPUT36), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G1986), .B2(new_n819), .ZN(new_n821));
  OR4_X1    g396(.A1(new_n804), .A2(new_n805), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n719), .B(new_n784), .C1(new_n785), .C2(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n822), .A2(new_n785), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(G311));
  INV_X1    g400(.A(G311), .ZN(G150));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n510), .B2(new_n511), .ZN(new_n828));
  NAND2_X1  g403(.A1(G80), .A2(G543), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT96), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n832), .B(new_n829), .C1(new_n543), .C2(new_n827), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n833), .A3(G651), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT98), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT97), .B(G55), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n521), .B1(new_n504), .B2(G543), .ZN(new_n837));
  INV_X1    g412(.A(new_n522), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n531), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n835), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n836), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n520), .B2(new_n522), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n845), .A2(KEYINPUT98), .A3(new_n841), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n834), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT99), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n849), .B(new_n834), .C1(new_n843), .C2(new_n846), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n734), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(KEYINPUT99), .A3(new_n549), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT38), .Z(new_n854));
  NOR2_X1   g429(.A1(new_n603), .A2(new_n613), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n857));
  AOI21_X1  g432(.A(G860), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n856), .ZN(new_n859));
  INV_X1    g434(.A(new_n834), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n839), .A2(new_n835), .A3(new_n842), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT98), .B1(new_n845), .B2(new_n841), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n550), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(new_n865), .ZN(G145));
  MUX2_X1   g441(.A(new_n729), .B(new_n730), .S(new_n776), .Z(new_n867));
  XNOR2_X1  g442(.A(G164), .B(new_n752), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n814), .B(new_n629), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n481), .A2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n474), .A2(G130), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n462), .A2(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n871), .B(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n867), .A2(new_n868), .ZN(new_n879));
  OR3_X1    g454(.A1(new_n870), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n878), .B1(new_n870), .B2(new_n879), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n624), .B(G160), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G162), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n880), .A2(new_n881), .A3(new_n885), .A4(new_n882), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g466(.A1(new_n847), .A2(new_n609), .ZN(new_n892));
  AOI21_X1  g467(.A(G288), .B1(new_n592), .B2(new_n593), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n592), .A2(G288), .A3(new_n593), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n897));
  NAND2_X1  g472(.A1(G303), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n506), .A2(KEYINPUT102), .A3(new_n514), .A4(new_n516), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n898), .A2(G305), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G305), .B1(new_n898), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n899), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n786), .ZN(new_n904));
  INV_X1    g479(.A(new_n895), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(new_n893), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n898), .A2(G305), .A3(new_n899), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n902), .A2(new_n908), .A3(KEYINPUT103), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT103), .B1(new_n902), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n902), .A2(new_n908), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(KEYINPUT42), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n912), .B1(KEYINPUT104), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(KEYINPUT104), .B2(new_n912), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n853), .B(new_n616), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n603), .A2(G299), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n607), .A2(new_n598), .A3(new_n602), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g495(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n920), .B2(KEYINPUT41), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n920), .B2(new_n917), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n916), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n892), .B1(new_n926), .B2(new_n609), .ZN(G295));
  OAI21_X1  g502(.A(new_n892), .B1(new_n926), .B2(new_n609), .ZN(G331));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n930));
  INV_X1    g505(.A(new_n920), .ZN(new_n931));
  OAI21_X1  g506(.A(G171), .B1(new_n568), .B2(new_n572), .ZN(new_n932));
  INV_X1    g507(.A(G168), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(G301), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n851), .A2(new_n935), .A3(new_n852), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n935), .B1(new_n851), .B2(new_n852), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n932), .A2(new_n934), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n850), .A2(new_n734), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n863), .A2(new_n849), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n852), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n851), .A2(new_n935), .A3(new_n852), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT41), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n920), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n944), .A2(new_n945), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n938), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n911), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n930), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI211_X1 g527(.A(KEYINPUT106), .B(new_n911), .C1(new_n938), .C2(new_n949), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n944), .A2(new_n923), .A3(new_n945), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT105), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n944), .A2(new_n923), .A3(new_n957), .A4(new_n945), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n956), .A2(new_n911), .A3(new_n938), .A4(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n959), .A2(new_n888), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n954), .A2(new_n960), .A3(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n888), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n938), .A2(new_n958), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n911), .B1(new_n964), .B2(new_n956), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n962), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n929), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n954), .A2(new_n960), .A3(new_n962), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT43), .B1(new_n963), .B2(new_n965), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT107), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n947), .A2(new_n948), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n936), .A2(new_n937), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n920), .B1(new_n944), .B2(new_n945), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n951), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT106), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n950), .A2(new_n930), .A3(new_n951), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n978), .A2(new_n962), .A3(new_n963), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n964), .A2(new_n956), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n951), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT43), .B1(new_n960), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT44), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n978), .A2(KEYINPUT43), .A3(new_n963), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n962), .B1(new_n960), .B2(new_n981), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n929), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n971), .A2(new_n988), .ZN(G397));
  INV_X1    g564(.A(G2067), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n752), .B(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT45), .B1(new_n497), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT108), .B(G40), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n463), .A2(new_n471), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n991), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n729), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n996), .B1(G1996), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n730), .B2(G1996), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n998), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n999), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n814), .B(new_n816), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n996), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n996), .ZN(new_n1007));
  XNOR2_X1  g582(.A(G290), .B(G1986), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n497), .A2(new_n992), .A3(new_n995), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(G8), .ZN(new_n1011));
  OR2_X1    g586(.A1(G305), .A2(G1981), .ZN(new_n1012));
  INV_X1    g587(.A(new_n581), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n535), .B1(new_n582), .B2(new_n583), .ZN(new_n1014));
  OAI21_X1  g589(.A(G1981), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(KEYINPUT49), .A3(new_n1015), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(G8), .A3(new_n1010), .A4(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G288), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(new_n796), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1011), .B1(new_n1022), .B2(new_n1012), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n497), .A2(new_n992), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n497), .A2(new_n1026), .A3(new_n992), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n995), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT110), .B1(new_n1028), .B2(G2090), .ZN(new_n1029));
  INV_X1    g604(.A(new_n995), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n993), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n800), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1030), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n1036));
  INV_X1    g611(.A(G2090), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1027), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1029), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G8), .ZN(new_n1040));
  INV_X1    g615(.A(G8), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G166), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1043), .A2(KEYINPUT111), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(KEYINPUT111), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1040), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1021), .A2(G1976), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT112), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(new_n1010), .A3(G8), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT52), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n796), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1051), .A2(new_n1010), .A3(G8), .A4(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1020), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT113), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1020), .A2(new_n1053), .A3(new_n1058), .A4(new_n1055), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1023), .B1(new_n1049), .B2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1062));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1033), .B2(G2078), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1024), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n995), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT114), .B1(new_n993), .B2(new_n1030), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1063), .A2(G2078), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1032), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1028), .A2(new_n710), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(KEYINPUT124), .A3(new_n1073), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1065), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(G301), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1071), .A2(G40), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n461), .A2(KEYINPUT125), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(new_n462), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n461), .A2(KEYINPUT125), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n471), .B(new_n1080), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1067), .A2(new_n1032), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1064), .A2(new_n1073), .A3(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1086), .A2(G171), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1062), .B1(new_n1079), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  INV_X1    g664(.A(G1956), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1028), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(G2072), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1031), .A2(new_n1032), .A3(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n607), .B(KEYINPUT57), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1091), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1089), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1095), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1091), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(KEYINPUT61), .A3(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT58), .B(G1341), .Z(new_n1104));
  NAND2_X1  g679(.A1(new_n1010), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1033), .B2(G1996), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n734), .A2(KEYINPUT119), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(KEYINPUT59), .A3(new_n1107), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1098), .A2(new_n1103), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1010), .A2(G2067), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n1028), .B2(new_n769), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT60), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT121), .B1(new_n1116), .B2(new_n603), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(KEYINPUT60), .A3(new_n603), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1115), .A2(new_n1122), .A3(new_n604), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1117), .A2(new_n1120), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1114), .A2(KEYINPUT60), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1112), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1114), .A2(new_n603), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1101), .B1(new_n1127), .B2(new_n1096), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1088), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1078), .A2(G301), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1086), .A2(G171), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(KEYINPUT54), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1028), .A2(G2090), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1971), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1134));
  OAI21_X1  g709(.A(G8), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1056), .B1(new_n1135), .B2(new_n1048), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1039), .A2(G8), .A3(new_n1047), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1069), .A2(new_n1032), .A3(new_n1070), .ZN(new_n1140));
  INV_X1    g715(.A(G1966), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1028), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT115), .B(G2084), .Z(new_n1143));
  AOI22_X1  g718(.A1(new_n1140), .A2(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1041), .B1(new_n1144), .B2(G168), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT122), .B(KEYINPUT51), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1144), .A2(new_n1041), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n933), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1151), .A2(KEYINPUT122), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1150), .B1(new_n1145), .B2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1132), .B(new_n1139), .C1(new_n1148), .C2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1061), .B1(new_n1129), .B2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1144), .A2(new_n1041), .A3(G286), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT116), .B1(new_n1138), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT116), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1156), .A2(new_n1136), .A3(new_n1160), .A4(new_n1137), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1156), .A2(KEYINPUT63), .A3(new_n1137), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1040), .A2(new_n1048), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1164), .A2(new_n1060), .A3(KEYINPUT117), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT117), .B1(new_n1164), .B2(new_n1060), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1163), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1162), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT62), .B1(new_n1153), .B2(new_n1148), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1145), .A2(new_n1152), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1170), .A2(new_n1171), .A3(new_n1147), .A4(new_n1150), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1138), .A2(new_n1078), .A3(G301), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1169), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1168), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1009), .B1(new_n1155), .B2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1004), .A2(new_n816), .A3(new_n806), .A4(new_n813), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n753), .A2(new_n990), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n996), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n996), .B1(new_n991), .B2(new_n1000), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT46), .B1(new_n996), .B2(G1996), .ZN(new_n1184));
  OR3_X1    g759(.A1(new_n996), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT47), .Z(new_n1187));
  NOR3_X1   g762(.A1(new_n996), .A2(G1986), .A3(G290), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT48), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1187), .B1(new_n1006), .B2(new_n1189), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1181), .A2(new_n1182), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1176), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g767(.A(new_n458), .B1(new_n647), .B2(new_n648), .ZN(new_n1194));
  OR2_X1    g768(.A1(G227), .A2(new_n1194), .ZN(new_n1195));
  AOI211_X1 g769(.A(KEYINPUT127), .B(new_n1195), .C1(new_n698), .C2(new_n699), .ZN(new_n1196));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n1197));
  INV_X1    g771(.A(new_n1195), .ZN(new_n1198));
  AOI21_X1  g772(.A(new_n1197), .B1(new_n700), .B2(new_n1198), .ZN(new_n1199));
  OAI221_X1 g773(.A(new_n890), .B1(new_n985), .B2(new_n984), .C1(new_n1196), .C2(new_n1199), .ZN(G225));
  INV_X1    g774(.A(G225), .ZN(G308));
endmodule


