//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n202), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  AND2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G141gat), .B(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(G155gat), .B2(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(G148gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G155gat), .B(G162gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT2), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n214), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225));
  XOR2_X1   g024(.A(G211gat), .B(G218gat), .Z(new_n226));
  AOI21_X1  g025(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n227));
  OR2_X1    g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT72), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(G197gat), .A2(G204gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(G197gat), .A2(G204gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT72), .B1(new_n235), .B2(new_n227), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n226), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n235), .A2(KEYINPUT72), .A3(new_n227), .ZN(new_n238));
  INV_X1    g037(.A(new_n226), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n225), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n224), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n203), .A2(new_n204), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n214), .A2(new_n223), .A3(new_n242), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n225), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n229), .ZN(new_n248));
  INV_X1    g047(.A(new_n227), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n231), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n239), .B1(new_n238), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n226), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n244), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(G22gat), .B1(new_n243), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n214), .A2(new_n223), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT29), .B1(new_n251), .B2(new_n252), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g057(.A(G22gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n237), .A2(new_n240), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n260), .A2(new_n246), .B1(new_n204), .B2(new_n203), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT31), .B(G50gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n255), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n255), .B2(new_n262), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n207), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n255), .A2(new_n262), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n263), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n255), .A2(new_n262), .A3(new_n264), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n206), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G227gat), .A2(G233gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n275));
  INV_X1    g074(.A(G183gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT27), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT27), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(G183gat), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n275), .B1(new_n281), .B2(KEYINPUT67), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n281), .A2(KEYINPUT66), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(KEYINPUT67), .ZN(new_n284));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n288));
  OR3_X1    g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n286), .B2(new_n287), .ZN(new_n290));
  INV_X1    g089(.A(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n289), .B(new_n290), .C1(KEYINPUT26), .C2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT67), .B1(new_n281), .B2(KEYINPUT66), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n275), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n284), .A2(new_n285), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(G134gat), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G127gat), .ZN(new_n302));
  OAI22_X1  g101(.A1(new_n298), .A2(KEYINPUT1), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G120gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G113gat), .ZN(new_n305));
  INV_X1    g104(.A(G113gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G120gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G127gat), .B(G134gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n303), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(G183gat), .B2(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316));
  INV_X1    g115(.A(new_n285), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(KEYINPUT65), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT65), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n285), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n315), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n293), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n324));
  NAND2_X1  g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(new_n326), .A3(KEYINPUT25), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n314), .B1(new_n316), .B2(new_n285), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n297), .A2(new_n312), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n312), .B1(new_n297), .B2(new_n332), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n274), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT32), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G15gat), .B(G43gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT69), .ZN(new_n340));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n336), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n281), .A2(KEYINPUT67), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT28), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n296), .B1(new_n295), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n294), .A2(new_n285), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n332), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n303), .A2(new_n311), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n297), .A2(new_n312), .A3(new_n332), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n273), .A3(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n352), .B(new_n354), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n342), .A2(KEYINPUT70), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n342), .A2(KEYINPUT70), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(KEYINPUT33), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n335), .A2(new_n358), .A3(KEYINPUT32), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n273), .B1(new_n350), .B2(new_n351), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT32), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n342), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n361), .A2(KEYINPUT33), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n359), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n352), .B(new_n353), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n272), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n348), .B2(new_n225), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n297), .B2(new_n332), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n260), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n348), .A2(new_n370), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n297), .B2(new_n332), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n374), .B(new_n253), .C1(new_n375), .C2(new_n370), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n373), .A2(new_n380), .A3(new_n376), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XOR2_X1   g184(.A(KEYINPUT73), .B(KEYINPUT30), .Z(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT74), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(KEYINPUT74), .A3(new_n386), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n312), .A2(new_n224), .A3(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n303), .A2(new_n214), .A3(new_n311), .A4(new_n223), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n395), .A3(KEYINPUT76), .ZN(new_n396));
  OR3_X1    g195(.A1(new_n394), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n220), .B1(new_n222), .B2(new_n219), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT3), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n349), .A3(new_n245), .ZN(new_n401));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(KEYINPUT5), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n396), .A2(new_n397), .A3(new_n401), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n392), .B1(new_n312), .B2(new_n224), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n402), .B(new_n401), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n349), .A2(new_n256), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n394), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n411), .B2(new_n403), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n408), .A2(KEYINPUT75), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT75), .B1(new_n408), .B2(new_n412), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n405), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G1gat), .B(G29gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT0), .ZN(new_n418));
  XNOR2_X1  g217(.A(G57gat), .B(G85gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n420), .B(new_n405), .C1(new_n414), .C2(new_n415), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n416), .A2(KEYINPUT6), .A3(new_n421), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT35), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n368), .A2(new_n391), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n405), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n412), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n429), .B1(new_n432), .B2(new_n413), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n423), .B1(new_n433), .B2(new_n420), .ZN(new_n434));
  INV_X1    g233(.A(new_n424), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT77), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT77), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n422), .A2(new_n437), .A3(new_n423), .A4(new_n424), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n438), .A3(new_n426), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(new_n391), .A3(new_n368), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT35), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n440), .B2(KEYINPUT35), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n428), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT37), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n373), .A2(new_n445), .A3(new_n376), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT79), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n373), .A2(KEYINPUT79), .A3(new_n376), .A4(new_n445), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n377), .A2(KEYINPUT37), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT81), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n381), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n445), .B1(new_n373), .B2(new_n376), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT81), .B1(new_n454), .B2(new_n380), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT38), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n425), .A2(new_n426), .A3(new_n384), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n454), .A2(KEYINPUT38), .A3(new_n380), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n450), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n450), .A2(new_n459), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT80), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n457), .A2(new_n458), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n396), .A2(new_n401), .A3(new_n397), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n403), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n410), .A2(new_n394), .A3(new_n402), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(KEYINPUT39), .A3(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n468), .B(new_n420), .C1(KEYINPUT39), .C2(new_n466), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n422), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n469), .A2(new_n470), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n389), .A2(new_n390), .ZN(new_n475));
  INV_X1    g274(.A(new_n385), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n272), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n464), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n439), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n272), .B1(new_n480), .B2(new_n477), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n367), .A2(KEYINPUT36), .A3(new_n360), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT36), .B1(new_n367), .B2(new_n360), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n444), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT83), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n444), .A2(new_n485), .A3(KEYINPUT83), .ZN(new_n489));
  NAND2_X1  g288(.A1(G229gat), .A2(G233gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT13), .ZN(new_n491));
  INV_X1    g290(.A(G8gat), .ZN(new_n492));
  INV_X1    g291(.A(G1gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT16), .ZN(new_n494));
  XOR2_X1   g293(.A(G15gat), .B(G22gat), .Z(new_n495));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT85), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n494), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n492), .B1(new_n500), .B2(KEYINPUT86), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n498), .B(KEYINPUT85), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(G1gat), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  OAI221_X1 g303(.A(new_n500), .B1(KEYINPUT86), .B2(new_n492), .C1(G1gat), .C2(new_n502), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G43gat), .B(G50gat), .Z(new_n508));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n512));
  INV_X1    g311(.A(G29gat), .ZN(new_n513));
  INV_X1    g312(.A(G36gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT14), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT14), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(G29gat), .A2(G36gat), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n510), .A2(new_n512), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(KEYINPUT15), .A3(new_n511), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n522), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n506), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n491), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n490), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT87), .B1(new_n523), .B2(KEYINPUT17), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT87), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n525), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI211_X1 g332(.A(KEYINPUT84), .B(KEYINPUT17), .C1(new_n520), .C2(new_n522), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT84), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n535), .B1(new_n525), .B2(new_n532), .ZN(new_n536));
  OAI22_X1  g335(.A1(new_n530), .A2(new_n533), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n526), .B(new_n529), .C1(new_n537), .C2(new_n506), .ZN(new_n538));
  INV_X1    g337(.A(new_n536), .ZN(new_n539));
  INV_X1    g338(.A(new_n534), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n523), .A2(KEYINPUT87), .A3(KEYINPUT17), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n531), .B1(new_n525), .B2(new_n532), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(new_n507), .A3(KEYINPUT88), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n528), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n527), .B1(new_n545), .B2(KEYINPUT18), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT18), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n545), .B2(KEYINPUT89), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT89), .ZN(new_n549));
  AOI211_X1 g348(.A(new_n549), .B(new_n528), .C1(new_n538), .C2(new_n544), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n546), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G197gat), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT11), .B(G169gat), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT12), .Z(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT90), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(new_n546), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  OAI221_X1 g359(.A(new_n546), .B1(new_n558), .B2(new_n557), .C1(new_n548), .C2(new_n550), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT94), .ZN(new_n564));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT7), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT93), .B1(new_n537), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT93), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n571), .B(new_n572), .Z(new_n576));
  NAND3_X1  g375(.A1(new_n543), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n576), .B2(new_n523), .ZN(new_n581));
  OAI211_X1 g380(.A(KEYINPUT95), .B(new_n564), .C1(new_n578), .C2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n581), .B1(new_n574), .B2(new_n577), .ZN(new_n584));
  INV_X1    g383(.A(new_n564), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G134gat), .B(G162gat), .Z(new_n587));
  NOR2_X1   g386(.A1(new_n579), .A2(KEYINPUT41), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n584), .B2(new_n585), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n582), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT96), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT96), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n582), .A2(new_n586), .A3(new_n590), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n584), .B(new_n585), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n589), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G57gat), .B(G64gat), .Z(new_n599));
  INV_X1    g398(.A(KEYINPUT9), .ZN(new_n600));
  INV_X1    g399(.A(G71gat), .ZN(new_n601));
  INV_X1    g400(.A(G78gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n599), .A2(KEYINPUT91), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G71gat), .B(G78gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n607));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  AOI21_X1  g408(.A(new_n506), .B1(KEYINPUT21), .B2(new_n606), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT92), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n611), .B(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n598), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n604), .B(new_n605), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n576), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n573), .A2(new_n606), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n573), .A2(new_n606), .A3(KEYINPUT10), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G230gat), .ZN(new_n627));
  INV_X1    g426(.A(G233gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n621), .A2(new_n623), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n632), .B2(new_n630), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n631), .B(new_n636), .C1(new_n632), .C2(new_n630), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(KEYINPUT97), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n633), .A2(new_n641), .A3(new_n637), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n619), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n488), .A2(new_n489), .A3(new_n562), .A4(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n439), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(new_n493), .ZN(G1324gat));
  XNOR2_X1  g448(.A(KEYINPUT16), .B(G8gat), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n647), .A2(new_n391), .A3(new_n650), .ZN(new_n651));
  OR3_X1    g450(.A1(new_n651), .A2(KEYINPUT98), .A3(KEYINPUT42), .ZN(new_n652));
  OAI21_X1  g451(.A(G8gat), .B1(new_n647), .B2(new_n391), .ZN(new_n653));
  OAI21_X1  g452(.A(KEYINPUT42), .B1(new_n651), .B2(KEYINPUT98), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(G1325gat));
  NOR3_X1   g454(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT99), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT36), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n365), .A2(new_n366), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n355), .B1(new_n359), .B2(new_n343), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n367), .A2(KEYINPUT36), .A3(new_n360), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G15gat), .B1(new_n647), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n367), .A2(new_n360), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(G15gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n647), .B2(new_n668), .ZN(G1326gat));
  INV_X1    g468(.A(new_n272), .ZN(new_n670));
  OR3_X1    g469(.A1(new_n647), .A2(KEYINPUT100), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT100), .B1(new_n647), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  INV_X1    g474(.A(new_n618), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n643), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n598), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n488), .A2(new_n489), .A3(new_n562), .A4(new_n679), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(G29gat), .A3(new_n439), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT45), .Z(new_n682));
  NAND4_X1  g481(.A1(new_n488), .A2(KEYINPUT44), .A3(new_n489), .A4(new_n598), .ZN(new_n683));
  INV_X1    g482(.A(new_n428), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n440), .A2(KEYINPUT35), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT82), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT35), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n664), .A2(new_n479), .A3(new_n481), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n598), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n562), .A2(new_n677), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G29gat), .B1(new_n695), .B2(new_n439), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n682), .A2(new_n696), .ZN(G1328gat));
  NOR3_X1   g496(.A1(new_n680), .A2(G36gat), .A3(new_n391), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT46), .ZN(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n695), .B2(new_n391), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1329gat));
  INV_X1    g500(.A(new_n664), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n683), .A2(new_n702), .A3(new_n692), .A4(new_n694), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G43gat), .ZN(new_n704));
  OR3_X1    g503(.A1(new_n680), .A2(G43gat), .A3(new_n667), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g506(.A(KEYINPUT48), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n683), .A2(new_n272), .A3(new_n692), .A4(new_n694), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G50gat), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n708), .B1(new_n710), .B2(KEYINPUT101), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n680), .A2(G50gat), .A3(new_n670), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(G50gat), .B2(new_n709), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n711), .B(new_n713), .ZN(G1331gat));
  NAND3_X1  g513(.A1(new_n664), .A2(new_n479), .A3(new_n481), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n444), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n562), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n716), .A2(new_n717), .A3(new_n619), .A4(new_n643), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT102), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(KEYINPUT102), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n439), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT103), .B(G57gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1332gat));
  XNOR2_X1  g523(.A(KEYINPUT105), .B(KEYINPUT106), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n719), .A2(new_n720), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n391), .A2(KEYINPUT104), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n391), .A2(KEYINPUT104), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n727), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n729), .B1(new_n727), .B2(new_n733), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n726), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n727), .A2(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n728), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n727), .A2(new_n729), .A3(new_n733), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n725), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n736), .A2(new_n740), .ZN(G1333gat));
  XNOR2_X1  g540(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G71gat), .B1(new_n721), .B2(new_n664), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n721), .A2(G71gat), .A3(new_n667), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n746), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(new_n744), .A3(new_n742), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(G1334gat));
  NOR2_X1   g549(.A1(new_n721), .A2(new_n670), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(new_n602), .ZN(G1335gat));
  NOR2_X1   g551(.A1(new_n562), .A2(new_n676), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n592), .A2(new_n594), .B1(new_n596), .B2(new_n589), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n444), .B2(new_n715), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n754), .B1(new_n756), .B2(KEYINPUT108), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n690), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n762), .A2(new_n568), .A3(new_n480), .A4(new_n643), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n754), .A2(new_n644), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n693), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765), .B2(new_n439), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(G1336gat));
  NOR3_X1   g566(.A1(new_n732), .A2(G92gat), .A3(new_n644), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  INV_X1    g569(.A(new_n732), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n693), .A2(new_n771), .A3(new_n764), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G92gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775));
  OAI211_X1 g574(.A(KEYINPUT108), .B(new_n598), .C1(new_n688), .C2(new_n689), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n753), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT108), .B1(new_n716), .B2(new_n598), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n761), .A2(KEYINPUT109), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(new_n757), .B2(new_n759), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n768), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n683), .A2(new_n477), .A3(new_n692), .A4(new_n764), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G92gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n775), .B1(new_n786), .B2(KEYINPUT52), .ZN(new_n787));
  AOI211_X1 g586(.A(KEYINPUT110), .B(new_n770), .C1(new_n783), .C2(new_n785), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n774), .B1(new_n787), .B2(new_n788), .ZN(G1337gat));
  XOR2_X1   g588(.A(KEYINPUT111), .B(G99gat), .Z(new_n790));
  NAND4_X1  g589(.A1(new_n762), .A2(new_n666), .A3(new_n643), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n765), .A2(new_n664), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n790), .ZN(G1338gat));
  NAND3_X1  g592(.A1(new_n693), .A2(new_n272), .A3(new_n764), .ZN(new_n794));
  XNOR2_X1  g593(.A(KEYINPUT112), .B(G106gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n644), .A2(G106gat), .A3(new_n670), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n762), .A2(new_n799), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n781), .A2(new_n782), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n801), .A2(new_n799), .B1(new_n794), .B2(new_n795), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n798), .A2(new_n800), .B1(new_n802), .B2(new_n797), .ZN(G1339gat));
  INV_X1    g602(.A(new_n368), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n631), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n629), .B1(new_n624), .B2(new_n625), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n636), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n807), .A2(KEYINPUT55), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT55), .B1(new_n807), .B2(new_n810), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI211_X1 g613(.A(KEYINPUT113), .B(KEYINPUT55), .C1(new_n807), .C2(new_n810), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n639), .B(new_n811), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n562), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n538), .A2(new_n528), .A3(new_n544), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n538), .A2(KEYINPUT114), .A3(new_n528), .A4(new_n544), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n524), .A2(new_n526), .A3(new_n491), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n555), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n546), .B(new_n557), .C1(new_n548), .C2(new_n550), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n824), .A2(KEYINPUT115), .A3(new_n555), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n827), .A2(new_n643), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n598), .B1(new_n818), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n755), .A2(new_n832), .A3(new_n816), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n805), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  AND4_X1   g633(.A1(new_n643), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n816), .B1(new_n561), .B2(new_n560), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n755), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n832), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n598), .A3(new_n817), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(KEYINPUT116), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n834), .A2(new_n840), .A3(new_n618), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n619), .A2(new_n717), .A3(new_n644), .ZN(new_n842));
  AOI211_X1 g641(.A(new_n439), .B(new_n804), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n732), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n306), .A3(new_n562), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n272), .B1(new_n841), .B2(new_n842), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n771), .A2(new_n439), .A3(new_n667), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n562), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n846), .B1(new_n851), .B2(G113gat), .ZN(new_n852));
  AOI211_X1 g651(.A(KEYINPUT117), .B(new_n306), .C1(new_n850), .C2(new_n562), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n845), .B1(new_n852), .B2(new_n853), .ZN(G1340gat));
  NOR3_X1   g653(.A1(new_n849), .A2(new_n304), .A3(new_n644), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n844), .A2(new_n643), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n304), .ZN(G1341gat));
  NAND3_X1  g656(.A1(new_n844), .A2(new_n299), .A3(new_n676), .ZN(new_n858));
  OAI21_X1  g657(.A(G127gat), .B1(new_n849), .B2(new_n618), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1342gat));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n301), .A3(new_n391), .A4(new_n598), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n849), .B2(new_n755), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  NAND2_X1  g664(.A1(new_n841), .A2(new_n842), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n272), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n732), .A2(new_n664), .A3(new_n480), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n811), .A2(new_n639), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n812), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n562), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n830), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n755), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n676), .B1(new_n874), .B2(new_n839), .ZN(new_n875));
  INV_X1    g674(.A(new_n842), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n272), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n869), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n868), .A2(new_n878), .A3(new_n562), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G141gat), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n664), .A2(new_n272), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT118), .Z(new_n884));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n480), .A3(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n717), .A2(G141gat), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n866), .A2(KEYINPUT119), .A3(new_n480), .A4(new_n884), .ZN(new_n889));
  AND4_X1   g688(.A1(new_n732), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n732), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(G141gat), .B2(new_n879), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n882), .A2(new_n890), .B1(new_n893), .B2(new_n881), .ZN(G1344gat));
  NOR2_X1   g693(.A1(new_n644), .A2(G148gat), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n887), .A2(new_n732), .A3(new_n889), .A4(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n868), .A2(new_n878), .ZN(new_n897));
  AOI211_X1 g696(.A(KEYINPUT59), .B(new_n217), .C1(new_n897), .C2(new_n643), .ZN(new_n898));
  XNOR2_X1  g697(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT121), .B1(new_n875), .B2(new_n876), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n598), .B1(new_n872), .B2(new_n830), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n618), .B1(new_n901), .B2(new_n833), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n903), .A3(new_n842), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n670), .A2(KEYINPUT57), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n900), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n869), .A2(new_n644), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n670), .B1(new_n841), .B2(new_n842), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n906), .B(new_n907), .C1(new_n867), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n899), .B1(new_n909), .B2(G148gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n896), .B1(new_n898), .B2(new_n910), .ZN(G1345gat));
  NAND2_X1  g710(.A1(new_n897), .A2(new_n676), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G155gat), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n618), .A2(G155gat), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n887), .A2(new_n732), .A3(new_n889), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1346gat));
  NAND3_X1  g715(.A1(new_n868), .A2(new_n878), .A3(new_n598), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G162gat), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n755), .A2(G162gat), .A3(new_n477), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n887), .A2(new_n889), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n918), .A2(new_n920), .A3(KEYINPUT122), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n480), .A2(new_n391), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n667), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n847), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(new_n291), .A3(new_n717), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n480), .B1(new_n841), .B2(new_n842), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n732), .A2(new_n804), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n562), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n930), .B1(new_n291), .B2(new_n935), .ZN(G1348gat));
  OAI21_X1  g735(.A(G176gat), .B1(new_n929), .B2(new_n644), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n643), .A2(new_n292), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n933), .B2(new_n938), .ZN(G1349gat));
  NAND3_X1  g738(.A1(new_n676), .A2(new_n277), .A3(new_n279), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n933), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(G183gat), .B1(new_n929), .B2(new_n618), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n934), .A2(new_n280), .A3(new_n598), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n847), .A2(new_n598), .A3(new_n928), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n946), .A2(new_n947), .A3(G190gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n946), .B2(G190gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  OAI21_X1  g749(.A(new_n906), .B1(new_n908), .B2(new_n867), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT124), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n906), .B(new_n953), .C1(new_n908), .C2(new_n867), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n702), .A2(new_n927), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n952), .A2(new_n562), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  XOR2_X1   g755(.A(KEYINPUT123), .B(G197gat), .Z(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n883), .A2(new_n732), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n931), .A2(new_n562), .A3(new_n957), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(G1352gat));
  NAND4_X1  g761(.A1(new_n952), .A2(new_n643), .A3(new_n954), .A4(new_n955), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G204gat), .ZN(new_n964));
  AOI211_X1 g763(.A(G204gat), .B(new_n644), .C1(KEYINPUT125), .C2(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n931), .A2(new_n960), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n964), .A2(new_n968), .ZN(G1353gat));
  NOR2_X1   g768(.A1(new_n618), .A2(G211gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n931), .A2(new_n960), .A3(new_n970), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n971), .B(KEYINPUT126), .Z(new_n972));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n676), .ZN(new_n973));
  OAI21_X1  g772(.A(G211gat), .B1(new_n951), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT63), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT63), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n976), .B(G211gat), .C1(new_n951), .C2(new_n973), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n972), .A2(new_n975), .A3(new_n977), .ZN(G1354gat));
  INV_X1    g777(.A(G218gat), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n755), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n952), .A2(new_n954), .A3(new_n955), .A4(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n931), .A2(new_n598), .A3(new_n960), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(new_n979), .ZN(new_n983));
  OR2_X1    g782(.A1(new_n983), .A2(KEYINPUT127), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(KEYINPUT127), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(G1355gat));
endmodule


