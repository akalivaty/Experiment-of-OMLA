

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U555 ( .A(n774), .B(KEYINPUT100), .Z(n521) );
  INV_X1 U556 ( .A(n739), .ZN(n716) );
  AND2_X1 U557 ( .A1(G160), .A2(G40), .ZN(n694) );
  NAND2_X1 U558 ( .A1(n775), .A2(n521), .ZN(n776) );
  NOR2_X1 U559 ( .A1(G651), .A2(n631), .ZN(n654) );
  INV_X1 U560 ( .A(G2105), .ZN(n529) );
  AND2_X1 U561 ( .A1(n529), .A2(G2104), .ZN(n874) );
  NAND2_X1 U562 ( .A1(G101), .A2(n874), .ZN(n522) );
  XNOR2_X1 U563 ( .A(n522), .B(KEYINPUT23), .ZN(n523) );
  XNOR2_X1 U564 ( .A(KEYINPUT65), .B(n523), .ZN(n527) );
  NAND2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  XOR2_X2 U566 ( .A(KEYINPUT66), .B(n524), .Z(n879) );
  NAND2_X1 U567 ( .A1(n879), .A2(G113), .ZN(n525) );
  XOR2_X1 U568 ( .A(KEYINPUT67), .B(n525), .Z(n526) );
  NAND2_X1 U569 ( .A1(n527), .A2(n526), .ZN(n533) );
  NOR2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XOR2_X1 U571 ( .A(KEYINPUT17), .B(n528), .Z(n872) );
  NAND2_X1 U572 ( .A1(G137), .A2(n872), .ZN(n531) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n529), .ZN(n878) );
  NAND2_X1 U574 ( .A1(G125), .A2(n878), .ZN(n530) );
  NAND2_X1 U575 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X2 U576 ( .A1(n533), .A2(n532), .ZN(G160) );
  XOR2_X1 U577 ( .A(G2443), .B(G2446), .Z(n535) );
  XNOR2_X1 U578 ( .A(G2427), .B(G2451), .ZN(n534) );
  XNOR2_X1 U579 ( .A(n535), .B(n534), .ZN(n541) );
  XOR2_X1 U580 ( .A(G2430), .B(G2454), .Z(n537) );
  XNOR2_X1 U581 ( .A(G1341), .B(G1348), .ZN(n536) );
  XNOR2_X1 U582 ( .A(n537), .B(n536), .ZN(n539) );
  XOR2_X1 U583 ( .A(G2435), .B(G2438), .Z(n538) );
  XNOR2_X1 U584 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U585 ( .A(n541), .B(n540), .Z(n542) );
  AND2_X1 U586 ( .A1(G14), .A2(n542), .ZN(G401) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n631) );
  NAND2_X1 U588 ( .A1(n654), .A2(G52), .ZN(n546) );
  INV_X1 U589 ( .A(G651), .ZN(n547) );
  NOR2_X1 U590 ( .A1(G543), .A2(n547), .ZN(n543) );
  XOR2_X1 U591 ( .A(KEYINPUT68), .B(n543), .Z(n544) );
  XNOR2_X1 U592 ( .A(KEYINPUT1), .B(n544), .ZN(n647) );
  NAND2_X1 U593 ( .A1(G64), .A2(n647), .ZN(n545) );
  NAND2_X1 U594 ( .A1(n546), .A2(n545), .ZN(n552) );
  NOR2_X1 U595 ( .A1(n631), .A2(n547), .ZN(n650) );
  NAND2_X1 U596 ( .A1(G77), .A2(n650), .ZN(n549) );
  NOR2_X1 U597 ( .A1(G651), .A2(G543), .ZN(n646) );
  NAND2_X1 U598 ( .A1(G90), .A2(n646), .ZN(n548) );
  NAND2_X1 U599 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n550), .Z(n551) );
  NOR2_X1 U601 ( .A1(n552), .A2(n551), .ZN(G171) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U603 ( .A(G132), .ZN(G219) );
  INV_X1 U604 ( .A(G82), .ZN(G220) );
  INV_X1 U605 ( .A(G120), .ZN(G236) );
  INV_X1 U606 ( .A(G69), .ZN(G235) );
  INV_X1 U607 ( .A(G108), .ZN(G238) );
  NAND2_X1 U608 ( .A1(G63), .A2(n647), .ZN(n553) );
  XOR2_X1 U609 ( .A(KEYINPUT75), .B(n553), .Z(n555) );
  NAND2_X1 U610 ( .A1(n654), .A2(G51), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U612 ( .A(KEYINPUT6), .B(n556), .ZN(n563) );
  NAND2_X1 U613 ( .A1(n650), .A2(G76), .ZN(n557) );
  XNOR2_X1 U614 ( .A(KEYINPUT74), .B(n557), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n646), .A2(G89), .ZN(n558) );
  XNOR2_X1 U616 ( .A(KEYINPUT4), .B(n558), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U618 ( .A(n561), .B(KEYINPUT5), .Z(n562) );
  NOR2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U620 ( .A(KEYINPUT7), .B(n564), .Z(n565) );
  XNOR2_X1 U621 ( .A(KEYINPUT76), .B(n565), .ZN(G168) );
  XOR2_X1 U622 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U624 ( .A(n566), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U625 ( .A(G223), .ZN(n827) );
  NAND2_X1 U626 ( .A1(n827), .A2(G567), .ZN(n567) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  NAND2_X1 U628 ( .A1(G56), .A2(n647), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT14), .B(n568), .Z(n576) );
  NAND2_X1 U630 ( .A1(n646), .A2(G81), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT12), .B(n569), .Z(n572) );
  NAND2_X1 U632 ( .A1(n650), .A2(G68), .ZN(n570) );
  XOR2_X1 U633 ( .A(n570), .B(KEYINPUT70), .Z(n571) );
  NOR2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT71), .B(n573), .Z(n574) );
  XNOR2_X1 U636 ( .A(n574), .B(KEYINPUT13), .ZN(n575) );
  NOR2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U638 ( .A1(n654), .A2(G43), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n912) );
  INV_X1 U640 ( .A(G860), .ZN(n601) );
  OR2_X1 U641 ( .A1(n912), .A2(n601), .ZN(G153) );
  INV_X1 U642 ( .A(G171), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U644 ( .A1(n647), .A2(G66), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n579), .B(KEYINPUT72), .ZN(n586) );
  NAND2_X1 U646 ( .A1(G79), .A2(n650), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G92), .A2(n646), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G54), .A2(n654), .ZN(n582) );
  XNOR2_X1 U650 ( .A(KEYINPUT73), .B(n582), .ZN(n583) );
  NOR2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U653 ( .A(KEYINPUT15), .B(n587), .Z(n931) );
  INV_X1 U654 ( .A(G868), .ZN(n604) );
  NAND2_X1 U655 ( .A1(n931), .A2(n604), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U657 ( .A1(G78), .A2(n650), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G91), .A2(n646), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U660 ( .A1(G65), .A2(n647), .ZN(n592) );
  XNOR2_X1 U661 ( .A(KEYINPUT69), .B(n592), .ZN(n593) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n654), .A2(G53), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n596), .A2(n595), .ZN(G299) );
  NOR2_X1 U665 ( .A1(G286), .A2(n604), .ZN(n597) );
  XOR2_X1 U666 ( .A(KEYINPUT77), .B(n597), .Z(n600) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n598) );
  XNOR2_X1 U668 ( .A(KEYINPUT78), .B(n598), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n601), .A2(G559), .ZN(n602) );
  INV_X1 U671 ( .A(n931), .ZN(n899) );
  NAND2_X1 U672 ( .A1(n602), .A2(n899), .ZN(n603) );
  XNOR2_X1 U673 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(G559), .A2(n604), .ZN(n605) );
  NAND2_X1 U675 ( .A1(n899), .A2(n605), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n606), .B(KEYINPUT79), .ZN(n608) );
  NOR2_X1 U677 ( .A1(n912), .A2(G868), .ZN(n607) );
  NOR2_X1 U678 ( .A1(n608), .A2(n607), .ZN(G282) );
  XNOR2_X1 U679 ( .A(G2100), .B(KEYINPUT81), .ZN(n618) );
  NAND2_X1 U680 ( .A1(G123), .A2(n878), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n609), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G99), .A2(n874), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT80), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U685 ( .A1(G135), .A2(n872), .ZN(n614) );
  NAND2_X1 U686 ( .A1(G111), .A2(n879), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n988) );
  XNOR2_X1 U689 ( .A(n988), .B(G2096), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U691 ( .A1(n899), .A2(G559), .ZN(n667) );
  XNOR2_X1 U692 ( .A(n912), .B(n667), .ZN(n619) );
  NOR2_X1 U693 ( .A1(n619), .A2(G860), .ZN(n626) );
  NAND2_X1 U694 ( .A1(n654), .A2(G55), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G67), .A2(n647), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G80), .A2(n650), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G93), .A2(n646), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n660) );
  XNOR2_X1 U701 ( .A(n626), .B(n660), .ZN(G145) );
  NAND2_X1 U702 ( .A1(G49), .A2(n654), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U705 ( .A(KEYINPUT82), .B(n629), .ZN(n630) );
  NOR2_X1 U706 ( .A1(n647), .A2(n630), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n631), .A2(G87), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(G288) );
  AND2_X1 U709 ( .A1(G60), .A2(n647), .ZN(n637) );
  NAND2_X1 U710 ( .A1(G72), .A2(n650), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G85), .A2(n646), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n654), .A2(G47), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(G290) );
  NAND2_X1 U716 ( .A1(G75), .A2(n650), .ZN(n641) );
  NAND2_X1 U717 ( .A1(G88), .A2(n646), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n654), .A2(G50), .ZN(n643) );
  NAND2_X1 U720 ( .A1(G62), .A2(n647), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U722 ( .A1(n645), .A2(n644), .ZN(G166) );
  NAND2_X1 U723 ( .A1(n646), .A2(G86), .ZN(n649) );
  NAND2_X1 U724 ( .A1(G61), .A2(n647), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n650), .A2(G73), .ZN(n651) );
  XOR2_X1 U727 ( .A(KEYINPUT2), .B(n651), .Z(n652) );
  NOR2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n654), .A2(G48), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n656), .A2(n655), .ZN(G305) );
  NOR2_X1 U731 ( .A1(G868), .A2(n660), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n657), .B(KEYINPUT85), .ZN(n670) );
  XOR2_X1 U733 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n658) );
  XNOR2_X1 U734 ( .A(G288), .B(n658), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n660), .B(n659), .ZN(n662) );
  XNOR2_X1 U736 ( .A(G290), .B(G166), .ZN(n661) );
  XNOR2_X1 U737 ( .A(n662), .B(n661), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n912), .B(G299), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(G305), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n665), .B(n664), .ZN(n902) );
  XOR2_X1 U741 ( .A(n902), .B(KEYINPUT84), .Z(n666) );
  XNOR2_X1 U742 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U743 ( .A1(G868), .A2(n668), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n672), .ZN(n674) );
  XNOR2_X1 U748 ( .A(KEYINPUT86), .B(KEYINPUT21), .ZN(n673) );
  XNOR2_X1 U749 ( .A(n674), .B(n673), .ZN(n675) );
  NAND2_X1 U750 ( .A1(G2072), .A2(n675), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U752 ( .A1(G235), .A2(G236), .ZN(n676) );
  XOR2_X1 U753 ( .A(KEYINPUT88), .B(n676), .Z(n677) );
  NOR2_X1 U754 ( .A1(G238), .A2(n677), .ZN(n678) );
  NAND2_X1 U755 ( .A1(G57), .A2(n678), .ZN(n833) );
  NAND2_X1 U756 ( .A1(G567), .A2(n833), .ZN(n679) );
  XNOR2_X1 U757 ( .A(n679), .B(KEYINPUT89), .ZN(n685) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n680) );
  XNOR2_X1 U759 ( .A(KEYINPUT22), .B(n680), .ZN(n681) );
  NAND2_X1 U760 ( .A1(n681), .A2(G96), .ZN(n682) );
  NOR2_X1 U761 ( .A1(G218), .A2(n682), .ZN(n683) );
  XNOR2_X1 U762 ( .A(KEYINPUT87), .B(n683), .ZN(n834) );
  AND2_X1 U763 ( .A1(G2106), .A2(n834), .ZN(n684) );
  NOR2_X1 U764 ( .A1(n685), .A2(n684), .ZN(G319) );
  INV_X1 U765 ( .A(G319), .ZN(n687) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U767 ( .A1(n687), .A2(n686), .ZN(n832) );
  NAND2_X1 U768 ( .A1(n832), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(G102), .A2(n874), .ZN(n689) );
  NAND2_X1 U770 ( .A1(G138), .A2(n872), .ZN(n688) );
  NAND2_X1 U771 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U772 ( .A1(n878), .A2(G126), .ZN(n691) );
  NAND2_X1 U773 ( .A1(G114), .A2(n879), .ZN(n690) );
  NAND2_X1 U774 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U775 ( .A1(n693), .A2(n692), .ZN(G164) );
  INV_X1 U776 ( .A(G166), .ZN(G303) );
  NOR2_X1 U777 ( .A1(G164), .A2(G1384), .ZN(n758) );
  NAND2_X1 U778 ( .A1(n758), .A2(n694), .ZN(n739) );
  NAND2_X1 U779 ( .A1(G1348), .A2(n739), .ZN(n696) );
  NAND2_X1 U780 ( .A1(G2067), .A2(n716), .ZN(n695) );
  NAND2_X1 U781 ( .A1(n696), .A2(n695), .ZN(n703) );
  NOR2_X1 U782 ( .A1(n931), .A2(n703), .ZN(n702) );
  INV_X1 U783 ( .A(G1996), .ZN(n940) );
  NOR2_X1 U784 ( .A1(n739), .A2(n940), .ZN(n697) );
  XOR2_X1 U785 ( .A(n697), .B(KEYINPUT26), .Z(n699) );
  NAND2_X1 U786 ( .A1(n739), .A2(G1341), .ZN(n698) );
  NAND2_X1 U787 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U788 ( .A1(n700), .A2(n912), .ZN(n701) );
  NOR2_X1 U789 ( .A1(n702), .A2(n701), .ZN(n705) );
  AND2_X1 U790 ( .A1(n931), .A2(n703), .ZN(n704) );
  NOR2_X1 U791 ( .A1(n705), .A2(n704), .ZN(n710) );
  NAND2_X1 U792 ( .A1(n716), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U793 ( .A(KEYINPUT27), .B(n706), .ZN(n708) );
  AND2_X1 U794 ( .A1(G1956), .A2(n739), .ZN(n707) );
  OR2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n711) );
  NOR2_X1 U796 ( .A1(G299), .A2(n711), .ZN(n709) );
  NOR2_X1 U797 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U798 ( .A1(G299), .A2(n711), .ZN(n712) );
  XOR2_X1 U799 ( .A(n712), .B(KEYINPUT28), .Z(n713) );
  NOR2_X1 U800 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U801 ( .A(n715), .B(KEYINPUT29), .ZN(n721) );
  XOR2_X1 U802 ( .A(G2078), .B(KEYINPUT25), .Z(n948) );
  NOR2_X1 U803 ( .A1(n948), .A2(n739), .ZN(n718) );
  NOR2_X1 U804 ( .A1(n716), .A2(G1961), .ZN(n717) );
  NOR2_X1 U805 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U806 ( .A(KEYINPUT97), .B(n719), .ZN(n725) );
  NAND2_X1 U807 ( .A1(G171), .A2(n725), .ZN(n720) );
  NAND2_X1 U808 ( .A1(n721), .A2(n720), .ZN(n735) );
  NAND2_X1 U809 ( .A1(G8), .A2(n739), .ZN(n784) );
  NOR2_X1 U810 ( .A1(G1966), .A2(n784), .ZN(n729) );
  NOR2_X1 U811 ( .A1(G2084), .A2(n739), .ZN(n731) );
  NOR2_X1 U812 ( .A1(n729), .A2(n731), .ZN(n722) );
  NAND2_X1 U813 ( .A1(G8), .A2(n722), .ZN(n723) );
  XNOR2_X1 U814 ( .A(KEYINPUT30), .B(n723), .ZN(n724) );
  NOR2_X1 U815 ( .A1(G168), .A2(n724), .ZN(n727) );
  NOR2_X1 U816 ( .A1(G171), .A2(n725), .ZN(n726) );
  NOR2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U818 ( .A(KEYINPUT31), .B(n728), .Z(n736) );
  AND2_X1 U819 ( .A1(n735), .A2(n736), .ZN(n730) );
  NOR2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U821 ( .A1(G8), .A2(n731), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U823 ( .A(n734), .B(KEYINPUT98), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n738) );
  AND2_X1 U825 ( .A1(G286), .A2(G8), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n738), .A2(n737), .ZN(n746) );
  INV_X1 U827 ( .A(G8), .ZN(n744) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n784), .ZN(n741) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U830 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U831 ( .A1(n742), .A2(G303), .ZN(n743) );
  OR2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  AND2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U834 ( .A(n747), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U835 ( .A1(n749), .A2(n748), .ZN(n780) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n772) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U838 ( .A1(n772), .A2(n750), .ZN(n919) );
  NAND2_X1 U839 ( .A1(n780), .A2(n919), .ZN(n751) );
  XNOR2_X1 U840 ( .A(n751), .B(KEYINPUT99), .ZN(n754) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n918) );
  INV_X1 U842 ( .A(n784), .ZN(n752) );
  NAND2_X1 U843 ( .A1(n918), .A2(n752), .ZN(n753) );
  NOR2_X1 U844 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U845 ( .A(n755), .B(KEYINPUT64), .ZN(n756) );
  NOR2_X1 U846 ( .A1(KEYINPUT33), .A2(n756), .ZN(n777) );
  XOR2_X1 U847 ( .A(G1981), .B(G305), .Z(n925) );
  XNOR2_X1 U848 ( .A(G1986), .B(G290), .ZN(n914) );
  NAND2_X1 U849 ( .A1(G160), .A2(G40), .ZN(n757) );
  NOR2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n823) );
  NAND2_X1 U851 ( .A1(n914), .A2(n823), .ZN(n759) );
  XNOR2_X1 U852 ( .A(n759), .B(KEYINPUT90), .ZN(n771) );
  NAND2_X1 U853 ( .A1(G104), .A2(n874), .ZN(n761) );
  NAND2_X1 U854 ( .A1(G140), .A2(n872), .ZN(n760) );
  NAND2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n763) );
  XOR2_X1 U856 ( .A(KEYINPUT34), .B(KEYINPUT91), .Z(n762) );
  XNOR2_X1 U857 ( .A(n763), .B(n762), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n878), .A2(G128), .ZN(n765) );
  NAND2_X1 U859 ( .A1(G116), .A2(n879), .ZN(n764) );
  NAND2_X1 U860 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U861 ( .A(KEYINPUT35), .B(n766), .Z(n767) );
  NOR2_X1 U862 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U863 ( .A(n769), .B(KEYINPUT36), .ZN(n770) );
  XNOR2_X1 U864 ( .A(n770), .B(KEYINPUT92), .ZN(n895) );
  XNOR2_X1 U865 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NOR2_X1 U866 ( .A1(n895), .A2(n820), .ZN(n989) );
  NAND2_X1 U867 ( .A1(n823), .A2(n989), .ZN(n817) );
  AND2_X1 U868 ( .A1(n771), .A2(n817), .ZN(n788) );
  AND2_X1 U869 ( .A1(n925), .A2(n788), .ZN(n775) );
  NAND2_X1 U870 ( .A1(KEYINPUT33), .A2(n772), .ZN(n773) );
  NOR2_X1 U871 ( .A1(n784), .A2(n773), .ZN(n774) );
  NOR2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n790) );
  NOR2_X1 U873 ( .A1(G2090), .A2(G303), .ZN(n778) );
  NAND2_X1 U874 ( .A1(G8), .A2(n778), .ZN(n779) );
  NAND2_X1 U875 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U876 ( .A1(n781), .A2(n784), .ZN(n786) );
  NOR2_X1 U877 ( .A1(G1981), .A2(G305), .ZN(n782) );
  XOR2_X1 U878 ( .A(n782), .B(KEYINPUT24), .Z(n783) );
  OR2_X1 U879 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U880 ( .A1(n786), .A2(n785), .ZN(n787) );
  AND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n789) );
  OR2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n810) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(KEYINPUT94), .Z(n792) );
  NAND2_X1 U884 ( .A1(G105), .A2(n874), .ZN(n791) );
  XNOR2_X1 U885 ( .A(n792), .B(n791), .ZN(n796) );
  NAND2_X1 U886 ( .A1(G141), .A2(n872), .ZN(n794) );
  NAND2_X1 U887 ( .A1(G117), .A2(n879), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n878), .A2(G129), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n885) );
  NAND2_X1 U892 ( .A1(G1996), .A2(n885), .ZN(n806) );
  XOR2_X1 U893 ( .A(KEYINPUT93), .B(G1991), .Z(n947) );
  NAND2_X1 U894 ( .A1(G95), .A2(n874), .ZN(n800) );
  NAND2_X1 U895 ( .A1(G131), .A2(n872), .ZN(n799) );
  NAND2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n878), .A2(G119), .ZN(n802) );
  NAND2_X1 U898 ( .A1(G107), .A2(n879), .ZN(n801) );
  NAND2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n803) );
  OR2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n869) );
  NAND2_X1 U901 ( .A1(n947), .A2(n869), .ZN(n805) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n1000) );
  XOR2_X1 U903 ( .A(n823), .B(KEYINPUT95), .Z(n807) );
  NAND2_X1 U904 ( .A1(n1000), .A2(n807), .ZN(n808) );
  XOR2_X1 U905 ( .A(KEYINPUT96), .B(n808), .Z(n813) );
  INV_X1 U906 ( .A(n813), .ZN(n809) );
  NAND2_X1 U907 ( .A1(n810), .A2(n809), .ZN(n825) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n885), .ZN(n995) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U910 ( .A1(n947), .A2(n869), .ZN(n990) );
  NOR2_X1 U911 ( .A1(n811), .A2(n990), .ZN(n812) );
  NOR2_X1 U912 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U913 ( .A1(n995), .A2(n814), .ZN(n815) );
  XOR2_X1 U914 ( .A(KEYINPUT39), .B(n815), .Z(n816) );
  XNOR2_X1 U915 ( .A(KEYINPUT101), .B(n816), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U917 ( .A(n819), .B(KEYINPUT102), .ZN(n821) );
  NAND2_X1 U918 ( .A1(n895), .A2(n820), .ZN(n1002) );
  NAND2_X1 U919 ( .A1(n821), .A2(n1002), .ZN(n822) );
  NAND2_X1 U920 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U922 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n827), .ZN(G217) );
  NAND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n829) );
  INV_X1 U925 ( .A(G661), .ZN(n828) );
  NOR2_X1 U926 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n830), .B(KEYINPUT103), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XOR2_X1 U934 ( .A(KEYINPUT43), .B(G2678), .Z(n836) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(KEYINPUT104), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U937 ( .A(KEYINPUT105), .B(G2090), .Z(n838) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U940 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2096), .B(G2100), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n844) );
  XOR2_X1 U943 ( .A(G2078), .B(G2084), .Z(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1981), .B(G1971), .Z(n846) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1961), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U948 ( .A(n847), .B(G2474), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1956), .B(G1976), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1966), .Z(n851) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U955 ( .A1(G124), .A2(n878), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n874), .A2(G100), .ZN(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G136), .A2(n872), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G112), .A2(n879), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U962 ( .A1(n860), .A2(n859), .ZN(G162) );
  NAND2_X1 U963 ( .A1(n878), .A2(G130), .ZN(n862) );
  NAND2_X1 U964 ( .A1(G118), .A2(n879), .ZN(n861) );
  NAND2_X1 U965 ( .A1(n862), .A2(n861), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G106), .A2(n874), .ZN(n864) );
  NAND2_X1 U967 ( .A1(G142), .A2(n872), .ZN(n863) );
  NAND2_X1 U968 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U969 ( .A(KEYINPUT45), .B(n865), .Z(n866) );
  NOR2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n871) );
  XOR2_X1 U971 ( .A(G162), .B(n988), .Z(n868) );
  XNOR2_X1 U972 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n887) );
  NAND2_X1 U974 ( .A1(G139), .A2(n872), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n873), .B(KEYINPUT108), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G103), .A2(n874), .ZN(n875) );
  XOR2_X1 U977 ( .A(KEYINPUT107), .B(n875), .Z(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n884) );
  NAND2_X1 U979 ( .A1(n878), .A2(G127), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G115), .A2(n879), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n1005) );
  XNOR2_X1 U984 ( .A(n885), .B(n1005), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n894) );
  XOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n889) );
  XNOR2_X1 U987 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U989 ( .A(n890), .B(KEYINPUT109), .Z(n892) );
  XNOR2_X1 U990 ( .A(G160), .B(KEYINPUT106), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U992 ( .A(n894), .B(n893), .Z(n897) );
  XNOR2_X1 U993 ( .A(G164), .B(n895), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U995 ( .A1(G37), .A2(n898), .ZN(G395) );
  XNOR2_X1 U996 ( .A(G286), .B(KEYINPUT112), .ZN(n901) );
  XNOR2_X1 U997 ( .A(G171), .B(n899), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n904), .ZN(G397) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n906), .ZN(n907) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n907), .ZN(n910) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(KEYINPUT113), .B(n908), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(KEYINPUT114), .B(n911), .ZN(G308) );
  INV_X1 U1009 ( .A(G308), .ZN(G225) );
  INV_X1 U1010 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1011 ( .A(KEYINPUT56), .B(G16), .ZN(n939) );
  XOR2_X1 U1012 ( .A(n912), .B(G1341), .Z(n924) );
  AND2_X1 U1013 ( .A1(G303), .A2(G1971), .ZN(n913) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(G1956), .B(KEYINPUT123), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n915), .B(G299), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(KEYINPUT124), .B(n922), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n929) );
  XNOR2_X1 U1022 ( .A(G1966), .B(G168), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1024 ( .A(KEYINPUT57), .B(n927), .Z(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n937) );
  XNOR2_X1 U1026 ( .A(G171), .B(G1961), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(n930), .B(KEYINPUT121), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(G1348), .B(KEYINPUT120), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n932), .B(n931), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(n935), .B(KEYINPUT122), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n1020) );
  XNOR2_X1 U1034 ( .A(G32), .B(n940), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n941), .A2(G28), .ZN(n946) );
  XNOR2_X1 U1036 ( .A(G2067), .B(G26), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(G2072), .B(G33), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(n944), .B(KEYINPUT119), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n952) );
  XNOR2_X1 U1041 ( .A(n947), .B(G25), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G27), .B(n948), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(n953), .B(KEYINPUT53), .ZN(n956) );
  XOR2_X1 U1046 ( .A(G2084), .B(G34), .Z(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT54), .B(n954), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(G35), .B(G2090), .ZN(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(KEYINPUT55), .B(n959), .ZN(n961) );
  INV_X1 U1052 ( .A(G29), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1054 ( .A1(n962), .A2(G11), .ZN(n1018) );
  XOR2_X1 U1055 ( .A(G1961), .B(G5), .Z(n970) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G22), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(G23), .B(G1976), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1059 ( .A(KEYINPUT126), .B(n965), .Z(n967) );
  XNOR2_X1 U1060 ( .A(G1986), .B(G24), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(KEYINPUT58), .B(n968), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n983) );
  XOR2_X1 U1064 ( .A(G1966), .B(G21), .Z(n981) );
  XOR2_X1 U1065 ( .A(G1348), .B(KEYINPUT59), .Z(n971) );
  XNOR2_X1 U1066 ( .A(G4), .B(n971), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(G6), .B(G1981), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(G1341), .B(G19), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(G1956), .B(G20), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n978), .B(KEYINPUT60), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(n979), .B(KEYINPUT125), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1077 ( .A(KEYINPUT61), .B(n984), .Z(n985) );
  NOR2_X1 U1078 ( .A1(G16), .A2(n985), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(KEYINPUT127), .B(n986), .ZN(n1016) );
  XOR2_X1 U1080 ( .A(G2084), .B(G160), .Z(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(KEYINPUT115), .B(n993), .ZN(n998) );
  XOR2_X1 U1085 ( .A(G2090), .B(G162), .Z(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1087 ( .A(KEYINPUT51), .B(n996), .Z(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(n1001), .B(KEYINPUT116), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1092 ( .A(KEYINPUT117), .B(n1004), .Z(n1010) );
  XOR2_X1 U1093 ( .A(G2072), .B(n1005), .Z(n1007) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1008), .Z(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(KEYINPUT52), .B(n1011), .Z(n1012) );
  NOR2_X1 U1099 ( .A1(KEYINPUT55), .A2(n1012), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(KEYINPUT118), .B(n1013), .Z(n1014) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(G29), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1021), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

