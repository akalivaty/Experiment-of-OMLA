//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1154;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT66), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT66), .B(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(new_n473), .A3(G137), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n466), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n471), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n463), .A2(new_n473), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n463), .A2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(G124), .A2(new_n479), .B1(new_n480), .B2(G136), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n473), .C2(G112), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT67), .Z(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND3_X1  g060(.A1(new_n472), .A2(G126), .A3(G2105), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT68), .ZN(new_n491));
  OAI21_X1  g066(.A(G138), .B1(new_n461), .B2(new_n462), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(new_n470), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n490), .A2(KEYINPUT68), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(KEYINPUT4), .C1(new_n492), .C2(new_n470), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n489), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  AOI211_X1 g076(.A(new_n501), .B(new_n489), .C1(new_n496), .C2(new_n498), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n500), .A2(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n510), .A2(new_n513), .ZN(G166));
  NAND3_X1  g089(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n515));
  XOR2_X1   g090(.A(new_n515), .B(KEYINPUT70), .Z(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  INV_X1    g094(.A(G89), .ZN(new_n520));
  OAI221_X1 g095(.A(new_n518), .B1(new_n508), .B2(new_n519), .C1(new_n520), .C2(new_n506), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n516), .A2(new_n521), .ZN(G168));
  INV_X1    g097(.A(G52), .ZN(new_n523));
  INV_X1    g098(.A(G90), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n523), .A2(new_n508), .B1(new_n506), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n512), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(G171));
  AOI22_X1  g103(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT71), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n530), .A2(G651), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  INV_X1    g110(.A(new_n506), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT73), .B(G81), .Z(new_n537));
  INV_X1    g112(.A(new_n508), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(G43), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n534), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  NAND2_X1  g120(.A1(new_n538), .A2(G53), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT9), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(KEYINPUT74), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n546), .B(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n512), .ZN(new_n552));
  INV_X1    g127(.A(G91), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n506), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  INV_X1    g132(.A(G168), .ZN(G286));
  INV_X1    g133(.A(G166), .ZN(G303));
  OAI21_X1  g134(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n560));
  INV_X1    g135(.A(G49), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n508), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(G87), .B2(new_n536), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(G288));
  NAND3_X1  g139(.A1(new_n504), .A2(G48), .A3(G543), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n505), .A2(G61), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n567), .A2(new_n568), .B1(G73), .B2(G543), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n505), .A2(KEYINPUT75), .A3(G61), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n566), .B1(new_n571), .B2(G651), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n505), .A2(new_n504), .A3(G86), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(G85), .A2(new_n536), .B1(new_n538), .B2(G47), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n512), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n578), .B(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n505), .A2(new_n504), .A3(G92), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT10), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n505), .A2(G66), .ZN(new_n584));
  NAND2_X1  g159(.A1(G79), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n512), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(G54), .B2(new_n538), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n581), .B1(new_n589), .B2(G868), .ZN(G284));
  OAI21_X1  g165(.A(new_n581), .B1(new_n589), .B2(G868), .ZN(G321));
  NAND2_X1  g166(.A1(G286), .A2(G868), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(new_n555), .B2(G868), .ZN(G297));
  OAI21_X1  g168(.A(new_n592), .B1(new_n555), .B2(G868), .ZN(G280));
  INV_X1    g169(.A(G860), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n588), .B1(G559), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT77), .ZN(G148));
  NOR2_X1   g172(.A1(new_n588), .A2(G559), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n540), .B2(G868), .ZN(G323));
  XOR2_X1   g176(.A(KEYINPUT78), .B(KEYINPUT11), .Z(new_n602));
  XNOR2_X1  g177(.A(G323), .B(new_n602), .ZN(G282));
  NAND2_X1  g178(.A1(new_n472), .A2(new_n475), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT13), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G2100), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT80), .Z(new_n609));
  AOI22_X1  g184(.A1(G123), .A2(new_n479), .B1(new_n480), .B2(G135), .ZN(new_n610));
  OAI221_X1 g185(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n473), .C2(G111), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(G2096), .Z(new_n613));
  OAI211_X1 g188(.A(new_n609), .B(new_n613), .C1(G2100), .C2(new_n607), .ZN(G156));
  XNOR2_X1  g189(.A(G2427), .B(G2430), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT82), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT81), .B(G2438), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT14), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2451), .B(G2454), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT16), .ZN(new_n624));
  XOR2_X1   g199(.A(G1341), .B(G1348), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n622), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2443), .B(G2446), .Z(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(G14), .A3(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(G401));
  INV_X1    g207(.A(KEYINPUT18), .ZN(new_n633));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT17), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n634), .A2(new_n635), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2100), .ZN(new_n640));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n636), .B2(KEYINPUT18), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2096), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(G227));
  XOR2_X1   g219(.A(G1971), .B(G1976), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT19), .ZN(new_n646));
  XOR2_X1   g221(.A(G1956), .B(G2474), .Z(new_n647));
  XOR2_X1   g222(.A(G1961), .B(G1966), .Z(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n646), .A2(new_n651), .A3(new_n649), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n651), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n654));
  AOI211_X1 g229(.A(new_n650), .B(new_n652), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n653), .B2(new_n654), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1991), .B(G1996), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1981), .B(G1986), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G229));
  INV_X1    g238(.A(G29), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(G25), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n479), .A2(G119), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT84), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n473), .A2(G107), .ZN(new_n668));
  OAI21_X1  g243(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  AOI22_X1  g245(.A1(new_n668), .A2(new_n670), .B1(new_n480), .B2(G131), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n665), .B1(new_n672), .B2(new_n664), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT35), .B(G1991), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n676), .A2(G24), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(G290), .B2(G16), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  OAI211_X1 g255(.A(KEYINPUT87), .B(new_n675), .C1(new_n680), .C2(G1986), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(G1986), .B2(new_n680), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n676), .A2(G6), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G305), .B2(G16), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT32), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n676), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n676), .ZN(new_n691));
  INV_X1    g266(.A(G1971), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n676), .A2(G23), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n563), .B2(new_n676), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT33), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n688), .A2(new_n689), .A3(new_n693), .A4(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT34), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(KEYINPUT34), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n682), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT36), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n664), .A2(G35), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G162), .B2(new_n664), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT29), .B(G2090), .Z(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  AOI22_X1  g282(.A1(new_n480), .A2(G141), .B1(G105), .B2(new_n475), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n479), .A2(G129), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT26), .Z(new_n711));
  NAND3_X1  g286(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT92), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G29), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G29), .B2(G32), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT27), .B(G1996), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT93), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(KEYINPUT94), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(KEYINPUT94), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n707), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n664), .A2(G26), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n480), .A2(G140), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT88), .ZN(new_n726));
  OAI221_X1 g301(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n473), .C2(G116), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n479), .A2(G128), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n724), .B1(new_n729), .B2(G29), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT90), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2067), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  NAND2_X1  g308(.A1(G164), .A2(G29), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G27), .B2(G29), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n732), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT91), .B(KEYINPUT25), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n480), .A2(G139), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n739), .B(new_n740), .C1(new_n473), .C2(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G33), .B(new_n742), .S(G29), .Z(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(G2072), .Z(new_n744));
  NOR2_X1   g319(.A1(G4), .A2(G16), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n589), .B2(G16), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n744), .B1(new_n746), .B2(G1348), .ZN(new_n747));
  NOR2_X1   g322(.A1(G5), .A2(G16), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G171), .B2(G16), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT24), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(G34), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(G34), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n477), .B2(G29), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n751), .B1(new_n752), .B2(new_n758), .C1(new_n717), .C2(new_n715), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n676), .A2(G20), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT23), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n555), .B2(new_n676), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1956), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n676), .A2(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G168), .B2(new_n676), .ZN(new_n765));
  INV_X1    g340(.A(G1966), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n746), .A2(G1348), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n664), .B1(new_n770), .B2(G28), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n771), .A2(KEYINPUT95), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(G28), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n771), .B2(KEYINPUT95), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n769), .B1(new_n772), .B2(new_n774), .C1(new_n612), .C2(new_n664), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n752), .B2(new_n758), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n767), .A2(new_n768), .A3(new_n776), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n747), .A2(new_n759), .A3(new_n763), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n540), .A2(G16), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G16), .B2(G19), .ZN(new_n780));
  INV_X1    g355(.A(G1341), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n735), .A2(new_n733), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n721), .A2(new_n736), .A3(new_n778), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n701), .B2(new_n702), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n703), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(G311));
  INV_X1    g364(.A(KEYINPUT96), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n788), .B(new_n790), .ZN(G150));
  INV_X1    g366(.A(G93), .ZN(new_n792));
  INV_X1    g367(.A(G55), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n506), .A2(new_n792), .B1(new_n508), .B2(new_n793), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(new_n512), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(new_n595), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT37), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n589), .A2(G559), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT38), .Z(new_n801));
  NAND3_X1  g376(.A1(new_n534), .A2(new_n535), .A3(new_n539), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(new_n797), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n801), .B(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(KEYINPUT39), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT97), .Z(new_n807));
  OAI21_X1  g382(.A(new_n595), .B1(new_n805), .B2(KEYINPUT39), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n799), .B1(new_n807), .B2(new_n808), .ZN(G145));
  AOI22_X1  g384(.A1(G130), .A2(new_n479), .B1(new_n480), .B2(G142), .ZN(new_n810));
  OAI221_X1 g385(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n473), .C2(G118), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(new_n606), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(new_n672), .ZN(new_n814));
  INV_X1    g389(.A(new_n489), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n472), .A2(new_n473), .A3(G138), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n494), .B1(new_n816), .B2(new_n491), .ZN(new_n817));
  INV_X1    g392(.A(new_n498), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n729), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n713), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n742), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n742), .A2(new_n712), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n820), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n820), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n827), .B(new_n824), .C1(new_n822), .C2(new_n742), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n814), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n826), .A2(new_n814), .A3(new_n828), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n612), .B(new_n477), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n484), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(G37), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(KEYINPUT99), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n829), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n834), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n836), .A2(new_n838), .A3(new_n831), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n835), .A2(new_n840), .A3(KEYINPUT100), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT40), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT40), .B1(new_n843), .B2(new_n844), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(G395));
  INV_X1    g422(.A(new_n797), .ZN(new_n848));
  INV_X1    g423(.A(G868), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n803), .B(KEYINPUT101), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n598), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n803), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n599), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n555), .A2(new_n588), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n589), .B1(new_n550), .B2(new_n554), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT106), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n857), .B2(new_n858), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n857), .A2(new_n864), .A3(new_n858), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n555), .A2(KEYINPUT102), .A3(new_n588), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n863), .B1(new_n867), .B2(new_n862), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n852), .A2(new_n855), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n860), .A2(new_n861), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n861), .B1(new_n860), .B2(new_n869), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n563), .B(KEYINPUT103), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G290), .ZN(new_n873));
  XNOR2_X1  g448(.A(G305), .B(G303), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n878), .A3(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n870), .B1(new_n871), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n882), .B(KEYINPUT42), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n886), .A2(new_n861), .A3(new_n860), .A4(new_n869), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n850), .B1(new_n888), .B2(new_n849), .ZN(G295));
  OAI21_X1  g464(.A(new_n850), .B1(new_n888), .B2(new_n849), .ZN(G331));
  NAND2_X1  g465(.A1(new_n803), .A2(G301), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n540), .A2(new_n797), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n802), .A2(new_n848), .ZN(new_n893));
  OAI21_X1  g468(.A(G171), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n891), .A2(G168), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n803), .A2(G301), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n892), .A2(G171), .A3(new_n893), .ZN(new_n897));
  OAI21_X1  g472(.A(G286), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n867), .A2(KEYINPUT108), .A3(KEYINPUT41), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n859), .A2(KEYINPUT107), .A3(new_n862), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT41), .B1(new_n857), .B2(new_n858), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n901), .A2(KEYINPUT107), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT108), .B1(new_n867), .B2(KEYINPUT41), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n895), .B(new_n898), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n891), .A2(G168), .A3(new_n894), .ZN(new_n906));
  AOI21_X1  g481(.A(G168), .B1(new_n891), .B2(new_n894), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n859), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n880), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  INV_X1    g487(.A(new_n880), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n898), .A2(new_n868), .A3(new_n895), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n912), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n913), .B1(new_n908), .B2(new_n914), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n913), .B1(new_n905), .B2(new_n908), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n917), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(KEYINPUT109), .B(KEYINPUT43), .C1(new_n917), .C2(new_n922), .ZN(new_n926));
  OR3_X1    g501(.A1(new_n917), .A2(KEYINPUT43), .A3(new_n918), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n921), .B1(new_n928), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g504(.A(G1384), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n819), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n932));
  INV_X1    g507(.A(G40), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n477), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n935), .A2(KEYINPUT110), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(KEYINPUT110), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G1996), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(KEYINPUT46), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT126), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT46), .B1(new_n938), .B2(new_n939), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n936), .A2(new_n937), .ZN(new_n943));
  INV_X1    g518(.A(new_n712), .ZN(new_n944));
  INV_X1    g519(.A(G2067), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n729), .B(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT47), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n713), .A2(new_n939), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n946), .B(new_n951), .C1(new_n939), .C2(new_n944), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n672), .B(new_n674), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(new_n943), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n943), .A2(G1986), .A3(G290), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(KEYINPUT48), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(KEYINPUT48), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n672), .A2(new_n674), .ZN(new_n960));
  OAI22_X1  g535(.A1(new_n952), .A2(new_n960), .B1(G2067), .B2(new_n729), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n958), .A2(new_n959), .B1(new_n938), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n950), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT127), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT127), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n950), .A2(new_n965), .A3(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n819), .A2(KEYINPUT112), .A3(new_n930), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n499), .B2(G1384), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n972), .A2(new_n934), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n819), .A2(new_n501), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n499), .A2(KEYINPUT69), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT113), .B1(new_n976), .B2(new_n971), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n930), .B1(new_n500), .B2(new_n502), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT50), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n973), .A2(new_n977), .A3(new_n752), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT112), .B1(new_n819), .B2(new_n930), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n499), .A2(new_n969), .A3(G1384), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n932), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(KEYINPUT45), .B(new_n930), .C1(new_n500), .C2(new_n502), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n934), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n766), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n981), .A2(G168), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(G8), .ZN(new_n989));
  AOI21_X1  g564(.A(G168), .B1(new_n981), .B2(new_n987), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n981), .B2(new_n987), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT51), .B1(new_n993), .B2(KEYINPUT123), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n981), .A2(new_n987), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G8), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT123), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n989), .B1(new_n999), .B2(KEYINPUT51), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT62), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n989), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n994), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT62), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1003), .B(new_n1004), .C1(new_n994), .C2(new_n991), .ZN(new_n1005));
  INV_X1    g580(.A(G2090), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n973), .A2(new_n977), .A3(new_n1006), .A4(new_n980), .ZN(new_n1007));
  INV_X1    g582(.A(new_n934), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n499), .A2(G1384), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(KEYINPUT45), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n976), .B2(KEYINPUT45), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n692), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(G303), .A2(G8), .B1(KEYINPUT114), .B2(KEYINPUT55), .ZN(new_n1014));
  NOR2_X1   g589(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT115), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1014), .B(new_n1016), .Z(new_n1017));
  NAND3_X1  g592(.A1(new_n1013), .A2(G8), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT49), .ZN(new_n1019));
  INV_X1    g594(.A(G1981), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT117), .B(G86), .Z(new_n1021));
  NAND2_X1  g596(.A1(new_n536), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1020), .B1(new_n572), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n512), .B1(new_n569), .B2(new_n570), .ZN(new_n1024));
  NOR4_X1   g599(.A1(new_n1024), .A2(G1981), .A3(new_n573), .A4(new_n566), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1019), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n572), .A2(new_n1020), .A3(new_n574), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n536), .A2(new_n1021), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1024), .A2(new_n566), .A3(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1027), .B(KEYINPUT49), .C1(new_n1020), .C2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n968), .A2(new_n970), .A3(new_n934), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1026), .A2(new_n1030), .A3(G8), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n563), .A2(G1976), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(G8), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1031), .A2(G8), .A3(new_n1033), .A4(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT116), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1039), .A2(KEYINPUT116), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1036), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n976), .A2(KEYINPUT118), .A3(new_n971), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n971), .B(new_n930), .C1(new_n500), .C2(new_n502), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n968), .A2(new_n970), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1008), .B1(new_n1048), .B2(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1006), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n992), .B1(new_n1050), .B2(new_n1012), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1018), .B(new_n1042), .C1(new_n1017), .C2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n973), .A2(new_n980), .A3(new_n977), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n750), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n1011), .B2(G2078), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n733), .A2(KEYINPUT53), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n986), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(G171), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1052), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1001), .A2(new_n1005), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n992), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1042), .A2(new_n1017), .A3(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1032), .A2(new_n1037), .A3(new_n563), .ZN(new_n1065));
  OAI211_X1 g640(.A(G8), .B(new_n1031), .C1(new_n1065), .C2(new_n1025), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT63), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n993), .A2(G168), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(new_n1052), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1068), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1063), .A2(new_n1017), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1071), .A2(new_n1018), .A3(new_n1042), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1067), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1062), .A2(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1059), .A2(G171), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT53), .B1(new_n1078), .B2(G2078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n1078), .B2(G2078), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1010), .B(new_n1080), .C1(KEYINPUT45), .C2(new_n1009), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1054), .A2(new_n1056), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1077), .B1(new_n1082), .B2(G171), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1052), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1054), .A2(G301), .A3(new_n1056), .A4(new_n1081), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1060), .A2(KEYINPUT125), .A3(new_n1085), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1085), .A2(KEYINPUT125), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(new_n1077), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1003), .B1(new_n994), .B2(new_n991), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n554), .B2(KEYINPUT120), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n555), .B(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT119), .B(G1956), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1010), .B(new_n1097), .C1(new_n976), .C2(KEYINPUT45), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1094), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n979), .B1(new_n978), .B2(KEYINPUT50), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n972), .A2(new_n934), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1348), .B1(new_n1103), .B2(new_n980), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1031), .A2(G2067), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1100), .B1(new_n1106), .B2(new_n588), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1096), .A2(new_n1094), .A3(new_n1099), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT61), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT118), .B1(new_n976), .B2(new_n971), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1049), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1095), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1093), .B1(new_n1116), .B2(new_n1098), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1111), .B1(new_n1117), .B2(new_n1108), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n934), .B1(new_n931), .B2(new_n932), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n932), .B2(new_n978), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  AOI22_X1  g696(.A1(new_n1120), .A2(new_n939), .B1(new_n1031), .B2(new_n1121), .ZN(new_n1122));
  OR3_X1    g697(.A1(new_n1122), .A2(KEYINPUT59), .A3(new_n802), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT59), .B1(new_n1122), .B2(new_n802), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1127));
  INV_X1    g702(.A(G1348), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1053), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1105), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(KEYINPUT60), .A3(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n589), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1106), .A2(KEYINPUT60), .A3(new_n588), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1118), .A2(new_n1125), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1116), .A2(new_n1135), .A3(new_n1093), .A4(new_n1098), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(KEYINPUT61), .A3(new_n1100), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1108), .A2(new_n1135), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1110), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1090), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT122), .B(new_n1110), .C1(new_n1134), .C2(new_n1139), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1075), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g719(.A1(G290), .A2(G1986), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n956), .B1(new_n938), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT111), .ZN(new_n1147));
  OR2_X1    g722(.A1(new_n1147), .A2(new_n955), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n967), .B1(new_n1144), .B2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g724(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1151));
  NAND2_X1  g725(.A1(new_n662), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g726(.A(new_n1152), .B1(new_n843), .B2(new_n844), .ZN(new_n1153));
  NAND2_X1  g727(.A1(new_n916), .A2(new_n919), .ZN(new_n1154));
  AND2_X1   g728(.A1(new_n1153), .A2(new_n1154), .ZN(G308));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(G225));
endmodule


