//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(new_n189), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n193), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G104), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G107), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT78), .A3(G101), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n197), .A3(G104), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .A4(new_n200), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n209), .A2(new_n213), .A3(G143), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n211), .B(G146), .C1(new_n209), .C2(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT78), .ZN(new_n219));
  XNOR2_X1  g033(.A(G104), .B(G107), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(new_n206), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n208), .A2(KEYINPUT10), .A3(new_n218), .A4(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n203), .A2(new_n205), .A3(new_n200), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G101), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT4), .A3(new_n207), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT0), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n209), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n212), .A2(new_n214), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n212), .A2(new_n214), .A3(new_n228), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n223), .A2(new_n232), .A3(G101), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n225), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n218), .A2(new_n221), .A3(new_n207), .A4(new_n202), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT10), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n222), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT64), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI22_X1  g054(.A1(new_n239), .A2(KEYINPUT11), .B1(new_n240), .B2(G137), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT11), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT64), .A4(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n239), .A2(KEYINPUT11), .B1(new_n240), .B2(G137), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n246), .B1(new_n245), .B2(new_n247), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT79), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND4_X1   g064(.A1(KEYINPUT64), .A2(new_n242), .A3(new_n243), .A4(G134), .ZN(new_n251));
  AOI22_X1  g065(.A1(KEYINPUT64), .A2(new_n242), .B1(new_n243), .B2(G134), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n247), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G131), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n246), .B(new_n247), .C1(new_n251), .C2(new_n252), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n196), .B1(new_n238), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT81), .ZN(new_n260));
  INV_X1    g074(.A(new_n218), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n202), .A2(new_n207), .ZN(new_n262));
  INV_X1    g076(.A(new_n221), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n235), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n254), .A2(new_n256), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT12), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n265), .A2(KEYINPUT12), .A3(new_n266), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n272), .B(new_n196), .C1(new_n238), .C2(new_n258), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n260), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n196), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n238), .A2(new_n266), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n238), .A2(new_n258), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT80), .B(G469), .Z(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n192), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n269), .A2(new_n270), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n275), .B1(new_n283), .B2(new_n277), .ZN(new_n284));
  OR2_X1    g098(.A1(new_n276), .A2(new_n259), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(G469), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n190), .B1(new_n282), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT92), .ZN(new_n288));
  XOR2_X1   g102(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G140), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G125), .ZN(new_n292));
  INV_X1    g106(.A(G125), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G140), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT19), .ZN(new_n296));
  XNOR2_X1  g110(.A(G125), .B(G140), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT76), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n213), .B(new_n296), .C1(new_n298), .C2(KEYINPUT19), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n292), .A2(new_n294), .A3(KEYINPUT75), .A4(KEYINPUT16), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n292), .A2(new_n294), .A3(KEYINPUT16), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n292), .B2(KEYINPUT16), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n300), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G146), .ZN(new_n305));
  INV_X1    g119(.A(G237), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(new_n194), .A3(G214), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT87), .A2(G143), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n211), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n307), .A2(new_n308), .ZN(new_n312));
  OAI21_X1  g126(.A(G131), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n307), .A2(new_n308), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n310), .A2(new_n308), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n246), .B(new_n314), .C1(new_n315), .C2(new_n307), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n299), .A2(new_n305), .A3(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n295), .A2(KEYINPUT76), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n297), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n213), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n295), .A2(G146), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OR3_X1    g138(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT18), .ZN(new_n325));
  OAI211_X1 g139(.A(KEYINPUT18), .B(G131), .C1(new_n311), .C2(new_n312), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n324), .A2(new_n316), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G113), .B(G122), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT88), .B(G104), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n318), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n213), .B(new_n300), .C1(new_n301), .C2(new_n303), .ZN(new_n333));
  OAI211_X1 g147(.A(KEYINPUT17), .B(G131), .C1(new_n311), .C2(new_n312), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n305), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT89), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n317), .A2(KEYINPUT17), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n305), .A2(new_n338), .A3(new_n333), .A4(new_n334), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n327), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n332), .B1(new_n341), .B2(new_n330), .ZN(new_n342));
  NOR2_X1   g156(.A1(G475), .A2(G902), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n290), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n331), .B1(new_n340), .B2(new_n327), .ZN(new_n345));
  INV_X1    g159(.A(new_n343), .ZN(new_n346));
  NOR4_X1   g160(.A1(new_n345), .A2(KEYINPUT20), .A3(new_n346), .A4(new_n332), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT90), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n344), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n331), .A2(KEYINPUT91), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n341), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n340), .A2(KEYINPUT91), .A3(new_n327), .A4(new_n331), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n189), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G475), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n342), .A2(new_n348), .A3(new_n355), .A4(new_n343), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n288), .B1(new_n349), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n347), .A2(new_n348), .B1(new_n353), .B2(G475), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n341), .A2(new_n330), .ZN(new_n360));
  INV_X1    g174(.A(new_n332), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n360), .A2(new_n355), .A3(new_n343), .A4(new_n361), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n345), .A2(new_n346), .A3(new_n332), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n362), .B(KEYINPUT90), .C1(new_n363), .C2(new_n290), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n359), .A2(new_n364), .A3(KEYINPUT92), .ZN(new_n365));
  XNOR2_X1  g179(.A(G128), .B(G143), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT13), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n211), .A2(G128), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n367), .B(G134), .C1(KEYINPUT13), .C2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G116), .B(G122), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(new_n197), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n366), .A2(new_n240), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n366), .B(new_n240), .ZN(new_n374));
  INV_X1    g188(.A(G116), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(KEYINPUT14), .A3(G122), .ZN(new_n376));
  INV_X1    g190(.A(new_n370), .ZN(new_n377));
  OAI211_X1 g191(.A(G107), .B(new_n376), .C1(new_n377), .C2(KEYINPUT14), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n370), .A2(new_n197), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n188), .A2(G217), .A3(new_n194), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n189), .ZN(new_n384));
  INV_X1    g198(.A(G478), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(KEYINPUT15), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n386), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n194), .A2(G952), .ZN(new_n390));
  NAND2_X1  g204(.A1(G234), .A2(G237), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(KEYINPUT21), .B(G898), .Z(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(G902), .A3(G953), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  AND4_X1   g211(.A1(new_n287), .A2(new_n358), .A3(new_n365), .A4(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT68), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT31), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n229), .A2(new_n230), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n254), .B2(new_n256), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n243), .A2(G134), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n240), .A2(G137), .ZN(new_n404));
  OAI21_X1  g218(.A(G131), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n256), .A2(new_n218), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT2), .ZN(new_n407));
  INV_X1    g221(.A(G113), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT66), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT66), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(KEYINPUT2), .B2(G113), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n409), .A2(new_n411), .B1(KEYINPUT2), .B2(G113), .ZN(new_n412));
  INV_X1    g226(.A(G119), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G116), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n375), .A2(G119), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n412), .B(new_n417), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n402), .A2(new_n406), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT30), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n420), .A2(KEYINPUT65), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(KEYINPUT65), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n421), .B(new_n422), .C1(new_n402), .C2(new_n406), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n231), .B1(new_n248), .B2(new_n249), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n256), .A2(new_n218), .A3(new_n405), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n424), .A2(KEYINPUT65), .A3(new_n420), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n419), .B1(new_n427), .B2(new_n418), .ZN(new_n428));
  NOR2_X1   g242(.A1(G237), .A2(G953), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G210), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(G101), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n400), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n412), .B(new_n416), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n423), .B2(new_n426), .ZN(new_n436));
  INV_X1    g250(.A(new_n433), .ZN(new_n437));
  NOR4_X1   g251(.A1(new_n436), .A2(KEYINPUT31), .A3(new_n419), .A4(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n435), .B1(new_n424), .B2(new_n425), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT28), .B1(new_n419), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n424), .A2(new_n435), .A3(new_n425), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT28), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n433), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n434), .A2(new_n438), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(G472), .A2(G902), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT67), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n399), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n427), .A2(new_n418), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n441), .A3(new_n433), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT31), .ZN(new_n451));
  INV_X1    g265(.A(new_n444), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n428), .A2(new_n400), .A3(new_n433), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n447), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n454), .A2(KEYINPUT32), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT32), .B1(new_n454), .B2(new_n455), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n448), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n418), .B1(new_n402), .B2(new_n406), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n441), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT70), .B1(new_n460), .B2(KEYINPUT28), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT70), .ZN(new_n462));
  AOI211_X1 g276(.A(new_n462), .B(new_n442), .C1(new_n459), .C2(new_n441), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n464), .A2(KEYINPUT29), .A3(new_n443), .A4(new_n433), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n189), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n440), .A2(new_n443), .A3(new_n433), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT69), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT69), .B1(new_n428), .B2(new_n433), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n470), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G472), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n454), .A2(new_n455), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n399), .A3(KEYINPUT32), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n458), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT72), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n209), .A2(G119), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT23), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(KEYINPUT72), .B(KEYINPUT23), .C1(new_n209), .C2(G119), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(KEYINPUT73), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n413), .A2(G128), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n483), .B(new_n479), .C1(new_n477), .C2(KEYINPUT73), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(G110), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT74), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n305), .A2(new_n333), .ZN(new_n489));
  XOR2_X1   g303(.A(KEYINPUT24), .B(G110), .Z(new_n490));
  INV_X1    g304(.A(new_n478), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n484), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT74), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n485), .A2(new_n493), .A3(G110), .A4(new_n486), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n488), .A2(new_n489), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(G110), .B1(new_n485), .B2(new_n486), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n490), .B1(new_n484), .B2(new_n491), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n305), .B(new_n322), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT22), .B(G137), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT77), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n495), .A2(new_n498), .A3(new_n502), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n189), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT25), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G234), .ZN(new_n510));
  OAI21_X1  g324(.A(G217), .B1(new_n510), .B2(G902), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT71), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n505), .A2(new_n506), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n512), .A2(G902), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n509), .A2(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XOR2_X1   g330(.A(G110), .B(G122), .Z(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n418), .A2(new_n233), .A3(new_n225), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n375), .A2(G119), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT5), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n408), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n414), .A2(new_n415), .A3(KEYINPUT5), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n412), .A2(new_n417), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n208), .A2(new_n524), .A3(new_n221), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n518), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n526), .A2(KEYINPUT6), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n225), .A2(new_n233), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n525), .B(new_n518), .C1(new_n528), .C2(new_n435), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT82), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT82), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n519), .A2(new_n531), .A3(new_n525), .A4(new_n518), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n526), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT6), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n527), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n231), .A2(G125), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n218), .A2(new_n293), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n194), .A2(G224), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n539), .B1(new_n536), .B2(new_n537), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n535), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G210), .B1(G237), .B2(G902), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n545), .B(KEYINPUT85), .Z(new_n546));
  NOR2_X1   g360(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n541), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n538), .A2(KEYINPUT7), .A3(new_n540), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n262), .A2(new_n263), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT84), .ZN(new_n552));
  OR3_X1    g366(.A1(new_n551), .A2(new_n552), .A3(new_n524), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n552), .B1(new_n551), .B2(new_n524), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n412), .A2(new_n417), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT83), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n522), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n522), .A2(new_n556), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n523), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n551), .B(new_n555), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n553), .A2(new_n554), .A3(new_n560), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n517), .B(KEYINPUT8), .Z(new_n562));
  AOI22_X1  g376(.A1(new_n561), .A2(new_n562), .B1(new_n530), .B2(new_n532), .ZN(new_n563));
  AOI21_X1  g377(.A(G902), .B1(new_n550), .B2(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n544), .A2(new_n546), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n546), .B1(new_n544), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(G214), .B1(G237), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n398), .A2(new_n476), .A3(new_n516), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G101), .ZN(G3));
  INV_X1    g385(.A(new_n384), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(G478), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT93), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n383), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT33), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n383), .A2(new_n574), .A3(KEYINPUT33), .ZN(new_n578));
  AOI21_X1  g392(.A(G902), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n573), .B1(new_n579), .B2(G478), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n358), .B2(new_n365), .ZN(new_n581));
  OAI21_X1  g395(.A(G472), .B1(new_n445), .B2(G902), .ZN(new_n582));
  INV_X1    g396(.A(new_n190), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n274), .A2(new_n278), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n189), .A3(new_n281), .ZN(new_n585));
  INV_X1    g399(.A(new_n192), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n286), .A3(new_n586), .ZN(new_n587));
  AND4_X1   g401(.A1(new_n474), .A2(new_n582), .A3(new_n583), .A4(new_n587), .ZN(new_n588));
  NOR4_X1   g402(.A1(new_n565), .A2(new_n566), .A3(new_n568), .A4(new_n396), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n581), .A2(new_n588), .A3(new_n516), .A4(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT34), .B(G104), .Z(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  INV_X1    g406(.A(G472), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n454), .B2(new_n189), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n445), .A2(new_n447), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n596), .A2(new_n516), .A3(new_n287), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n363), .A2(new_n290), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n354), .B1(new_n598), .B2(new_n344), .ZN(new_n599));
  INV_X1    g413(.A(new_n389), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n597), .A2(new_n589), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G107), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  INV_X1    g419(.A(new_n566), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n544), .A2(new_n546), .A3(new_n564), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n515), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT36), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n503), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n495), .A2(new_n498), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n613), .B1(new_n495), .B2(new_n498), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n611), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n616), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n614), .A3(new_n610), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n609), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n509), .B2(new_n512), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n608), .A2(new_n621), .A3(new_n568), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n398), .A2(new_n596), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT37), .B(G110), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G12));
  INV_X1    g439(.A(KEYINPUT96), .ZN(new_n626));
  OR3_X1    g440(.A1(new_n394), .A2(new_n626), .A3(G900), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n626), .B1(new_n394), .B2(G900), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n392), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT97), .Z(new_n630));
  NOR2_X1   g444(.A1(new_n601), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n476), .A2(new_n631), .A3(new_n622), .A4(new_n287), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT98), .B(G128), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G30));
  INV_X1    g448(.A(new_n428), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n433), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n189), .B1(new_n460), .B2(new_n433), .ZN(new_n638));
  OAI21_X1  g452(.A(G472), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n458), .A2(new_n475), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n630), .B(KEYINPUT39), .Z(new_n642));
  AND2_X1   g456(.A1(new_n287), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n621), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n641), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n359), .A2(new_n364), .A3(KEYINPUT92), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT92), .B1(new_n359), .B2(new_n364), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n650), .A2(new_n568), .A3(new_n600), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n643), .A2(new_n644), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n608), .B(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n647), .A2(new_n651), .A3(new_n652), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G143), .ZN(G45));
  AOI211_X1 g471(.A(new_n580), .B(new_n630), .C1(new_n358), .C2(new_n365), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n658), .A2(new_n476), .A3(new_n287), .A4(new_n622), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G146), .ZN(G48));
  INV_X1    g474(.A(new_n516), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT32), .ZN(new_n662));
  AOI211_X1 g476(.A(KEYINPUT68), .B(new_n662), .C1(new_n454), .C2(new_n455), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n662), .B1(new_n445), .B2(new_n447), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n454), .A2(KEYINPUT32), .A3(new_n455), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n663), .B1(new_n666), .B2(new_n448), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n661), .B1(new_n667), .B2(new_n473), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n585), .B(new_n583), .C1(new_n191), .C2(new_n279), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n279), .A2(new_n191), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n672), .A2(KEYINPUT100), .A3(new_n583), .A4(new_n585), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n668), .A2(new_n581), .A3(new_n589), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  AND3_X1   g491(.A1(new_n671), .A2(new_n569), .A3(new_n673), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n661), .A2(new_n396), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n476), .A3(new_n602), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  AND3_X1   g495(.A1(new_n358), .A2(new_n365), .A3(new_n397), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n678), .A2(new_n476), .A3(new_n682), .A4(new_n646), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G119), .ZN(G21));
  OAI211_X1 g498(.A(new_n569), .B(new_n389), .C1(new_n648), .C2(new_n649), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n358), .A2(new_n365), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n688), .A2(KEYINPUT103), .A3(new_n569), .A4(new_n389), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n464), .B2(new_n443), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n440), .A2(new_n462), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n460), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n693), .A2(new_n691), .A3(new_n443), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n437), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n451), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT102), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n699), .B(new_n451), .C1(new_n692), .C2(new_n696), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n453), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n594), .B1(new_n701), .B2(new_n455), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n702), .A2(new_n516), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n690), .A2(new_n703), .A3(new_n395), .A4(new_n674), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  NAND4_X1  g519(.A1(new_n658), .A2(new_n702), .A3(new_n678), .A4(new_n646), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  NAND3_X1  g521(.A1(new_n473), .A2(new_n664), .A3(new_n665), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n516), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT105), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(new_n711), .A3(new_n516), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n580), .ZN(new_n714));
  INV_X1    g528(.A(new_n630), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n688), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n568), .B1(new_n606), .B2(new_n607), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT104), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n286), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n284), .A2(KEYINPUT104), .A3(G469), .A4(new_n285), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n282), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n717), .A2(new_n583), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n713), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(KEYINPUT42), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n721), .A2(new_n583), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n567), .B1(new_n565), .B2(new_n566), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n476), .A2(new_n728), .A3(new_n516), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n725), .A2(KEYINPUT106), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  INV_X1    g547(.A(new_n731), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n713), .B2(new_n723), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n733), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  NAND2_X1  g553(.A1(new_n729), .A2(new_n631), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n688), .A2(new_n580), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n742), .B1(new_n743), .B2(KEYINPUT107), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n745), .B(KEYINPUT43), .C1(new_n688), .C2(new_n580), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n596), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(KEYINPUT44), .A3(new_n748), .A4(new_n646), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n284), .A2(new_n285), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n284), .A2(KEYINPUT45), .A3(new_n285), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(G469), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT46), .B1(new_n754), .B2(new_n586), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n586), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n585), .A3(new_n757), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n758), .A2(new_n583), .A3(new_n642), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n744), .A2(new_n746), .A3(new_n748), .A4(new_n646), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n749), .A2(new_n717), .A3(new_n759), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  XNOR2_X1  g578(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n586), .ZN(new_n767));
  INV_X1    g581(.A(new_n585), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n767), .A2(new_n755), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n766), .B1(new_n769), .B2(new_n190), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n758), .A2(new_n583), .A3(new_n765), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n667), .A2(new_n473), .A3(new_n661), .A4(new_n717), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n772), .A2(new_n716), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n291), .ZN(G42));
  AOI211_X1 g589(.A(new_n594), .B(new_n621), .C1(new_n701), .C2(new_n455), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n717), .A2(new_n671), .A3(new_n673), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n779));
  INV_X1    g593(.A(new_n392), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n747), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n744), .A2(new_n746), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT115), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n777), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT116), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n672), .A2(new_n585), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n190), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n727), .B1(new_n772), .B2(new_n792), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n780), .A2(new_n703), .A3(new_n746), .A4(new_n744), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n782), .A2(new_n661), .A3(new_n640), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n688), .A2(new_n714), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n793), .A2(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n655), .A2(new_n567), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(new_n674), .A3(new_n798), .ZN(new_n799));
  XOR2_X1   g613(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(KEYINPUT113), .A2(KEYINPUT50), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n794), .A2(new_n674), .A3(new_n802), .A4(new_n798), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n797), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n789), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n287), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n667), .B2(new_n473), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n621), .A2(new_n599), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n389), .A2(new_n630), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n813), .B(new_n567), .C1(new_n565), .C2(new_n566), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n810), .A2(new_n811), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n476), .A2(new_n287), .A3(new_n812), .A4(new_n815), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT110), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n729), .A2(new_n631), .B1(new_n723), .B2(new_n776), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT111), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT111), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n819), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n597), .A2(new_n650), .A3(new_n389), .A4(new_n589), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n683), .A2(new_n826), .A3(new_n623), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT109), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n570), .A2(new_n828), .A3(new_n590), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n828), .B1(new_n570), .B2(new_n590), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n704), .B(new_n827), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n675), .A2(new_n680), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n825), .A2(new_n833), .A3(new_n738), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n640), .A2(new_n621), .A3(new_n715), .ZN(new_n836));
  INV_X1    g650(.A(new_n726), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n690), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n706), .A2(new_n659), .A3(new_n632), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n706), .A2(new_n632), .A3(new_n659), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n690), .A2(new_n836), .A3(new_n837), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT112), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n839), .B1(new_n838), .B2(new_n840), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n834), .A2(new_n835), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n842), .A2(KEYINPUT52), .A3(new_n843), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n825), .A2(new_n833), .A3(new_n738), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT53), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(KEYINPUT54), .A3(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n819), .A2(new_n820), .A3(new_n823), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n823), .B1(new_n819), .B2(new_n820), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n683), .A2(new_n826), .A3(new_n623), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n476), .A2(new_n516), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n650), .A2(new_n569), .A3(new_n287), .A4(new_n397), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n590), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT109), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n570), .A2(new_n828), .A3(new_n590), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n724), .A2(KEYINPUT42), .B1(new_n729), .B2(new_n730), .ZN(new_n866));
  INV_X1    g680(.A(new_n832), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n865), .A2(new_n704), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n858), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n849), .A2(new_n869), .A3(KEYINPUT53), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n853), .A2(new_n835), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n785), .A2(new_n787), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n713), .ZN(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n794), .A2(new_n678), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n795), .A2(new_n581), .ZN(new_n880));
  NAND2_X1  g694(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n390), .A3(new_n881), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n855), .A2(new_n873), .A3(new_n883), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n808), .A2(new_n884), .B1(G952), .B2(G953), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT49), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n743), .B1(new_n886), .B2(new_n791), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n886), .B2(new_n791), .ZN(new_n888));
  INV_X1    g702(.A(new_n655), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n640), .A2(new_n661), .A3(new_n568), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n888), .A2(new_n583), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n885), .A2(new_n891), .ZN(G75));
  XNOR2_X1  g706(.A(new_n535), .B(KEYINPUT119), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n543), .B(KEYINPUT55), .Z(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n546), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n189), .B(new_n897), .C1(new_n870), .C2(new_n871), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n898), .B2(KEYINPUT56), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n870), .A2(new_n871), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(G902), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n900), .B(new_n895), .C1(new_n902), .C2(new_n897), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n194), .A2(G952), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n899), .A2(new_n903), .A3(new_n905), .ZN(G51));
  XNOR2_X1  g720(.A(new_n192), .B(KEYINPUT57), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n870), .A2(new_n872), .A3(new_n871), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n872), .B1(new_n870), .B2(new_n871), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n584), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n902), .A2(new_n754), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n904), .B1(new_n911), .B2(new_n912), .ZN(G54));
  AOI21_X1  g727(.A(new_n189), .B1(new_n870), .B2(new_n871), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  INV_X1    g729(.A(new_n342), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .A4(new_n342), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n917), .A2(new_n905), .A3(new_n918), .ZN(G60));
  NAND2_X1  g733(.A1(new_n577), .A2(new_n578), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n855), .A2(new_n873), .ZN(new_n921));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT59), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n920), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n920), .A2(new_n923), .ZN(new_n925));
  INV_X1    g739(.A(new_n909), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n873), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n924), .A2(new_n927), .A3(new_n904), .ZN(G63));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n617), .A2(new_n619), .ZN(new_n930));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT60), .Z(new_n932));
  NAND3_X1  g746(.A1(new_n901), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n905), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n514), .B1(new_n901), .B2(new_n932), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n929), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n901), .A2(new_n932), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n513), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n938), .A2(KEYINPUT61), .A3(new_n905), .A4(new_n933), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n936), .A2(new_n939), .ZN(G66));
  AOI21_X1  g754(.A(new_n194), .B1(new_n393), .B2(G224), .ZN(new_n941));
  INV_X1    g755(.A(new_n833), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(new_n194), .ZN(new_n943));
  INV_X1    g757(.A(G898), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n893), .B1(new_n944), .B2(G953), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n943), .B(new_n945), .ZN(G69));
  NAND2_X1  g760(.A1(new_n840), .A2(KEYINPUT123), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n706), .A2(new_n659), .A3(new_n632), .A4(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n656), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n947), .A2(new_n656), .A3(new_n949), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n774), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n581), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n688), .B2(new_n600), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n958), .A2(new_n668), .A3(new_n643), .A4(new_n717), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n763), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(G953), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n427), .B(KEYINPUT120), .Z(new_n963));
  OAI21_X1  g777(.A(new_n296), .B1(new_n298), .B2(KEYINPUT19), .ZN(new_n964));
  XNOR2_X1  g778(.A(KEYINPUT121), .B(KEYINPUT122), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n964), .B(new_n965), .Z(new_n966));
  XNOR2_X1  g780(.A(new_n963), .B(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OR3_X1    g782(.A1(new_n961), .A2(new_n962), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(G900), .A2(G953), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n749), .A2(new_n717), .A3(new_n762), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n690), .A2(new_n713), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n759), .ZN(new_n974));
  INV_X1    g788(.A(new_n740), .ZN(new_n975));
  AOI211_X1 g789(.A(new_n975), .B(new_n774), .C1(new_n737), .C2(new_n732), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n947), .A2(new_n949), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n968), .B(new_n970), .C1(new_n978), .C2(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n962), .B1(new_n961), .B2(new_n968), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n969), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n982), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n969), .A2(new_n979), .A3(new_n980), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(G72));
  NAND4_X1  g800(.A1(new_n974), .A2(new_n976), .A3(new_n833), .A4(new_n977), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT126), .Z(new_n990));
  NAND2_X1  g804(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n635), .A2(new_n433), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n987), .A2(KEYINPUT127), .A3(new_n990), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n850), .A2(new_n854), .ZN(new_n997));
  INV_X1    g811(.A(new_n994), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n997), .A2(new_n636), .A3(new_n989), .A4(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n956), .A2(new_n833), .A3(new_n960), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n990), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n637), .ZN(new_n1002));
  AND4_X1   g816(.A1(new_n905), .A2(new_n996), .A3(new_n999), .A4(new_n1002), .ZN(G57));
endmodule


