//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1' ..
//Module:
 module locked_locked_c2670( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6,
    G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26,
    G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48,
    G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64,
    G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80,
    G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126,
    G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140,
    G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184,
    G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198,
    G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210,
    G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245,
    G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
    G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273,
    G274, G275, G276, G277, G278, G279, G452, G483, G543, G559, G567, G651,
    G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966,
    G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078,
    G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435,
    G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  , KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64);
input KEYINPUT64;
input KEYINPUT65;
input KEYINPUT66;
input KEYINPUT67;
input KEYINPUT68;
input KEYINPUT69;
input KEYINPUT70;
input KEYINPUT71;
input KEYINPUT72;
input KEYINPUT73;
input KEYINPUT74;
input KEYINPUT75;
input KEYINPUT76;
input KEYINPUT77;
input KEYINPUT78;
input KEYINPUT79;
input KEYINPUT80;
input KEYINPUT81;
input KEYINPUT82;
input KEYINPUT83;
input KEYINPUT84;
input KEYINPUT85;
input KEYINPUT86;
input KEYINPUT87;
input KEYINPUT88;
input KEYINPUT89;
input KEYINPUT90;
input KEYINPUT91;
input KEYINPUT92;
input KEYINPUT93;
input KEYINPUT94;
input KEYINPUT95;
input KEYINPUT96;
input KEYINPUT97;
input KEYINPUT98;
input KEYINPUT99;
input KEYINPUT100;
input KEYINPUT101;
input KEYINPUT102;
input KEYINPUT103;
input KEYINPUT104;
input KEYINPUT105;
input KEYINPUT106;
input KEYINPUT107;
input KEYINPUT108;
input KEYINPUT109;
input KEYINPUT110;
input KEYINPUT111;
input KEYINPUT112;
input KEYINPUT113;
input KEYINPUT114;
input KEYINPUT115;
input KEYINPUT116;
input KEYINPUT117;
input KEYINPUT118;
input KEYINPUT119;
input KEYINPUT120;
input KEYINPUT121;
input KEYINPUT122;
input KEYINPUT123;
input KEYINPUT124;
input KEYINPUT125;
input KEYINPUT126;
input KEYINPUT127;
//Header:
   input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3,
    G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24,
    G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44,
    G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62,
    G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78,
    G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94,
    G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138,
    G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182,
    G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196,
    G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208,
    G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243,
    G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255,
    G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271,
    G272, G273, G274, G275, G276, G277, G278, G279, G452, G483, G543, G559,
    G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961,
    G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072,
    G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430,
    G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n382, new_n386, new_n387, new_n388, new_n389, new_n392, new_n393,
    new_n394, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n410, new_n411, new_n412, new_n413, new_n414, new_n415, new_n416,
    new_n417, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451, new_n452, new_n453, new_n454,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n462, new_n463,
    new_n464, new_n465, new_n466, new_n467, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n489, new_n490, new_n491,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n500,
    new_n501, new_n502, new_n503, new_n504, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n518, new_n519, new_n522, new_n524, new_n525, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n975, new_n976,
    new_n977;
wire RLL_wire_A_64;
wire RLL_wire_A_65;
wire RLL_wire_A_66;
wire RLL_wire_A_67;
wire RLL_wire_A_68;
wire RLL_wire_A_69;
wire RLL_wire_A_70;
wire RLL_wire_A_71;
wire RLL_wire_A_72;
wire RLL_wire_A_73;
wire RLL_wire_A_74;
wire RLL_wire_A_75;
wire RLL_wire_A_76;
wire RLL_wire_A_77;
wire RLL_wire_A_78;
wire RLL_wire_A_79;
wire RLL_wire_A_80;
wire RLL_wire_A_81;
wire RLL_wire_A_82;
wire RLL_wire_A_83;
wire RLL_wire_A_84;
wire RLL_wire_A_85;
wire RLL_wire_A_86;
wire RLL_wire_A_87;
wire RLL_wire_A_88;
wire RLL_wire_A_89;
wire RLL_wire_A_90;
wire RLL_wire_A_91;
wire RLL_wire_A_92;
wire RLL_wire_A_93;
wire RLL_wire_A_94;
wire RLL_wire_A_95;
wire RLL_wire_A_96;
wire RLL_wire_A_97;
wire RLL_wire_A_98;
wire RLL_wire_A_99;
wire RLL_wire_A_100;
wire RLL_wire_A_101;
wire RLL_wire_A_102;
wire RLL_wire_A_103;
wire RLL_wire_A_104;
wire RLL_wire_A_105;
wire RLL_wire_A_106;
wire RLL_wire_A_107;
wire RLL_wire_A_108;
wire RLL_wire_A_109;
wire RLL_wire_A_110;
wire RLL_wire_A_111;
wire RLL_wire_A_112;
wire RLL_wire_A_113;
wire RLL_wire_A_114;
wire RLL_wire_A_115;
wire RLL_wire_A_116;
wire RLL_wire_A_117;
wire RLL_wire_A_118;
wire RLL_wire_A_119;
wire RLL_wire_A_120;
wire RLL_wire_A_121;
wire RLL_wire_A_122;
wire RLL_wire_A_123;
wire RLL_wire_A_124;
wire RLL_wire_A_125;
wire RLL_wire_A_126;
wire RLL_wire_A_127;

//Body:
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(RLL_wire_A_64));
  XNOR2_X1 RLL_XNOR_64 (.A(RLL_wire_A_64), .B(KEYINPUT64), .ZN(G337) );
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(RLL_wire_A_65));
  XOR2_X1 RLL_XOR_65 (.A(RLL_wire_A_65), .B(KEYINPUT65), .Z(G219) );
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n382));
  XOR2_X1   g021(.A(new_n382), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n386));
  XOR2_X1   g025(.A(new_n386), .B(KEYINPUT2), .Z(new_n387));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n388));
  INV_X1    g027(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g028(.A1(new_n387), .A2(new_n389), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n387), .A2(G2106), .ZN(new_n392));
  NAND2_X1  g031(.A1(new_n389), .A2(G567), .ZN(new_n393));
  NAND2_X1  g032(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g033(.A(new_n394), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n396));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(RLL_wire_A_66));
  XNOR2_X1 RLL_XNOR_66 (.A(RLL_wire_A_66), .B(KEYINPUT66), .ZN(new_n397) );
  NAND2_X1  g036(.A1(new_n397), .A2(G125), .ZN(new_n398));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n399));
  AOI21_X1  g038(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g039(.A(G2104), .ZN(new_n401));
  NAND2_X1  g040(.A1(new_n401), .A2(KEYINPUT3), .ZN(new_n402));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n403));
  NAND2_X1  g042(.A1(new_n403), .A2(G2104), .ZN(new_n404));
  NAND4_X1  g043(.A1(new_n402), .A2(new_n404), .A3(G137), .A4(new_n396), .ZN(new_n405));
  NOR2_X1   g044(.A1(new_n401), .A2(G2105), .ZN(new_n406));
  NAND2_X1  g045(.A1(new_n406), .A2(G101), .ZN(new_n407));
  NAND2_X1  g046(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g047(.A1(new_n400), .A2(new_n408), .ZN(G160));
  NAND2_X1  g048(.A1(new_n402), .A2(new_n404), .ZN(new_n410));
  NOR2_X1   g049(.A1(new_n410), .A2(G2105), .ZN(new_n411));
  NAND2_X1  g050(.A1(new_n411), .A2(G136), .ZN(new_n412));
  NOR2_X1   g051(.A1(new_n410), .A2(new_n396), .ZN(new_n413));
  NAND2_X1  g052(.A1(new_n413), .A2(G124), .ZN(new_n414));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n415));
  OAI211_X1 g054(.A(new_n415), .B(G2104), .C1(G112), .C2(new_n396), .ZN(new_n416));
  NAND3_X1  g055(.A1(new_n412), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g056(.A(new_n417), .ZN(G162));
  NAND4_X1  g057(.A1(new_n402), .A2(new_n404), .A3(G126), .A4(G2105), .ZN(new_n419));
  INV_X1    g058(.A(G114), .ZN(RLL_wire_A_67));
  XOR2_X1 RLL_XOR_67 (.A(RLL_wire_A_67), .B(KEYINPUT67), .Z(new_n420) );
  NAND2_X1  g059(.A1(new_n420), .A2(G2105), .ZN(RLL_wire_A_68));
  XNOR2_X1 RLL_XNOR_68 (.A(RLL_wire_A_68), .B(KEYINPUT68), .ZN(new_n421) );
  OAI211_X1 g060(.A(new_n421), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n422));
  NAND2_X1  g061(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g062(.A1(new_n402), .A2(new_n404), .A3(G138), .A4(new_n396), .ZN(new_n424));
  NAND2_X1  g063(.A1(new_n424), .A2(KEYINPUT4), .ZN(new_n425));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n426));
  NAND4_X1  g065(.A1(new_n397), .A2(new_n426), .A3(G138), .A4(new_n396), .ZN(RLL_wire_A_69));
  XNOR2_X1 RLL_XNOR_69 (.A(RLL_wire_A_69), .B(KEYINPUT69), .ZN(new_n427) );
  AOI21_X1  g066(.A(new_n423), .B1(new_n425), .B2(new_n427), .ZN(G164));
  INV_X1    g067(.A(G651), .ZN(new_n429));
  NAND2_X1  g068(.A1(new_n429), .A2(KEYINPUT6), .ZN(RLL_wire_A_70));
  XNOR2_X1 RLL_XNOR_70 (.A(RLL_wire_A_70), .B(KEYINPUT70), .ZN(new_n430) );
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n431));
  NAND2_X1  g070(.A1(new_n431), .A2(G651), .ZN(new_n432));
  NAND4_X1  g071(.A1(new_n430), .A2(new_n432), .A3(G50), .A4(G543), .ZN(new_n433));
  INV_X1    g072(.A(G543), .ZN(new_n434));
  NAND2_X1  g073(.A1(new_n434), .A2(KEYINPUT5), .ZN(new_n435));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n436));
  NAND2_X1  g075(.A1(new_n436), .A2(G543), .ZN(new_n437));
  NAND4_X1  g076(.A1(new_n435), .A2(new_n437), .A3(new_n430), .A4(new_n432), .ZN(new_n438));
  INV_X1    g077(.A(G88), .ZN(new_n439));
  OAI21_X1  g078(.A(new_n433), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g079(.A1(new_n435), .A2(new_n437), .A3(G62), .ZN(new_n441));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n442));
  AOI21_X1  g081(.A(new_n429), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g082(.A1(new_n440), .A2(new_n443), .ZN(RLL_wire_A_71));
  XOR2_X1 RLL_XOR_71 (.A(RLL_wire_A_71), .B(KEYINPUT71), .Z(G166) );
  AND2_X1   g083(.A1(new_n435), .A2(new_n437), .ZN(new_n445));
  NAND3_X1  g084(.A1(new_n445), .A2(G63), .A3(G651), .ZN(new_n446));
  AND2_X1   g085(.A1(new_n430), .A2(new_n432), .ZN(new_n447));
  NAND2_X1  g086(.A1(new_n447), .A2(G543), .ZN(new_n448));
  INV_X1    g087(.A(G51), .ZN(new_n449));
  OAI21_X1  g088(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n451));
  XNOR2_X1  g090(.A(new_n451), .B(KEYINPUT7), .ZN(new_n452));
  INV_X1    g091(.A(G89), .ZN(RLL_wire_A_72));
  XNOR2_X1 RLL_XNOR_72 (.A(RLL_wire_A_72), .B(KEYINPUT72), .ZN(new_n453) );
  OAI21_X1  g092(.A(new_n452), .B1(new_n453), .B2(new_n438), .ZN(new_n454));
  NOR2_X1   g093(.A1(new_n450), .A2(new_n454), .ZN(G168));
  AOI22_X1  g094(.A1(new_n445), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n456));
  NOR2_X1   g095(.A1(new_n456), .A2(new_n429), .ZN(new_n457));
  INV_X1    g096(.A(G52), .ZN(new_n458));
  INV_X1    g097(.A(G90), .ZN(new_n459));
  OAI22_X1  g098(.A1(new_n448), .A2(new_n458), .B1(new_n459), .B2(new_n438), .ZN(new_n460));
  NOR2_X1   g099(.A1(new_n457), .A2(new_n460), .ZN(G171));
  AOI22_X1  g100(.A1(new_n445), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n462));
  NOR2_X1   g101(.A1(new_n462), .A2(new_n429), .ZN(new_n463));
  INV_X1    g102(.A(G43), .ZN(new_n464));
  INV_X1    g103(.A(G81), .ZN(new_n465));
  OAI22_X1  g104(.A1(new_n448), .A2(new_n464), .B1(new_n465), .B2(new_n438), .ZN(new_n466));
  NOR2_X1   g105(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g106(.A1(new_n467), .A2(G860), .ZN(G153));
  NAND4_X1  g107(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g108(.A1(G1), .A2(G3), .ZN(RLL_wire_A_73));
  XOR2_X1 RLL_XOR_73 (.A(RLL_wire_A_73), .B(KEYINPUT73), .Z(new_n470) );
  XNOR2_X1  g109(.A(new_n470), .B(KEYINPUT8), .ZN(RLL_wire_A_74));
  XNOR2_X1 RLL_XNOR_74 (.A(RLL_wire_A_74), .B(KEYINPUT74), .ZN(new_n471) );
  NAND4_X1  g110(.A1(G319), .A2(G483), .A3(G661), .A4(new_n471), .ZN(G188));
  NAND3_X1  g111(.A1(new_n447), .A2(G53), .A3(G543), .ZN(new_n473));
  NAND2_X1  g112(.A1(new_n473), .A2(KEYINPUT9), .ZN(new_n474));
  INV_X1    g113(.A(KEYINPUT9), .ZN(new_n475));
  NAND4_X1  g114(.A1(new_n447), .A2(new_n475), .A3(G53), .A4(G543), .ZN(RLL_wire_A_75));
  XNOR2_X1 RLL_XNOR_75 (.A(RLL_wire_A_75), .B(KEYINPUT75), .ZN(new_n476) );
  NAND2_X1  g115(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g116(.A(new_n438), .ZN(new_n478));
  NAND2_X1  g117(.A1(new_n478), .A2(G91), .ZN(RLL_wire_A_76));
  XOR2_X1 RLL_XOR_76 (.A(RLL_wire_A_76), .B(KEYINPUT76), .Z(new_n479) );
  NAND2_X1  g118(.A1(G78), .A2(G543), .ZN(new_n480));
  NAND2_X1  g119(.A1(new_n435), .A2(new_n437), .ZN(new_n481));
  INV_X1    g120(.A(G65), .ZN(new_n482));
  OAI21_X1  g121(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g122(.A1(new_n483), .A2(G651), .ZN(RLL_wire_A_77));
  XNOR2_X1 RLL_XNOR_77 (.A(RLL_wire_A_77), .B(KEYINPUT77), .ZN(new_n484) );
  NAND3_X1  g123(.A1(new_n477), .A2(new_n479), .A3(new_n484), .ZN(G299));
  INV_X1    g124(.A(G171), .ZN(G301));
  INV_X1    g125(.A(G168), .ZN(G286));
  INV_X1    g126(.A(G166), .ZN(G303));
  NAND2_X1  g127(.A1(new_n478), .A2(G87), .ZN(new_n489));
  NAND3_X1  g128(.A1(new_n447), .A2(G49), .A3(G543), .ZN(new_n490));
  OAI21_X1  g129(.A(G651), .B1(new_n445), .B2(G74), .ZN(new_n491));
  NAND3_X1  g130(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(G288));
  NAND3_X1  g131(.A1(new_n435), .A2(new_n437), .A3(G61), .ZN(new_n493));
  NAND2_X1  g132(.A1(G73), .A2(G543), .ZN(new_n494));
  AOI21_X1  g133(.A(new_n429), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g134(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g135(.A1(new_n478), .A2(G86), .ZN(new_n497));
  NAND4_X1  g136(.A1(new_n430), .A2(new_n432), .A3(G48), .A4(G543), .ZN(new_n498));
  NAND3_X1  g137(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(G305));
  AOI22_X1  g138(.A1(new_n445), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n500));
  NOR2_X1   g139(.A1(new_n500), .A2(new_n429), .ZN(new_n501));
  INV_X1    g140(.A(G47), .ZN(new_n502));
  INV_X1    g141(.A(G85), .ZN(new_n503));
  OAI22_X1  g142(.A1(new_n448), .A2(new_n502), .B1(new_n503), .B2(new_n438), .ZN(new_n504));
  OR2_X1    g143(.A1(new_n501), .A2(new_n504), .ZN(G290));
  NAND2_X1  g144(.A1(G301), .A2(G868), .ZN(new_n506));
  NAND2_X1  g145(.A1(new_n478), .A2(G92), .ZN(new_n507));
  XOR2_X1   g146(.A(new_n507), .B(KEYINPUT10), .Z(RLL_wire_A_78));
  XOR2_X1 RLL_XOR_78 (.A(RLL_wire_A_78), .B(KEYINPUT78), .Z(new_n508) );
  INV_X1    g147(.A(new_n448), .ZN(RLL_wire_A_79));
  XNOR2_X1 RLL_XNOR_79 (.A(RLL_wire_A_79), .B(KEYINPUT79), .ZN(new_n509) );
  NAND2_X1  g148(.A1(G79), .A2(G543), .ZN(RLL_wire_A_80));
  XNOR2_X1 RLL_XNOR_80 (.A(RLL_wire_A_80), .B(KEYINPUT80), .ZN(new_n510) );
  INV_X1    g149(.A(G66), .ZN(new_n511));
  OAI21_X1  g150(.A(new_n510), .B1(new_n481), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g151(.A1(new_n509), .A2(G54), .B1(new_n512), .B2(G651), .ZN(new_n513));
  NAND2_X1  g152(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  INV_X1    g153(.A(new_n514), .ZN(RLL_wire_A_81));
  XOR2_X1 RLL_XOR_81 (.A(RLL_wire_A_81), .B(KEYINPUT81), .Z(new_n515) );
  OAI21_X1  g154(.A(new_n506), .B1(new_n515), .B2(G868), .ZN(G284));
  OAI21_X1  g155(.A(new_n506), .B1(new_n515), .B2(G868), .ZN(G321));
  NAND2_X1  g156(.A1(G286), .A2(G868), .ZN(new_n518));
  INV_X1    g157(.A(G299), .ZN(new_n519));
  OAI21_X1  g158(.A(new_n518), .B1(new_n519), .B2(G868), .ZN(G297));
  OAI21_X1  g159(.A(new_n518), .B1(new_n519), .B2(G868), .ZN(G280));
  INV_X1    g160(.A(G559), .ZN(new_n522));
  OAI21_X1  g161(.A(new_n515), .B1(new_n522), .B2(G860), .ZN(RLL_wire_A_82));
  XNOR2_X1 RLL_XNOR_82 (.A(RLL_wire_A_82), .B(KEYINPUT82), .ZN(G148) );
  NAND2_X1  g162(.A1(new_n515), .A2(new_n522), .ZN(new_n524));
  NAND2_X1  g163(.A1(new_n524), .A2(G868), .ZN(new_n525));
  OAI21_X1  g164(.A(new_n525), .B1(G868), .B2(new_n467), .ZN(G323));
  XNOR2_X1  g165(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g166(.A1(new_n397), .A2(new_n406), .ZN(new_n528));
  XNOR2_X1  g167(.A(new_n528), .B(KEYINPUT12), .ZN(new_n529));
  XNOR2_X1  g168(.A(new_n529), .B(KEYINPUT13), .ZN(new_n530));
  INV_X1    g169(.A(G2100), .ZN(new_n531));
  OR2_X1    g170(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g171(.A1(new_n530), .A2(new_n531), .ZN(RLL_wire_A_83));
  XNOR2_X1 RLL_XNOR_83 (.A(RLL_wire_A_83), .B(KEYINPUT83), .ZN(new_n533) );
  NAND2_X1  g172(.A1(new_n411), .A2(G135), .ZN(new_n534));
  NAND2_X1  g173(.A1(new_n413), .A2(G123), .ZN(new_n535));
  NOR2_X1   g174(.A1(new_n396), .A2(G111), .ZN(new_n536));
  OAI21_X1  g175(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n537));
  OAI211_X1 g176(.A(new_n534), .B(new_n535), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  XOR2_X1   g177(.A(new_n538), .B(G2096), .Z(new_n539));
  NAND3_X1  g178(.A1(new_n532), .A2(new_n533), .A3(new_n539), .ZN(G156));
  XNOR2_X1  g179(.A(G2451), .B(G2454), .ZN(new_n541));
  XNOR2_X1  g180(.A(new_n541), .B(KEYINPUT16), .ZN(new_n542));
  XOR2_X1   g181(.A(G2443), .B(G2446), .Z(new_n543));
  XOR2_X1   g182(.A(new_n542), .B(new_n543), .Z(new_n544));
  INV_X1    g183(.A(KEYINPUT14), .ZN(new_n545));
  XNOR2_X1  g184(.A(KEYINPUT15), .B(G2435), .ZN(new_n546));
  XNOR2_X1  g185(.A(new_n546), .B(G2438), .ZN(new_n547));
  XNOR2_X1  g186(.A(G2427), .B(G2430), .ZN(new_n548));
  AOI21_X1  g187(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g188(.A(new_n549), .B1(new_n548), .B2(new_n547), .ZN(new_n550));
  XNOR2_X1  g189(.A(new_n544), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g190(.A(G1341), .B(G1348), .ZN(new_n552));
  OR2_X1    g191(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g192(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  NAND3_X1  g193(.A1(new_n553), .A2(G14), .A3(new_n554), .ZN(new_n555));
  INV_X1    g194(.A(new_n555), .ZN(G401));
  XOR2_X1   g195(.A(G2084), .B(G2090), .Z(new_n557));
  XNOR2_X1  g196(.A(G2067), .B(G2678), .ZN(new_n558));
  XNOR2_X1  g197(.A(G2072), .B(G2078), .ZN(new_n559));
  NAND3_X1  g198(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  XOR2_X1   g199(.A(new_n560), .B(KEYINPUT18), .Z(new_n561));
  INV_X1    g200(.A(new_n558), .ZN(new_n562));
  INV_X1    g201(.A(new_n559), .ZN(new_n563));
  AOI21_X1  g202(.A(new_n557), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XOR2_X1   g203(.A(new_n559), .B(KEYINPUT17), .Z(new_n565));
  OAI21_X1  g204(.A(new_n564), .B1(new_n565), .B2(new_n562), .ZN(new_n566));
  NAND3_X1  g205(.A1(new_n565), .A2(new_n562), .A3(new_n557), .ZN(RLL_wire_A_84));
  XOR2_X1 RLL_XOR_84 (.A(RLL_wire_A_84), .B(KEYINPUT84), .Z(new_n567) );
  NAND3_X1  g206(.A1(new_n561), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  XOR2_X1   g207(.A(G2096), .B(G2100), .Z(new_n569));
  XNOR2_X1  g208(.A(new_n568), .B(new_n569), .ZN(G227));
  XOR2_X1   g209(.A(G1971), .B(G1976), .Z(new_n571));
  XNOR2_X1  g210(.A(new_n571), .B(KEYINPUT19), .ZN(new_n572));
  XNOR2_X1  g211(.A(G1956), .B(G2474), .ZN(new_n573));
  XNOR2_X1  g212(.A(G1961), .B(G1966), .ZN(new_n574));
  NOR2_X1   g213(.A1(new_n573), .A2(new_n574), .ZN(RLL_wire_A_85));
  XNOR2_X1 RLL_XNOR_85 (.A(RLL_wire_A_85), .B(KEYINPUT85), .ZN(new_n575) );
  NAND2_X1  g214(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g215(.A(new_n576), .B(KEYINPUT20), .ZN(new_n577));
  NAND3_X1  g216(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n578));
  XNOR2_X1  g217(.A(new_n573), .B(new_n574), .ZN(new_n579));
  OAI211_X1 g218(.A(new_n577), .B(new_n578), .C1(new_n572), .C2(new_n579), .ZN(RLL_wire_A_86));
  XNOR2_X1 RLL_XNOR_86 (.A(RLL_wire_A_86), .B(KEYINPUT86), .ZN(new_n580) );
  XOR2_X1   g219(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n581));
  XNOR2_X1  g220(.A(G1981), .B(G1986), .ZN(RLL_wire_A_87));
  XNOR2_X1 RLL_XNOR_87 (.A(RLL_wire_A_87), .B(KEYINPUT87), .ZN(new_n582) );
  XNOR2_X1  g221(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g222(.A(new_n580), .B(new_n583), .ZN(new_n584));
  XOR2_X1   g223(.A(G1991), .B(G1996), .Z(new_n585));
  XNOR2_X1  g224(.A(new_n584), .B(new_n585), .ZN(G229));
  INV_X1    g225(.A(G29), .ZN(new_n587));
  NAND2_X1  g226(.A1(new_n587), .A2(G25), .ZN(new_n588));
  NAND2_X1  g227(.A1(new_n411), .A2(G131), .ZN(new_n589));
  NAND2_X1  g228(.A1(new_n413), .A2(G119), .ZN(new_n590));
  OR2_X1    g229(.A1(G95), .A2(G2105), .ZN(new_n591));
  OAI211_X1 g230(.A(new_n591), .B(G2104), .C1(G107), .C2(new_n396), .ZN(new_n592));
  NAND3_X1  g231(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  INV_X1    g232(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g233(.A(new_n588), .B1(new_n594), .B2(new_n587), .ZN(new_n595));
  XOR2_X1   g234(.A(KEYINPUT35), .B(G1991), .Z(new_n596));
  XOR2_X1   g235(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g236(.A(G16), .ZN(new_n598));
  NAND2_X1  g237(.A1(new_n598), .A2(G24), .ZN(new_n599));
  INV_X1    g238(.A(G290), .ZN(new_n600));
  OAI21_X1  g239(.A(new_n599), .B1(new_n600), .B2(new_n598), .ZN(RLL_wire_A_88));
  XOR2_X1 RLL_XOR_88 (.A(RLL_wire_A_88), .B(KEYINPUT88), .Z(new_n601) );
  XNOR2_X1  g240(.A(new_n601), .B(G1986), .ZN(RLL_wire_A_89));
  XOR2_X1 RLL_XOR_89 (.A(RLL_wire_A_89), .B(KEYINPUT89), .Z(new_n602) );
  INV_X1    g241(.A(KEYINPUT34), .ZN(RLL_wire_A_90));
  XOR2_X1 RLL_XOR_90 (.A(RLL_wire_A_90), .B(KEYINPUT90), .Z(new_n603) );
  MUX2_X1   g242(.A(G6), .B(G305), .S(G16), .Z(new_n604));
  XNOR2_X1  g243(.A(KEYINPUT32), .B(G1981), .ZN(new_n605));
  XNOR2_X1  g244(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NOR2_X1   g245(.A1(G16), .A2(G23), .ZN(new_n607));
  AND3_X1   g246(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n608));
  AOI21_X1  g247(.A(new_n607), .B1(new_n608), .B2(G16), .ZN(new_n609));
  XOR2_X1   g248(.A(KEYINPUT33), .B(G1976), .Z(new_n610));
  XNOR2_X1  g249(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g250(.A1(new_n598), .A2(G22), .ZN(new_n612));
  OAI21_X1  g251(.A(new_n612), .B1(G166), .B2(new_n598), .ZN(new_n613));
  XNOR2_X1  g252(.A(new_n613), .B(G1971), .ZN(new_n614));
  NOR3_X1   g253(.A1(new_n606), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  AOI211_X1 g254(.A(new_n597), .B(new_n602), .C1(new_n603), .C2(new_n615), .ZN(new_n616));
  OR2_X1    g255(.A1(new_n615), .A2(new_n603), .ZN(new_n617));
  NAND2_X1  g256(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g257(.A1(new_n618), .A2(KEYINPUT36), .ZN(new_n619));
  INV_X1    g258(.A(KEYINPUT36), .ZN(RLL_wire_A_91));
  XOR2_X1 RLL_XOR_91 (.A(RLL_wire_A_91), .B(KEYINPUT91), .Z(new_n620) );
  NAND3_X1  g259(.A1(new_n616), .A2(new_n620), .A3(new_n617), .ZN(new_n621));
  NAND2_X1  g260(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g261(.A1(G4), .A2(G16), .ZN(new_n623));
  AOI21_X1  g262(.A(new_n623), .B1(new_n515), .B2(G16), .ZN(RLL_wire_A_92));
  XOR2_X1 RLL_XOR_92 (.A(RLL_wire_A_92), .B(KEYINPUT92), .Z(new_n624) );
  INV_X1    g263(.A(G1348), .ZN(new_n625));
  XNOR2_X1  g264(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g265(.A1(new_n598), .A2(G19), .ZN(new_n627));
  OAI21_X1  g266(.A(new_n627), .B1(new_n467), .B2(new_n598), .ZN(new_n628));
  XOR2_X1   g267(.A(new_n628), .B(G1341), .Z(new_n629));
  NAND2_X1  g268(.A1(new_n411), .A2(G140), .ZN(new_n630));
  NAND2_X1  g269(.A1(new_n413), .A2(G128), .ZN(new_n631));
  OR2_X1    g270(.A1(G104), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g271(.A(new_n632), .B(G2104), .C1(G116), .C2(new_n396), .ZN(new_n633));
  NAND3_X1  g272(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(RLL_wire_A_93));
  XNOR2_X1 RLL_XNOR_93 (.A(RLL_wire_A_93), .B(KEYINPUT93), .ZN(new_n634) );
  NAND2_X1  g273(.A1(new_n634), .A2(G29), .ZN(new_n635));
  NAND2_X1  g274(.A1(new_n587), .A2(G26), .ZN(new_n636));
  XNOR2_X1  g275(.A(new_n636), .B(KEYINPUT28), .ZN(new_n637));
  NAND2_X1  g276(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g277(.A(new_n638), .B(G2067), .Z(new_n639));
  NAND3_X1  g278(.A1(new_n626), .A2(new_n629), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g279(.A1(G29), .A2(G33), .ZN(new_n641));
  NAND3_X1  g280(.A1(new_n396), .A2(G103), .A3(G2104), .ZN(new_n642));
  XOR2_X1   g281(.A(new_n642), .B(KEYINPUT25), .Z(new_n643));
  NAND2_X1  g282(.A1(new_n411), .A2(G139), .ZN(new_n644));
  NAND2_X1  g283(.A1(new_n643), .A2(new_n644), .ZN(RLL_wire_A_94));
  XOR2_X1 RLL_XOR_94 (.A(RLL_wire_A_94), .B(KEYINPUT94), .Z(new_n645) );
  AOI22_X1  g284(.A1(new_n397), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n646));
  NOR2_X1   g285(.A1(new_n646), .A2(new_n396), .ZN(new_n647));
  OR2_X1    g286(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g287(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g288(.A(new_n641), .B1(new_n649), .B2(G29), .ZN(new_n650));
  OR2_X1    g289(.A1(new_n650), .A2(G2072), .ZN(new_n651));
  INV_X1    g290(.A(KEYINPUT24), .ZN(new_n652));
  OAI21_X1  g291(.A(new_n587), .B1(new_n652), .B2(G34), .ZN(RLL_wire_A_95));
  XOR2_X1 RLL_XOR_95 (.A(RLL_wire_A_95), .B(KEYINPUT95), .Z(new_n653) );
  AOI21_X1  g292(.A(new_n653), .B1(new_n652), .B2(G34), .ZN(new_n654));
  AOI21_X1  g293(.A(new_n654), .B1(G160), .B2(G29), .ZN(new_n655));
  NAND2_X1  g294(.A1(new_n655), .A2(G2084), .ZN(new_n656));
  NAND2_X1  g295(.A1(new_n650), .A2(G2072), .ZN(new_n657));
  NAND2_X1  g296(.A1(new_n411), .A2(G141), .ZN(new_n658));
  NAND2_X1  g297(.A1(new_n413), .A2(G129), .ZN(new_n659));
  NAND2_X1  g298(.A1(new_n406), .A2(G105), .ZN(new_n660));
  NAND3_X1  g299(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n661));
  XOR2_X1   g300(.A(new_n661), .B(KEYINPUT26), .Z(new_n662));
  NAND4_X1  g301(.A1(new_n658), .A2(new_n659), .A3(new_n660), .A4(new_n662), .ZN(RLL_wire_A_96));
  XNOR2_X1 RLL_XNOR_96 (.A(RLL_wire_A_96), .B(KEYINPUT96), .ZN(new_n663) );
  INV_X1    g302(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g303(.A1(new_n664), .A2(G29), .ZN(new_n665));
  OAI21_X1  g304(.A(new_n665), .B1(G29), .B2(G32), .ZN(new_n666));
  XNOR2_X1  g305(.A(KEYINPUT27), .B(G1996), .ZN(new_n667));
  NAND2_X1  g306(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g307(.A1(new_n651), .A2(new_n656), .A3(new_n657), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g308(.A1(G168), .A2(G16), .ZN(RLL_wire_A_97));
  XNOR2_X1 RLL_XNOR_97 (.A(RLL_wire_A_97), .B(KEYINPUT97), .ZN(new_n670) );
  OAI21_X1  g309(.A(new_n670), .B1(G16), .B2(G21), .ZN(new_n671));
  INV_X1    g310(.A(G1966), .ZN(new_n672));
  OR2_X1    g311(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g312(.A(KEYINPUT31), .B(G11), .Z(new_n674));
  NOR2_X1   g313(.A1(new_n538), .A2(new_n587), .ZN(new_n675));
  INV_X1    g314(.A(G28), .ZN(new_n676));
  OR2_X1    g315(.A1(new_n676), .A2(KEYINPUT30), .ZN(new_n677));
  AOI21_X1  g316(.A(G29), .B1(new_n676), .B2(KEYINPUT30), .ZN(new_n678));
  AOI211_X1 g317(.A(new_n674), .B(new_n675), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  NAND2_X1  g318(.A1(new_n671), .A2(new_n672), .ZN(new_n680));
  NOR2_X1   g319(.A1(G5), .A2(G16), .ZN(new_n681));
  AOI21_X1  g320(.A(new_n681), .B1(G171), .B2(G16), .ZN(new_n682));
  NAND2_X1  g321(.A1(new_n682), .A2(G1961), .ZN(new_n683));
  NAND4_X1  g322(.A1(new_n673), .A2(new_n679), .A3(new_n680), .A4(new_n683), .ZN(new_n684));
  OR2_X1    g323(.A1(new_n655), .A2(G2084), .ZN(new_n685));
  OAI221_X1 g324(.A(new_n685), .B1(G1961), .B2(new_n682), .C1(new_n666), .C2(new_n667), .ZN(new_n686));
  NAND2_X1  g325(.A1(new_n587), .A2(G27), .ZN(new_n687));
  OAI21_X1  g326(.A(new_n687), .B1(G164), .B2(new_n587), .ZN(new_n688));
  XNOR2_X1  g327(.A(new_n688), .B(G2078), .ZN(new_n689));
  OR4_X1    g328(.A1(new_n669), .A2(new_n684), .A3(new_n686), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g329(.A1(new_n587), .A2(G35), .ZN(new_n691));
  OAI21_X1  g330(.A(new_n691), .B1(G162), .B2(new_n587), .ZN(new_n692));
  XNOR2_X1  g331(.A(new_n692), .B(KEYINPUT29), .ZN(new_n693));
  NOR2_X1   g332(.A1(new_n693), .A2(G2090), .ZN(new_n694));
  NAND2_X1  g333(.A1(new_n693), .A2(G2090), .ZN(RLL_wire_A_98));
  XOR2_X1 RLL_XOR_98 (.A(RLL_wire_A_98), .B(KEYINPUT98), .Z(new_n695) );
  NAND2_X1  g334(.A1(new_n598), .A2(G20), .ZN(new_n696));
  XOR2_X1   g335(.A(new_n696), .B(KEYINPUT23), .Z(new_n697));
  AOI21_X1  g336(.A(new_n697), .B1(G299), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g337(.A(new_n698), .B(G1956), .ZN(new_n699));
  NAND2_X1  g338(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NOR4_X1   g339(.A1(new_n640), .A2(new_n690), .A3(new_n694), .A4(new_n700), .ZN(new_n701));
  AND2_X1   g340(.A1(new_n622), .A2(new_n701), .ZN(G311));
  NAND2_X1  g341(.A1(new_n622), .A2(new_n701), .ZN(G150));
  NAND2_X1  g342(.A1(new_n515), .A2(G559), .ZN(new_n704));
  XNOR2_X1  g343(.A(new_n704), .B(KEYINPUT38), .ZN(RLL_wire_A_99));
  XOR2_X1 RLL_XOR_99 (.A(RLL_wire_A_99), .B(KEYINPUT99), .Z(new_n705) );
  AOI22_X1  g344(.A1(new_n445), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n706));
  NOR2_X1   g345(.A1(new_n706), .A2(new_n429), .ZN(new_n707));
  INV_X1    g346(.A(G55), .ZN(RLL_wire_A_100));
  XNOR2_X1 RLL_XNOR_100 (.A(RLL_wire_A_100), .B(KEYINPUT100), .ZN(new_n708) );
  INV_X1    g347(.A(G93), .ZN(new_n709));
  OAI22_X1  g348(.A1(new_n448), .A2(new_n708), .B1(new_n709), .B2(new_n438), .ZN(new_n710));
  OAI21_X1  g349(.A(new_n467), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g350(.A1(new_n707), .A2(new_n710), .ZN(new_n712));
  OAI21_X1  g351(.A(new_n712), .B1(new_n463), .B2(new_n466), .ZN(new_n713));
  NAND2_X1  g352(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g353(.A(new_n705), .B(new_n714), .ZN(new_n715));
  OR2_X1    g354(.A1(new_n715), .A2(KEYINPUT39), .ZN(new_n716));
  INV_X1    g355(.A(G860), .ZN(new_n717));
  NAND2_X1  g356(.A1(new_n715), .A2(KEYINPUT39), .ZN(new_n718));
  NAND3_X1  g357(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g358(.A1(new_n712), .A2(new_n717), .ZN(new_n720));
  XNOR2_X1  g359(.A(new_n720), .B(KEYINPUT37), .ZN(new_n721));
  NAND2_X1  g360(.A1(new_n719), .A2(new_n721), .ZN(G145));
  XNOR2_X1  g361(.A(new_n538), .B(G160), .ZN(new_n723));
  XNOR2_X1  g362(.A(new_n723), .B(G162), .ZN(new_n724));
  NAND2_X1  g363(.A1(new_n425), .A2(new_n427), .ZN(new_n725));
  AND2_X1   g364(.A1(new_n419), .A2(new_n422), .ZN(new_n726));
  NAND2_X1  g365(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g366(.A(new_n634), .B(new_n727), .ZN(new_n728));
  XNOR2_X1  g367(.A(new_n728), .B(new_n664), .ZN(new_n729));
  NAND2_X1  g368(.A1(new_n729), .A2(new_n649), .ZN(new_n730));
  XNOR2_X1  g369(.A(new_n728), .B(new_n663), .ZN(new_n731));
  NAND2_X1  g370(.A1(new_n731), .A2(new_n648), .ZN(new_n732));
  NAND2_X1  g371(.A1(new_n411), .A2(G142), .ZN(new_n733));
  NAND2_X1  g372(.A1(new_n413), .A2(G130), .ZN(new_n734));
  NOR2_X1   g373(.A1(new_n396), .A2(G118), .ZN(new_n735));
  OAI21_X1  g374(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n736));
  OAI211_X1 g375(.A(new_n733), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  XNOR2_X1  g376(.A(new_n737), .B(new_n593), .ZN(new_n738));
  XNOR2_X1  g377(.A(new_n738), .B(new_n529), .ZN(new_n739));
  INV_X1    g378(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g379(.A1(new_n730), .A2(new_n732), .A3(new_n740), .ZN(RLL_wire_A_101));
  XOR2_X1 RLL_XOR_101 (.A(RLL_wire_A_101), .B(KEYINPUT101), .Z(new_n741) );
  INV_X1    g380(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g381(.A(new_n740), .B1(new_n730), .B2(new_n732), .ZN(new_n743));
  OAI21_X1  g382(.A(new_n724), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g383(.A(G37), .ZN(new_n745));
  NAND2_X1  g384(.A1(new_n730), .A2(new_n732), .ZN(new_n746));
  NAND2_X1  g385(.A1(new_n746), .A2(new_n739), .ZN(new_n747));
  INV_X1    g386(.A(new_n724), .ZN(RLL_wire_A_102));
  XNOR2_X1 RLL_XNOR_102 (.A(RLL_wire_A_102), .B(KEYINPUT102), .ZN(new_n748) );
  NAND3_X1  g387(.A1(new_n747), .A2(new_n748), .A3(new_n741), .ZN(new_n749));
  NAND3_X1  g388(.A1(new_n744), .A2(new_n745), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g389(.A(new_n750), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g390(.A(new_n524), .B(new_n714), .ZN(new_n752));
  NAND3_X1  g391(.A1(new_n508), .A2(G299), .A3(new_n513), .ZN(new_n753));
  INV_X1    g392(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g393(.A(G299), .B1(new_n508), .B2(new_n513), .ZN(new_n755));
  NOR2_X1   g394(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g395(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  INV_X1    g396(.A(new_n755), .ZN(new_n758));
  AOI21_X1  g397(.A(KEYINPUT41), .B1(new_n758), .B2(new_n753), .ZN(new_n759));
  INV_X1    g398(.A(KEYINPUT41), .ZN(new_n760));
  NOR3_X1   g399(.A1(new_n754), .A2(new_n760), .A3(new_n755), .ZN(new_n761));
  OAI21_X1  g400(.A(new_n752), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g401(.A(G290), .B(new_n608), .ZN(new_n763));
  XNOR2_X1  g402(.A(G305), .B(G166), .ZN(new_n764));
  OR2_X1    g403(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g404(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  NAND2_X1  g405(.A1(new_n765), .A2(new_n766), .ZN(RLL_wire_A_103));
  XNOR2_X1 RLL_XNOR_103 (.A(RLL_wire_A_103), .B(KEYINPUT103), .ZN(new_n767) );
  NAND2_X1  g406(.A1(new_n767), .A2(KEYINPUT42), .ZN(new_n768));
  INV_X1    g407(.A(KEYINPUT42), .ZN(new_n769));
  NAND3_X1  g408(.A1(new_n765), .A2(new_n769), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g409(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  AND3_X1   g410(.A1(new_n757), .A2(new_n762), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g411(.A(new_n771), .B1(new_n757), .B2(new_n762), .ZN(new_n773));
  OAI21_X1  g412(.A(G868), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g413(.A(new_n774), .B1(G868), .B2(new_n712), .ZN(G295));
  OAI21_X1  g414(.A(new_n774), .B1(G868), .B2(new_n712), .ZN(G331));
  INV_X1    g415(.A(KEYINPUT44), .ZN(new_n777));
  INV_X1    g416(.A(KEYINPUT43), .ZN(RLL_wire_A_104));
  XNOR2_X1 RLL_XNOR_104 (.A(RLL_wire_A_104), .B(KEYINPUT104), .ZN(new_n778) );
  NAND2_X1  g417(.A1(G301), .A2(G168), .ZN(new_n779));
  NAND2_X1  g418(.A1(G286), .A2(G171), .ZN(new_n780));
  NAND2_X1  g419(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g420(.A1(new_n781), .A2(new_n714), .ZN(new_n782));
  AND2_X1   g421(.A1(new_n781), .A2(new_n714), .ZN(new_n783));
  OAI22_X1  g422(.A1(new_n759), .A2(new_n761), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OR2_X1    g423(.A1(new_n781), .A2(new_n714), .ZN(new_n785));
  NAND2_X1  g424(.A1(new_n781), .A2(new_n714), .ZN(new_n786));
  OAI211_X1 g425(.A(new_n785), .B(new_n786), .C1(new_n755), .C2(new_n754), .ZN(RLL_wire_A_105));
  XNOR2_X1 RLL_XNOR_105 (.A(RLL_wire_A_105), .B(KEYINPUT105), .ZN(new_n787) );
  NAND2_X1  g426(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g427(.A(new_n767), .ZN(RLL_wire_A_106));
  XOR2_X1 RLL_XOR_106 (.A(RLL_wire_A_106), .B(KEYINPUT106), .Z(new_n789) );
  AOI21_X1  g428(.A(G37), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g429(.A1(new_n784), .A2(new_n767), .A3(new_n787), .ZN(new_n791));
  AOI21_X1  g430(.A(new_n778), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g431(.A(new_n760), .B1(new_n754), .B2(new_n755), .ZN(new_n793));
  NAND3_X1  g432(.A1(new_n758), .A2(KEYINPUT41), .A3(new_n753), .ZN(new_n794));
  AOI22_X1  g433(.A1(new_n793), .A2(new_n794), .B1(new_n785), .B2(new_n786), .ZN(new_n795));
  NOR3_X1   g434(.A1(new_n783), .A2(new_n756), .A3(new_n782), .ZN(new_n796));
  OAI21_X1  g435(.A(new_n789), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND4_X1   g436(.A1(new_n778), .A2(new_n797), .A3(new_n791), .A4(new_n745), .ZN(new_n798));
  OAI21_X1  g437(.A(new_n777), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g438(.A1(new_n790), .A2(new_n778), .A3(new_n791), .ZN(new_n800));
  NAND3_X1  g439(.A1(new_n797), .A2(new_n791), .A3(new_n745), .ZN(RLL_wire_A_107));
  XOR2_X1 RLL_XOR_107 (.A(RLL_wire_A_107), .B(KEYINPUT107), .Z(new_n801) );
  NAND2_X1  g440(.A1(new_n801), .A2(KEYINPUT43), .ZN(new_n802));
  NAND3_X1  g441(.A1(new_n800), .A2(new_n802), .A3(KEYINPUT44), .ZN(new_n803));
  NAND2_X1  g442(.A1(new_n799), .A2(new_n803), .ZN(G397));
  INV_X1    g443(.A(G1384), .ZN(new_n805));
  NAND2_X1  g444(.A1(new_n727), .A2(new_n805), .ZN(new_n806));
  INV_X1    g445(.A(KEYINPUT45), .ZN(new_n807));
  INV_X1    g446(.A(G40), .ZN(new_n808));
  NOR3_X1   g447(.A1(new_n400), .A2(new_n808), .A3(new_n408), .ZN(new_n809));
  NAND3_X1  g448(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  OR2_X1    g449(.A1(G290), .A2(G1986), .ZN(new_n811));
  NAND2_X1  g450(.A1(G290), .A2(G1986), .ZN(new_n812));
  AOI21_X1  g451(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g452(.A1(new_n810), .A2(G1996), .ZN(new_n814));
  NAND2_X1  g453(.A1(new_n814), .A2(new_n664), .ZN(RLL_wire_A_108));
  XOR2_X1 RLL_XOR_108 (.A(RLL_wire_A_108), .B(KEYINPUT108), .Z(new_n815) );
  INV_X1    g454(.A(new_n810), .ZN(new_n816));
  NAND3_X1  g455(.A1(new_n816), .A2(G1996), .A3(new_n663), .ZN(new_n817));
  XNOR2_X1  g456(.A(new_n634), .B(G2067), .ZN(new_n818));
  NAND2_X1  g457(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g458(.A1(new_n815), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  XOR2_X1   g459(.A(new_n593), .B(new_n596), .Z(new_n821));
  AOI211_X1 g460(.A(new_n813), .B(new_n820), .C1(new_n816), .C2(new_n821), .ZN(new_n822));
  OAI21_X1  g461(.A(new_n807), .B1(G164), .B2(G1384), .ZN(new_n823));
  NAND3_X1  g462(.A1(new_n727), .A2(KEYINPUT45), .A3(new_n805), .ZN(new_n824));
  NAND3_X1  g463(.A1(new_n823), .A2(new_n824), .A3(new_n809), .ZN(new_n825));
  INV_X1    g464(.A(G1971), .ZN(new_n826));
  NAND2_X1  g465(.A1(new_n825), .A2(new_n826), .ZN(RLL_wire_A_109));
  XOR2_X1 RLL_XOR_109 (.A(RLL_wire_A_109), .B(KEYINPUT109), .Z(new_n827) );
  AOI21_X1  g466(.A(G1384), .B1(new_n725), .B2(new_n726), .ZN(new_n828));
  INV_X1    g467(.A(KEYINPUT50), .ZN(new_n829));
  NAND2_X1  g468(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g469(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n831));
  INV_X1    g470(.A(G2090), .ZN(new_n832));
  NAND4_X1  g471(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n809), .ZN(RLL_wire_A_110));
  XNOR2_X1 RLL_XNOR_110 (.A(RLL_wire_A_110), .B(KEYINPUT110), .ZN(new_n833) );
  NAND2_X1  g472(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g473(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n835));
  INV_X1    g474(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g475(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n837));
  NOR2_X1   g476(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g477(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g478(.A1(new_n834), .A2(G8), .A3(new_n839), .ZN(new_n840));
  INV_X1    g479(.A(G8), .ZN(new_n841));
  AOI21_X1  g480(.A(new_n841), .B1(new_n809), .B2(new_n828), .ZN(new_n842));
  NAND2_X1  g481(.A1(new_n608), .A2(G1976), .ZN(new_n843));
  NAND2_X1  g482(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g483(.A1(new_n844), .A2(KEYINPUT52), .ZN(new_n845));
  INV_X1    g484(.A(G1976), .ZN(RLL_wire_A_111));
  XNOR2_X1 RLL_XNOR_111 (.A(RLL_wire_A_111), .B(KEYINPUT111), .ZN(new_n846) );
  AOI21_X1  g485(.A(KEYINPUT52), .B1(G288), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g486(.A1(new_n842), .A2(new_n843), .A3(new_n847), .ZN(RLL_wire_A_112));
  XOR2_X1 RLL_XOR_112 (.A(RLL_wire_A_112), .B(KEYINPUT112), .Z(new_n848) );
  INV_X1    g487(.A(G1981), .ZN(new_n849));
  NAND4_X1  g488(.A1(new_n496), .A2(new_n497), .A3(new_n849), .A4(new_n498), .ZN(new_n850));
  INV_X1    g489(.A(G86), .ZN(new_n851));
  OAI21_X1  g490(.A(new_n498), .B1(new_n438), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g491(.A(G1981), .B1(new_n852), .B2(new_n495), .ZN(new_n853));
  NAND2_X1  g492(.A1(new_n850), .A2(new_n853), .ZN(RLL_wire_A_113));
  XOR2_X1 RLL_XOR_113 (.A(RLL_wire_A_113), .B(KEYINPUT113), .Z(new_n854) );
  INV_X1    g493(.A(KEYINPUT49), .ZN(new_n855));
  NAND2_X1  g494(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g495(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT49), .ZN(RLL_wire_A_114));
  XOR2_X1 RLL_XOR_114 (.A(RLL_wire_A_114), .B(KEYINPUT114), .Z(new_n857) );
  NAND3_X1  g496(.A1(new_n856), .A2(new_n842), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g497(.A1(new_n845), .A2(new_n848), .A3(new_n858), .ZN(new_n859));
  INV_X1    g498(.A(new_n842), .ZN(new_n860));
  INV_X1    g499(.A(new_n850), .ZN(RLL_wire_A_115));
  XOR2_X1 RLL_XOR_115 (.A(RLL_wire_A_115), .B(KEYINPUT115), .Z(new_n861) );
  NOR2_X1   g500(.A1(G288), .A2(G1976), .ZN(new_n862));
  AOI21_X1  g501(.A(new_n861), .B1(new_n858), .B2(new_n862), .ZN(RLL_wire_A_116));
  XOR2_X1 RLL_XOR_116 (.A(RLL_wire_A_116), .B(KEYINPUT116), .Z(new_n863) );
  OAI22_X1  g502(.A1(new_n840), .A2(new_n859), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g503(.A(new_n809), .B1(new_n828), .B2(new_n829), .ZN(new_n865));
  NOR3_X1   g504(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n866));
  NOR2_X1   g505(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI22_X1  g506(.A1(new_n867), .A2(new_n832), .B1(new_n825), .B2(new_n826), .ZN(new_n868));
  OAI21_X1  g507(.A(new_n838), .B1(new_n868), .B2(new_n841), .ZN(new_n869));
  AND3_X1   g508(.A1(new_n845), .A2(new_n848), .A3(new_n858), .ZN(new_n870));
  OAI21_X1  g509(.A(new_n809), .B1(new_n828), .B2(KEYINPUT45), .ZN(new_n871));
  NOR3_X1   g510(.A1(G164), .A2(new_n807), .A3(G1384), .ZN(new_n872));
  OAI21_X1  g511(.A(new_n672), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g512(.A(G2084), .ZN(new_n874));
  NAND4_X1  g513(.A1(new_n830), .A2(new_n831), .A3(new_n874), .A4(new_n809), .ZN(new_n875));
  AOI211_X1 g514(.A(new_n841), .B(G286), .C1(new_n873), .C2(new_n875), .ZN(new_n876));
  NAND4_X1  g515(.A1(new_n869), .A2(new_n840), .A3(new_n870), .A4(new_n876), .ZN(new_n877));
  INV_X1    g516(.A(KEYINPUT63), .ZN(new_n878));
  NAND2_X1  g517(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g518(.A1(new_n834), .A2(G8), .ZN(new_n880));
  AOI21_X1  g519(.A(new_n859), .B1(new_n880), .B2(new_n838), .ZN(new_n881));
  NAND4_X1  g520(.A1(new_n881), .A2(KEYINPUT63), .A3(new_n840), .A4(new_n876), .ZN(new_n882));
  AOI21_X1  g521(.A(new_n864), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  INV_X1    g522(.A(G1956), .ZN(new_n884));
  OAI21_X1  g523(.A(new_n884), .B1(new_n865), .B2(new_n866), .ZN(new_n885));
  INV_X1    g524(.A(KEYINPUT57), .ZN(new_n886));
  AND2_X1   g525(.A1(new_n474), .A2(new_n476), .ZN(RLL_wire_A_117));
  XOR2_X1 RLL_XOR_117 (.A(RLL_wire_A_117), .B(KEYINPUT117), .Z(new_n887) );
  NAND2_X1  g526(.A1(new_n484), .A2(new_n479), .ZN(new_n888));
  OAI21_X1  g527(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(RLL_wire_A_118));
  XOR2_X1 RLL_XOR_118 (.A(RLL_wire_A_118), .B(KEYINPUT118), .Z(new_n889) );
  NAND4_X1  g528(.A1(new_n477), .A2(KEYINPUT57), .A3(new_n479), .A4(new_n484), .ZN(new_n890));
  NAND2_X1  g529(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g530(.A(KEYINPUT56), .B(G2072), .ZN(new_n892));
  NAND4_X1  g531(.A1(new_n823), .A2(new_n824), .A3(new_n809), .A4(new_n892), .ZN(new_n893));
  AND3_X1   g532(.A1(new_n885), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g533(.A1(new_n809), .A2(new_n828), .ZN(new_n895));
  NOR2_X1   g534(.A1(new_n895), .A2(G2067), .ZN(new_n896));
  NAND3_X1  g535(.A1(new_n830), .A2(new_n831), .A3(new_n809), .ZN(new_n897));
  AOI21_X1  g536(.A(new_n896), .B1(new_n625), .B2(new_n897), .ZN(new_n898));
  OR2_X1    g537(.A1(new_n898), .A2(new_n514), .ZN(new_n899));
  NAND2_X1  g538(.A1(new_n885), .A2(new_n893), .ZN(new_n900));
  INV_X1    g539(.A(new_n891), .ZN(new_n901));
  NAND2_X1  g540(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g541(.A(new_n894), .B1(new_n899), .B2(new_n902), .ZN(RLL_wire_A_119));
  XOR2_X1 RLL_XOR_119 (.A(RLL_wire_A_119), .B(KEYINPUT119), .Z(new_n903) );
  INV_X1    g542(.A(G1996), .ZN(new_n904));
  NAND4_X1  g543(.A1(new_n823), .A2(new_n824), .A3(new_n904), .A4(new_n809), .ZN(new_n905));
  XOR2_X1   g544(.A(KEYINPUT58), .B(G1341), .Z(new_n906));
  NAND2_X1  g545(.A1(new_n895), .A2(new_n906), .ZN(RLL_wire_A_120));
  XNOR2_X1 RLL_XNOR_120 (.A(RLL_wire_A_120), .B(KEYINPUT120), .ZN(new_n907) );
  NAND2_X1  g546(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g547(.A1(new_n908), .A2(new_n467), .ZN(new_n909));
  NAND2_X1  g548(.A1(new_n909), .A2(KEYINPUT59), .ZN(new_n910));
  INV_X1    g549(.A(KEYINPUT59), .ZN(new_n911));
  NAND3_X1  g550(.A1(new_n908), .A2(new_n911), .A3(new_n467), .ZN(new_n912));
  NAND2_X1  g551(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g552(.A(KEYINPUT61), .ZN(new_n914));
  AOI21_X1  g553(.A(new_n891), .B1(new_n885), .B2(new_n893), .ZN(new_n915));
  OAI21_X1  g554(.A(new_n914), .B1(new_n894), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g555(.A1(new_n885), .A2(new_n891), .A3(new_n893), .ZN(new_n917));
  NAND3_X1  g556(.A1(new_n902), .A2(KEYINPUT61), .A3(new_n917), .ZN(new_n918));
  AND3_X1   g557(.A1(new_n913), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AND3_X1   g558(.A1(new_n898), .A2(KEYINPUT60), .A3(new_n514), .ZN(new_n920));
  AOI21_X1  g559(.A(new_n514), .B1(new_n898), .B2(KEYINPUT60), .ZN(new_n921));
  OAI22_X1  g560(.A1(new_n920), .A2(new_n921), .B1(KEYINPUT60), .B2(new_n898), .ZN(new_n922));
  AOI21_X1  g561(.A(new_n903), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g562(.A1(new_n873), .A2(new_n875), .ZN(new_n924));
  NOR2_X1   g563(.A1(G168), .A2(new_n841), .ZN(RLL_wire_A_121));
  XOR2_X1 RLL_XOR_121 (.A(RLL_wire_A_121), .B(KEYINPUT121), .Z(new_n925) );
  NAND2_X1  g564(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n927));
  NAND2_X1  g566(.A1(new_n924), .A2(G8), .ZN(new_n928));
  INV_X1    g567(.A(new_n925), .ZN(RLL_wire_A_122));
  XNOR2_X1 RLL_XNOR_122 (.A(RLL_wire_A_122), .B(KEYINPUT122), .ZN(new_n929) );
  AOI21_X1  g568(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g569(.A(new_n841), .B1(new_n873), .B2(new_n875), .ZN(new_n931));
  NOR3_X1   g570(.A1(new_n931), .A2(KEYINPUT51), .A3(new_n925), .ZN(new_n932));
  OAI21_X1  g571(.A(new_n926), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n934));
  NOR3_X1   g573(.A1(new_n871), .A2(new_n872), .A3(G2078), .ZN(new_n935));
  INV_X1    g574(.A(G1961), .ZN(new_n936));
  AOI22_X1  g575(.A1(new_n935), .A2(KEYINPUT53), .B1(new_n936), .B2(new_n897), .ZN(new_n937));
  INV_X1    g576(.A(KEYINPUT53), .ZN(RLL_wire_A_123));
  XNOR2_X1 RLL_XNOR_123 (.A(RLL_wire_A_123), .B(KEYINPUT123), .ZN(new_n938) );
  OAI21_X1  g577(.A(new_n938), .B1(new_n825), .B2(G2078), .ZN(new_n939));
  AOI21_X1  g578(.A(G301), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g579(.A1(new_n897), .A2(new_n936), .ZN(new_n941));
  INV_X1    g580(.A(new_n408), .ZN(new_n942));
  AND2_X1   g581(.A1(new_n398), .A2(new_n399), .ZN(new_n943));
  OAI211_X1 g582(.A(G40), .B(new_n942), .C1(new_n943), .C2(new_n396), .ZN(new_n944));
  AOI21_X1  g583(.A(new_n944), .B1(new_n806), .B2(new_n807), .ZN(new_n945));
  INV_X1    g584(.A(G2078), .ZN(new_n946));
  NAND4_X1  g585(.A1(new_n945), .A2(KEYINPUT53), .A3(new_n946), .A4(new_n824), .ZN(new_n947));
  AND4_X1   g586(.A1(G301), .A2(new_n939), .A3(new_n941), .A4(new_n947), .ZN(new_n948));
  OAI21_X1  g587(.A(new_n934), .B1(new_n940), .B2(new_n948), .ZN(RLL_wire_A_124));
  XOR2_X1 RLL_XOR_124 (.A(RLL_wire_A_124), .B(KEYINPUT124), .Z(new_n949) );
  AND3_X1   g588(.A1(new_n869), .A2(new_n840), .A3(new_n870), .ZN(new_n950));
  NAND3_X1  g589(.A1(new_n937), .A2(G301), .A3(new_n939), .ZN(new_n951));
  NAND3_X1  g590(.A1(new_n939), .A2(new_n947), .A3(new_n941), .ZN(new_n952));
  NAND2_X1  g591(.A1(new_n952), .A2(G171), .ZN(new_n953));
  NAND3_X1  g592(.A1(new_n951), .A2(new_n953), .A3(KEYINPUT54), .ZN(new_n954));
  NAND4_X1  g593(.A1(new_n933), .A2(new_n949), .A3(new_n950), .A4(new_n954), .ZN(new_n955));
  OAI21_X1  g594(.A(new_n883), .B1(new_n923), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g595(.A(new_n940), .B(new_n950), .C1(new_n933), .C2(KEYINPUT62), .ZN(RLL_wire_A_125));
  XOR2_X1 RLL_XOR_125 (.A(RLL_wire_A_125), .B(KEYINPUT125), .Z(new_n957) );
  AND2_X1   g596(.A1(new_n933), .A2(KEYINPUT62), .ZN(new_n958));
  NOR2_X1   g597(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g598(.A(new_n822), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g599(.A1(new_n594), .A2(new_n596), .ZN(new_n961));
  OAI22_X1  g600(.A1(new_n820), .A2(new_n961), .B1(G2067), .B2(new_n634), .ZN(new_n962));
  AND2_X1   g601(.A1(new_n962), .A2(new_n816), .ZN(new_n963));
  OR2_X1    g602(.A1(new_n814), .A2(KEYINPUT46), .ZN(new_n964));
  NAND2_X1  g603(.A1(new_n814), .A2(KEYINPUT46), .ZN(new_n965));
  OAI21_X1  g604(.A(new_n816), .B1(new_n818), .B2(new_n663), .ZN(new_n966));
  NAND3_X1  g605(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  XOR2_X1   g606(.A(new_n967), .B(KEYINPUT47), .Z(new_n968));
  AOI21_X1  g607(.A(new_n820), .B1(new_n816), .B2(new_n821), .ZN(RLL_wire_A_126));
  XOR2_X1 RLL_XOR_126 (.A(RLL_wire_A_126), .B(KEYINPUT126), .Z(new_n969) );
  NOR2_X1   g608(.A1(new_n811), .A2(new_n810), .ZN(RLL_wire_A_127));
  XNOR2_X1 RLL_XNOR_127 (.A(RLL_wire_A_127), .B(KEYINPUT127), .ZN(new_n970) );
  XOR2_X1   g609(.A(new_n970), .B(KEYINPUT48), .Z(new_n971));
  AOI211_X1 g610(.A(new_n963), .B(new_n968), .C1(new_n969), .C2(new_n971), .ZN(new_n972));
  NAND2_X1  g611(.A1(new_n960), .A2(new_n972), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g612(.A1(G227), .A2(new_n394), .ZN(new_n975));
  NAND2_X1  g613(.A1(new_n555), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g614(.A1(G229), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g615(.A(new_n750), .B(new_n977), .C1(new_n792), .C2(new_n798), .ZN(G225));
  INV_X1    g616(.A(G225), .ZN(G308));

endmodule
