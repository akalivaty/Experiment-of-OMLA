//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(G1gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT95), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n204), .B(new_n205), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n210), .B1(new_n209), .B2(new_n208), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT96), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n204), .A2(new_n208), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G8gat), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT93), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT15), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(new_n218), .B2(new_n217), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  OR3_X1    g020(.A1(new_n221), .A2(G29gat), .A3(G36gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G29gat), .A2(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT94), .B(G43gat), .Z(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G50gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(G43gat), .B2(new_n230), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n225), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n227), .B1(new_n234), .B2(new_n220), .ZN(new_n235));
  OR2_X1    g034(.A1(new_n216), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(KEYINPUT17), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n235), .A2(KEYINPUT17), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n216), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(KEYINPUT18), .A3(new_n241), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n216), .A2(new_n235), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n236), .A2(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n241), .B(KEYINPUT13), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(G113gat), .B(G141gat), .Z(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT92), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n253));
  XNOR2_X1  g052(.A(G169gat), .B(G197gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n252), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT12), .Z(new_n257));
  OR2_X1    g056(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n250), .A2(new_n257), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT21), .ZN(new_n261));
  XNOR2_X1  g060(.A(G57gat), .B(G64gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G71gat), .B(G78gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n216), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT99), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G127gat), .B(G155gat), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n268), .B(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G231gat), .A2(G233gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT98), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G183gat), .B(G211gat), .Z(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n273), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G85gat), .A2(G92gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT7), .ZN(new_n282));
  NAND2_X1  g081(.A1(G99gat), .A2(G106gat), .ZN(new_n283));
  INV_X1    g082(.A(G85gat), .ZN(new_n284));
  INV_X1    g083(.A(G92gat), .ZN(new_n285));
  AOI22_X1  g084(.A1(KEYINPUT8), .A2(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G99gat), .B(G106gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT101), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n238), .A2(new_n237), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G232gat), .A2(G233gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n292), .B(KEYINPUT100), .Z(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT41), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n291), .B(new_n295), .C1(new_n235), .C2(new_n290), .ZN(new_n296));
  XOR2_X1   g095(.A(G134gat), .B(G162gat), .Z(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n294), .A2(KEYINPUT41), .ZN(new_n299));
  XNOR2_X1  g098(.A(G190gat), .B(G218gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n301), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n280), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n289), .B(new_n266), .Z(new_n307));
  INV_X1    g106(.A(new_n266), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT10), .ZN(new_n309));
  OAI22_X1  g108(.A1(new_n307), .A2(KEYINPUT10), .B1(new_n290), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n310), .B(KEYINPUT102), .Z(new_n311));
  NAND2_X1  g110(.A1(G230gat), .A2(G233gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n307), .A2(G230gat), .A3(G233gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n314), .B(KEYINPUT103), .Z(new_n315));
  XNOR2_X1  g114(.A(G120gat), .B(G148gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(G176gat), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n317), .B(G204gat), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n310), .A2(new_n312), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n319), .B1(new_n315), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n306), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT89), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT25), .ZN(new_n327));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT65), .ZN(new_n329));
  NOR2_X1   g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330));
  OR2_X1    g129(.A1(new_n330), .A2(KEYINPUT23), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(KEYINPUT23), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT24), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n336), .A2(G183gat), .A3(G190gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT66), .B(G190gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(G183gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n333), .B1(KEYINPUT67), .B2(new_n340), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n340), .A2(KEYINPUT67), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n327), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n339), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT27), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n346), .B1(new_n347), .B2(G183gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT27), .B(G183gat), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n345), .B(new_n348), .C1(new_n346), .C2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n349), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n353), .A2(new_n351), .A3(new_n339), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n330), .B(KEYINPUT26), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n329), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n334), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT64), .ZN(new_n361));
  OR3_X1    g160(.A1(new_n361), .A2(G183gat), .A3(G190gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n361), .B1(G183gat), .B2(G190gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n338), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n333), .A2(KEYINPUT25), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n356), .A2(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G113gat), .ZN(new_n367));
  INV_X1    g166(.A(G120gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT1), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(G113gat), .B2(G120gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G127gat), .B(G134gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G127gat), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n375), .A2(G134gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(G134gat), .ZN(new_n377));
  OAI22_X1  g176(.A1(new_n369), .A2(new_n371), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n344), .A2(new_n366), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n379), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n364), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n354), .B1(new_n351), .B2(new_n350), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(new_n359), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n381), .B1(new_n384), .B2(new_n343), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G227gat), .ZN(new_n387));
  INV_X1    g186(.A(G233gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT32), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G71gat), .B(G99gat), .Z(new_n392));
  XNOR2_X1  g191(.A(G15gat), .B(G43gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n390), .B1(new_n380), .B2(new_n385), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n391), .B(new_n394), .C1(KEYINPUT33), .C2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n390), .A3(new_n385), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n397), .B(KEYINPUT34), .Z(new_n398));
  INV_X1    g197(.A(KEYINPUT32), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n394), .A2(KEYINPUT33), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT69), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT69), .ZN(new_n403));
  INV_X1    g202(.A(new_n401), .ZN(new_n404));
  NOR4_X1   g203(.A1(new_n395), .A2(new_n403), .A3(new_n399), .A4(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n396), .B(new_n398), .C1(new_n402), .C2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n403), .B1(new_n391), .B2(new_n404), .ZN(new_n408));
  INV_X1    g207(.A(new_n405), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n398), .B1(new_n410), .B2(new_n396), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n326), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT35), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n396), .B1(new_n402), .B2(new_n405), .ZN(new_n414));
  INV_X1    g213(.A(new_n398), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(KEYINPUT89), .A3(new_n406), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n384), .A2(new_n343), .ZN(new_n418));
  NAND2_X1  g217(.A1(G226gat), .A2(G233gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT71), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n344), .A2(new_n366), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT71), .B1(new_n384), .B2(new_n343), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT72), .B(KEYINPUT29), .Z(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(new_n419), .B(KEYINPUT70), .Z(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n420), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G197gat), .B(G204gat), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT22), .ZN(new_n431));
  INV_X1    g230(.A(G211gat), .ZN(new_n432));
  INV_X1    g231(.A(G218gat), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G211gat), .B(G218gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n430), .A3(new_n434), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n429), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n419), .B1(new_n418), .B2(KEYINPUT29), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(new_n440), .ZN(new_n445));
  XNOR2_X1  g244(.A(G8gat), .B(G36gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(G64gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(new_n285), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n442), .A2(KEYINPUT30), .A3(new_n445), .A4(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n445), .B1(new_n428), .B2(new_n440), .ZN(new_n450));
  INV_X1    g249(.A(new_n448), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n450), .B2(new_n451), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n449), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n412), .A2(new_n413), .A3(new_n417), .A4(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(G22gat), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n459));
  INV_X1    g258(.A(G228gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n460), .A2(new_n388), .ZN(new_n461));
  XNOR2_X1  g260(.A(G141gat), .B(G148gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT73), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT2), .ZN(new_n464));
  INV_X1    g263(.A(G141gat), .ZN(new_n465));
  INV_X1    g264(.A(G148gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT73), .ZN(new_n468));
  NAND2_X1  g267(.A1(G141gat), .A2(G148gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n463), .A2(new_n464), .A3(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(G155gat), .A2(G162gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT74), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n472), .B2(new_n473), .ZN(new_n477));
  INV_X1    g276(.A(G155gat), .ZN(new_n478));
  INV_X1    g277(.A(G162gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT74), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n464), .B1(G155gat), .B2(G162gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n462), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n483), .A2(KEYINPUT75), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT75), .B1(new_n483), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n475), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT29), .B1(new_n438), .B2(new_n439), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n488), .B1(KEYINPUT3), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT82), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n483), .A2(new_n485), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT75), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n483), .A2(KEYINPUT75), .A3(new_n485), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n440), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT3), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n497), .A2(new_n475), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(KEYINPUT82), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n461), .B1(new_n492), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n500), .B(new_n475), .C1(new_n486), .C2(new_n487), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n424), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT83), .B1(new_n505), .B2(new_n441), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT83), .ZN(new_n507));
  AOI211_X1 g306(.A(new_n507), .B(new_n440), .C1(new_n504), .C2(new_n424), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n459), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n505), .A2(new_n441), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n507), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n505), .A2(KEYINPUT83), .A3(new_n441), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n461), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n490), .A2(new_n491), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT82), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(KEYINPUT84), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n510), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n474), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT2), .B1(new_n462), .B2(KEYINPUT73), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(new_n470), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n495), .B2(new_n496), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT3), .B1(new_n440), .B2(new_n424), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n461), .B1(new_n511), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n458), .B1(new_n520), .B2(new_n528), .ZN(new_n529));
  AOI211_X1 g328(.A(G22gat), .B(new_n527), .C1(new_n510), .C2(new_n519), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT86), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n503), .A2(new_n509), .A3(new_n459), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT84), .B1(new_n514), .B2(new_n518), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n528), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G22gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT86), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n458), .A3(new_n528), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G78gat), .B(G106gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(new_n230), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n541));
  XOR2_X1   g340(.A(new_n540), .B(new_n541), .Z(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT85), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n543), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n531), .A2(new_n538), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT79), .ZN(new_n549));
  XOR2_X1   g348(.A(G1gat), .B(G29gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G57gat), .B(G85gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT5), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n475), .B(new_n379), .C1(new_n486), .C2(new_n487), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT4), .ZN(new_n556));
  NAND2_X1  g355(.A1(G225gat), .A2(G233gat), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n379), .B1(new_n488), .B2(KEYINPUT3), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n504), .ZN(new_n559));
  AND4_X1   g358(.A1(new_n554), .A2(new_n556), .A3(new_n557), .A4(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT77), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT76), .B1(new_n555), .B2(KEYINPUT4), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT76), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT4), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n524), .A2(new_n563), .A3(new_n564), .A4(new_n379), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n555), .A2(KEYINPUT4), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n381), .B1(new_n524), .B2(new_n500), .ZN(new_n568));
  INV_X1    g367(.A(new_n504), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n557), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n561), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n572), .A2(new_n559), .A3(KEYINPUT77), .A4(new_n557), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n488), .A2(new_n381), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n555), .ZN(new_n576));
  INV_X1    g375(.A(new_n557), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n554), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n560), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT87), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n578), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n582), .B1(new_n571), .B2(new_n573), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n583), .A2(KEYINPUT87), .A3(new_n560), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n553), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n553), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT6), .B1(new_n579), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n579), .A2(new_n586), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n585), .A2(new_n587), .B1(KEYINPUT6), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n545), .B1(new_n531), .B2(new_n538), .ZN(new_n590));
  NOR4_X1   g389(.A1(new_n457), .A2(new_n547), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT80), .B1(new_n579), .B2(new_n586), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT80), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n593), .B(new_n553), .C1(new_n583), .C2(new_n560), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n587), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n588), .A2(KEYINPUT6), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n455), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n542), .B1(new_n530), .B2(KEYINPUT85), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT86), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n407), .A2(new_n411), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n597), .A2(new_n601), .A3(new_n602), .A4(new_n546), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT35), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT90), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT90), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n603), .A2(new_n606), .A3(KEYINPUT35), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n591), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n442), .A2(new_n445), .A3(new_n448), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT37), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n610), .B(new_n445), .C1(new_n428), .C2(new_n440), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n611), .A2(KEYINPUT88), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n450), .A2(KEYINPUT37), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n448), .B1(new_n611), .B2(KEYINPUT88), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT38), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n429), .A2(new_n440), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n443), .A2(new_n444), .A3(new_n441), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n618), .A2(KEYINPUT37), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT38), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n612), .A2(new_n620), .A3(new_n614), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n589), .A2(new_n609), .A3(new_n616), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n547), .A2(new_n590), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n557), .B1(new_n556), .B2(new_n559), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n553), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT39), .B1(new_n576), .B2(new_n577), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT40), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n585), .A2(new_n455), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n622), .A2(new_n623), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n595), .A2(new_n596), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI22_X1  g432(.A1(new_n633), .A2(new_n455), .B1(new_n547), .B2(new_n590), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT36), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n407), .B2(new_n411), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n416), .A2(KEYINPUT36), .A3(new_n406), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n631), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n260), .B(new_n325), .C1(new_n608), .C2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n632), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n203), .ZN(G1324gat));
  OAI21_X1  g442(.A(G8gat), .B1(new_n641), .B2(new_n456), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT104), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT16), .B(G8gat), .ZN(new_n647));
  OR3_X1    g446(.A1(new_n641), .A2(new_n456), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT42), .Z(new_n649));
  OR3_X1    g448(.A1(new_n646), .A2(new_n649), .A3(KEYINPUT105), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT105), .B1(new_n646), .B2(new_n649), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(G1325gat));
  AND3_X1   g451(.A1(new_n636), .A2(KEYINPUT106), .A3(new_n637), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT106), .B1(new_n636), .B2(new_n637), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(G15gat), .B1(new_n641), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n412), .A2(new_n417), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(G15gat), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n641), .B2(new_n658), .ZN(G1326gat));
  NOR2_X1   g458(.A1(new_n641), .A2(new_n623), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT43), .B(G22gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT107), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n660), .B(new_n662), .ZN(G1327gat));
  INV_X1    g462(.A(new_n280), .ZN(new_n664));
  INV_X1    g463(.A(new_n324), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n305), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n667), .B(new_n260), .C1(new_n608), .C2(new_n640), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n668), .A2(G29gat), .A3(new_n632), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT45), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n304), .A2(KEYINPUT44), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n608), .B2(new_n640), .ZN(new_n673));
  INV_X1    g472(.A(new_n260), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n657), .A2(new_n455), .ZN(new_n676));
  INV_X1    g475(.A(new_n589), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n676), .A2(new_n623), .A3(new_n413), .A4(new_n677), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n603), .A2(new_n606), .A3(KEYINPUT35), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n606), .B1(new_n603), .B2(KEYINPUT35), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n631), .A2(new_n655), .A3(new_n634), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n305), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n673), .B(new_n675), .C1(new_n683), .C2(KEYINPUT44), .ZN(new_n684));
  OAI21_X1  g483(.A(G29gat), .B1(new_n684), .B2(new_n632), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n685), .ZN(G1328gat));
  NOR3_X1   g485(.A1(new_n668), .A2(G36gat), .A3(new_n456), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT46), .ZN(new_n688));
  OAI21_X1  g487(.A(G36gat), .B1(new_n684), .B2(new_n456), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1329gat));
  NOR2_X1   g489(.A1(new_n657), .A2(new_n229), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OR3_X1    g491(.A1(new_n668), .A2(KEYINPUT108), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT108), .B1(new_n668), .B2(new_n692), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n229), .B1(new_n684), .B2(new_n655), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n700), .B1(new_n684), .B2(new_n655), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n671), .B1(new_n681), .B2(new_n639), .ZN(new_n702));
  INV_X1    g501(.A(new_n682), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n304), .B1(new_n608), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n655), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n706), .A2(KEYINPUT109), .A3(new_n707), .A4(new_n675), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n701), .A2(new_n708), .A3(new_n229), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n698), .B1(new_n693), .B2(new_n694), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n709), .A2(KEYINPUT110), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT110), .B1(new_n709), .B2(new_n710), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n699), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT111), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n699), .B(new_n715), .C1(new_n711), .C2(new_n712), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1330gat));
  OAI21_X1  g516(.A(G50gat), .B1(new_n684), .B2(new_n623), .ZN(new_n718));
  INV_X1    g517(.A(new_n623), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n230), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n668), .B2(new_n720), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g521(.A1(new_n681), .A2(new_n682), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n306), .A2(new_n260), .A3(new_n665), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n633), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT112), .B(G57gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1332gat));
  INV_X1    g527(.A(new_n725), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n456), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(G1333gat));
  NAND3_X1  g533(.A1(new_n725), .A2(G71gat), .A3(new_n707), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT113), .Z(new_n736));
  INV_X1    g535(.A(KEYINPUT114), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n729), .A2(new_n737), .A3(new_n657), .ZN(new_n738));
  INV_X1    g537(.A(new_n657), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT114), .B1(new_n725), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n738), .A2(G71gat), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g542(.A1(new_n725), .A2(new_n719), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g544(.A1(new_n260), .A2(new_n280), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n683), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT51), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n665), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n284), .A3(new_n633), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n706), .A2(new_n324), .A3(new_n746), .ZN(new_n751));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751), .B2(new_n632), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1336gat));
  OAI21_X1  g552(.A(G92gat), .B1(new_n751), .B2(new_n456), .ZN(new_n754));
  NAND2_X1  g553(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n324), .A2(new_n285), .A3(new_n455), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n756), .B(KEYINPUT115), .Z(new_n757));
  OAI211_X1 g556(.A(new_n754), .B(new_n755), .C1(new_n748), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT116), .A2(KEYINPUT52), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT117), .Z(new_n760));
  XNOR2_X1  g559(.A(new_n758), .B(new_n760), .ZN(G1337gat));
  INV_X1    g560(.A(G99gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n749), .A2(new_n762), .A3(new_n739), .ZN(new_n763));
  OAI21_X1  g562(.A(G99gat), .B1(new_n751), .B2(new_n655), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1338gat));
  INV_X1    g564(.A(G106gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n766), .A3(new_n719), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G106gat), .B1(new_n751), .B2(new_n623), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(new_n771), .A3(KEYINPUT53), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n767), .B(new_n770), .C1(new_n768), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1339gat));
  NAND2_X1  g574(.A1(new_n325), .A2(new_n674), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n313), .B(KEYINPUT54), .C1(new_n312), .C2(new_n310), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n318), .B1(new_n322), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT55), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n321), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n674), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n240), .A2(new_n241), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n247), .A2(new_n248), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n256), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n258), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n305), .B1(new_n790), .B2(new_n665), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n304), .B1(new_n785), .B2(new_n790), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n664), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n776), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n623), .A2(new_n602), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n633), .A2(new_n456), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n795), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(G113gat), .B1(new_n801), .B2(new_n260), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n795), .A2(new_n623), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(new_n633), .A3(new_n676), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n674), .A2(new_n367), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n802), .B1(new_n805), .B2(new_n806), .ZN(G1340gat));
  AOI21_X1  g606(.A(G120gat), .B1(new_n801), .B2(new_n324), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n665), .A2(new_n368), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n805), .B2(new_n809), .ZN(G1341gat));
  OAI21_X1  g609(.A(G127gat), .B1(new_n804), .B2(new_n664), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n801), .A2(new_n375), .A3(new_n280), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1342gat));
  NOR3_X1   g612(.A1(new_n800), .A2(G134gat), .A3(new_n305), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n815), .A2(KEYINPUT56), .ZN(new_n816));
  OAI21_X1  g615(.A(G134gat), .B1(new_n804), .B2(new_n305), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(KEYINPUT56), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(G1343gat));
  NAND2_X1  g618(.A1(new_n795), .A2(new_n719), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n820), .A2(new_n707), .A3(new_n798), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n465), .A3(new_n260), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823));
  XNOR2_X1  g622(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n781), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n825), .A2(new_n321), .A3(new_n782), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n791), .B1(new_n826), .B2(new_n260), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828));
  OR3_X1    g627(.A1(new_n794), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n827), .B2(new_n794), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n776), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n823), .B1(new_n831), .B2(new_n719), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n707), .A2(new_n798), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n820), .B2(KEYINPUT57), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n832), .A2(new_n834), .A3(new_n674), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n822), .B1(new_n835), .B2(new_n465), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n466), .A3(new_n324), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n820), .A2(KEYINPUT57), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n776), .B1(new_n827), .B2(new_n794), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n823), .A3(new_n719), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n324), .A3(new_n833), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n466), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n839), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n834), .ZN(new_n849));
  AOI211_X1 g648(.A(KEYINPUT59), .B(new_n466), .C1(new_n849), .C2(new_n324), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n838), .B1(new_n848), .B2(new_n850), .ZN(G1345gat));
  AOI21_X1  g650(.A(G155gat), .B1(new_n821), .B2(new_n280), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n280), .A2(G155gat), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(KEYINPUT122), .Z(new_n854));
  AOI21_X1  g653(.A(new_n852), .B1(new_n849), .B2(new_n854), .ZN(G1346gat));
  NAND3_X1  g654(.A1(new_n821), .A2(new_n479), .A3(new_n304), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n832), .A2(new_n834), .A3(new_n305), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n479), .ZN(G1347gat));
  NAND4_X1  g657(.A1(new_n803), .A2(new_n632), .A3(new_n455), .A4(new_n739), .ZN(new_n859));
  INV_X1    g658(.A(G169gat), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n859), .A2(new_n860), .A3(new_n674), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n796), .A2(new_n456), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n795), .A2(new_n632), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT123), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(KEYINPUT123), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n260), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n861), .B1(new_n868), .B2(new_n860), .ZN(G1348gat));
  OAI21_X1  g668(.A(G176gat), .B1(new_n859), .B2(new_n665), .ZN(new_n870));
  INV_X1    g669(.A(new_n867), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n665), .A2(G176gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(G1349gat));
  NOR2_X1   g672(.A1(new_n664), .A2(new_n353), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT125), .B1(new_n867), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n859), .B2(new_n664), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(G183gat), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n859), .A2(new_n876), .A3(new_n664), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n875), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g680(.A1(new_n867), .A2(new_n345), .A3(new_n304), .ZN(new_n882));
  OAI21_X1  g681(.A(G190gat), .B1(new_n859), .B2(new_n305), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(KEYINPUT61), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(KEYINPUT61), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(G1351gat));
  NAND2_X1  g685(.A1(new_n865), .A2(new_n866), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n707), .A2(new_n456), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n623), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n674), .A2(G197gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT126), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n889), .A2(new_n633), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n843), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n260), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G197gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n893), .A2(new_n897), .ZN(G1352gat));
  AND2_X1   g697(.A1(new_n887), .A2(new_n890), .ZN(new_n899));
  XOR2_X1   g698(.A(KEYINPUT127), .B(G204gat), .Z(new_n900));
  NOR2_X1   g699(.A1(new_n665), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(KEYINPUT62), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n843), .A2(new_n324), .A3(new_n894), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n900), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(KEYINPUT62), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(G1353gat));
  NAND3_X1  g706(.A1(new_n899), .A2(new_n432), .A3(new_n280), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n895), .A2(new_n280), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT63), .B1(new_n909), .B2(G211gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1354gat));
  AOI21_X1  g711(.A(G218gat), .B1(new_n899), .B2(new_n304), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n305), .A2(new_n433), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n895), .B2(new_n914), .ZN(G1355gat));
endmodule


