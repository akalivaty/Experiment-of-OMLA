//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1126, new_n1127;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n452), .A2(G2106), .B1(KEYINPUT66), .B2(new_n458), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n464), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n476), .A2(new_n477), .A3(new_n478), .A4(new_n467), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n471), .B(new_n473), .C1(new_n474), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT68), .ZN(G160));
  XNOR2_X1  g056(.A(new_n479), .B(KEYINPUT69), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n478), .A2(G100), .ZN(new_n484));
  NAND2_X1  g059(.A1(G112), .A2(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n466), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND4_X1   g061(.A1(G2105), .A2(new_n476), .A3(new_n477), .A4(new_n467), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G124), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  MUX2_X1   g066(.A(G102), .B(G114), .S(G2105), .Z(new_n492));
  AOI22_X1  g067(.A1(new_n487), .A2(G126), .B1(G2104), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  OAI211_X1 g069(.A(KEYINPUT70), .B(KEYINPUT4), .C1(new_n479), .C2(new_n494), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(new_n465), .A3(new_n467), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT67), .B1(new_n464), .B2(G2104), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n464), .A2(G2104), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n501), .A2(G138), .A3(new_n478), .A4(new_n477), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT70), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n491), .B(new_n493), .C1(new_n498), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n479), .B2(new_n494), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(new_n495), .A3(new_n497), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n491), .B1(new_n509), .B2(new_n493), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n505), .A2(new_n510), .ZN(G164));
  AND3_X1   g086(.A1(KEYINPUT72), .A2(KEYINPUT6), .A3(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT6), .B1(KEYINPUT72), .B2(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI21_X1  g093(.A(G543), .B1(new_n512), .B2(new_n513), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n520), .A2(new_n523), .ZN(G166));
  INV_X1    g099(.A(new_n516), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n528), .B(new_n529), .C1(new_n530), .C2(new_n519), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n526), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(new_n515), .A2(G64), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n522), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n537), .B1(new_n536), .B2(new_n535), .ZN(new_n538));
  INV_X1    g113(.A(new_n519), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n525), .A2(G90), .B1(G52), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n516), .A2(new_n543), .B1(new_n544), .B2(new_n519), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n522), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n525), .A2(G91), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(KEYINPUT74), .A2(G53), .ZN(new_n557));
  OR3_X1    g132(.A1(new_n519), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n522), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n556), .B1(new_n519), .B2(new_n557), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n555), .A2(new_n558), .A3(new_n560), .A4(new_n561), .ZN(G299));
  XNOR2_X1  g137(.A(G168), .B(KEYINPUT75), .ZN(G286));
  INV_X1    g138(.A(G166), .ZN(G303));
  NAND2_X1  g139(.A1(new_n525), .A2(G87), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n539), .A2(G49), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(new_n539), .A2(G48), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  OAI221_X1 g146(.A(new_n569), .B1(new_n570), .B2(new_n516), .C1(new_n522), .C2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n522), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g154(.A(KEYINPUT78), .B(G85), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n525), .A2(new_n580), .B1(G47), .B2(new_n539), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n579), .A2(KEYINPUT79), .A3(new_n581), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G290));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G301), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n522), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n514), .A2(KEYINPUT80), .A3(G543), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n519), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G54), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n589), .B(new_n592), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n597), .B1(new_n593), .B2(new_n595), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT81), .B1(new_n599), .B2(new_n591), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n516), .A2(new_n601), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n598), .A2(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n588), .B1(new_n587), .B2(new_n605), .ZN(G284));
  AOI21_X1  g181(.A(new_n588), .B1(new_n587), .B2(new_n605), .ZN(G321));
  NAND2_X1  g182(.A1(G299), .A2(new_n587), .ZN(new_n608));
  INV_X1    g183(.A(G286), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n587), .ZN(G297));
  XNOR2_X1  g185(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT83), .Z(G148));
  NOR3_X1   g189(.A1(new_n545), .A2(G868), .A3(new_n547), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n598), .A2(new_n600), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n603), .A2(new_n604), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(G559), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n615), .B1(new_n619), .B2(G868), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n487), .A2(G123), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT86), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n482), .A2(G135), .ZN(new_n624));
  MUX2_X1   g199(.A(G99), .B(G111), .S(G2105), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G2104), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n478), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT84), .B(G2100), .Z(new_n634));
  AOI22_X1  g209(.A1(new_n633), .A2(KEYINPUT13), .B1(KEYINPUT85), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(KEYINPUT13), .B2(new_n633), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n634), .A2(KEYINPUT85), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n627), .A2(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n630), .A2(new_n638), .A3(new_n639), .ZN(G156));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT15), .B(G2435), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2427), .ZN(new_n644));
  INV_X1    g219(.A(G2430), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n647), .A2(new_n653), .ZN(new_n655));
  AND3_X1   g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT88), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n657), .A2(new_n658), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n660), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n668), .B(new_n659), .C1(new_n669), .C2(new_n665), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n629), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n678), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT89), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n675), .A2(new_n679), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(KEYINPUT20), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(KEYINPUT20), .ZN(new_n685));
  AOI211_X1 g260(.A(new_n680), .B(new_n682), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT90), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT91), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n689), .B(new_n693), .ZN(G229));
  NOR2_X1   g269(.A1(G6), .A2(G16), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n574), .B2(G16), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT93), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT32), .B(G1981), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(G288), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G16), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(G16), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n699), .A2(new_n700), .A3(new_n706), .A4(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT34), .ZN(new_n713));
  NOR2_X1   g288(.A1(G16), .A2(G24), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n584), .A2(new_n585), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G16), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT92), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1986), .ZN(new_n718));
  NOR2_X1   g293(.A1(G25), .A2(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n482), .A2(G131), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n478), .A2(G95), .ZN(new_n721));
  NAND2_X1  g296(.A1(G107), .A2(G2105), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n466), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n487), .B2(G119), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n719), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  XOR2_X1   g303(.A(new_n727), .B(new_n728), .Z(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n712), .A2(new_n713), .A3(new_n718), .A4(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(KEYINPUT36), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(KEYINPUT36), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n701), .A2(G21), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G168), .B2(new_n701), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n736), .A2(G1966), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT31), .B(G11), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT96), .B(G28), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(KEYINPUT30), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n738), .B1(new_n740), .B2(new_n743), .C1(new_n736), .C2(G1966), .ZN(new_n744));
  AND2_X1   g319(.A1(KEYINPUT24), .A2(G34), .ZN(new_n745));
  NOR2_X1   g320(.A1(KEYINPUT24), .A2(G34), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G160), .B2(G29), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n737), .B(new_n744), .C1(new_n749), .C2(G2084), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n701), .A2(G5), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G171), .B2(new_n701), .ZN(new_n752));
  AOI22_X1  g327(.A1(G1961), .A2(new_n752), .B1(new_n628), .B2(G29), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n750), .B(new_n753), .C1(G1961), .C2(new_n752), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n701), .A2(G20), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT98), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT23), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G1956), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n742), .A2(G32), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n482), .A2(G141), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n472), .A2(G105), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT26), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n763), .B(new_n765), .C1(new_n487), .C2(G129), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n761), .B1(new_n768), .B2(new_n742), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT27), .B(G1996), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G4), .A2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n605), .B2(G16), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G1348), .ZN(new_n774));
  NOR2_X1   g349(.A1(G29), .A2(G35), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G162), .B2(G29), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT29), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n774), .B1(new_n777), .B2(G2090), .ZN(new_n778));
  NOR4_X1   g353(.A1(new_n754), .A2(new_n760), .A3(new_n771), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n742), .A2(G27), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G164), .B2(new_n742), .ZN(new_n781));
  INV_X1    g356(.A(G2078), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n773), .A2(G1348), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n749), .A2(G2084), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT97), .Z(new_n786));
  AOI211_X1 g361(.A(new_n784), .B(new_n786), .C1(G2090), .C2(new_n777), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G19), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n548), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT94), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1341), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n482), .A2(G139), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n465), .A2(new_n467), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n793), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n794));
  AOI21_X1  g369(.A(KEYINPUT25), .B1(new_n472), .B2(G103), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n792), .B1(new_n478), .B2(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G33), .B(new_n797), .S(G29), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2072), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n742), .A2(G26), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT28), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n482), .A2(G140), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n487), .A2(G128), .ZN(new_n803));
  NOR2_X1   g378(.A1(G104), .A2(G2105), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT95), .Z(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(new_n478), .B2(G116), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n802), .B(new_n803), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n801), .B1(new_n807), .B2(G29), .ZN(new_n808));
  INV_X1    g383(.A(G2067), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n791), .A2(new_n799), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n779), .A2(new_n783), .A3(new_n787), .A4(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n734), .A2(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  XOR2_X1   g392(.A(KEYINPUT100), .B(G93), .Z(new_n818));
  INV_X1    g393(.A(G55), .ZN(new_n819));
  OAI22_X1  g394(.A1(new_n516), .A2(new_n818), .B1(new_n819), .B2(new_n519), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT101), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n522), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n548), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n605), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT102), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n829));
  AOI21_X1  g404(.A(G860), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n829), .B2(new_n828), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n823), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(G145));
  XNOR2_X1  g409(.A(new_n725), .B(new_n632), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n482), .A2(G142), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n478), .A2(G106), .ZN(new_n837));
  NAND2_X1  g412(.A1(G118), .A2(G2105), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n466), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n487), .B2(G130), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n835), .B(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n493), .B1(new_n498), .B2(new_n503), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n807), .B(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n842), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n797), .B(new_n767), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(G160), .B(new_n489), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n627), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(G37), .B1(new_n847), .B2(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g428(.A(G290), .B(G288), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n574), .B(G303), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT42), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n857), .A2(KEYINPUT106), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(KEYINPUT106), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n856), .B2(new_n859), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n824), .B(new_n619), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n605), .A2(G299), .ZN(new_n863));
  INV_X1    g438(.A(G299), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT103), .B1(new_n618), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n605), .A2(new_n866), .A3(G299), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n863), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n865), .A2(new_n867), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n605), .A2(KEYINPUT104), .A3(G299), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT104), .B1(new_n605), .B2(G299), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n870), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT105), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n877), .B(new_n870), .C1(new_n871), .C2(new_n874), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n868), .A2(KEYINPUT41), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n880), .A2(new_n862), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n861), .B1(new_n869), .B2(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n882), .A2(KEYINPUT107), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n861), .A2(new_n881), .A3(new_n869), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n882), .B2(KEYINPUT107), .ZN(new_n885));
  OAI21_X1  g460(.A(G868), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n823), .A2(new_n587), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(G295));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n887), .ZN(G331));
  NAND2_X1  g464(.A1(G286), .A2(G171), .ZN(new_n890));
  NAND3_X1  g465(.A1(G301), .A2(KEYINPUT108), .A3(G168), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n892));
  INV_X1    g467(.A(G168), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(G171), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n890), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n824), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n878), .A2(new_n879), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(new_n876), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n896), .A2(new_n868), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n856), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n880), .A2(new_n896), .ZN(new_n903));
  INV_X1    g478(.A(new_n856), .ZN(new_n904));
  INV_X1    g479(.A(new_n900), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n901), .A2(new_n902), .A3(new_n906), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT44), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n900), .B1(new_n880), .B2(new_n896), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n910), .B2(new_n904), .ZN(new_n911));
  OR3_X1    g486(.A1(new_n868), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT109), .B1(new_n868), .B2(KEYINPUT41), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n871), .A2(new_n874), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n912), .B(new_n913), .C1(new_n870), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n896), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n905), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n856), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n902), .B1(new_n911), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT110), .B1(new_n909), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n906), .A2(new_n907), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n904), .B1(new_n916), .B2(new_n905), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT44), .A4(new_n908), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n902), .B1(new_n921), .B2(new_n922), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n911), .A2(KEYINPUT43), .A3(new_n901), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n926), .A2(new_n931), .ZN(G397));
  INV_X1    g507(.A(G40), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n480), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(G1384), .B1(new_n509), .B2(new_n493), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT45), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n807), .B(new_n809), .ZN(new_n938));
  INV_X1    g513(.A(G1996), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n767), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n725), .B(new_n728), .Z(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(G290), .B(G1986), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n937), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n935), .B1(KEYINPUT45), .B2(new_n936), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n843), .A2(KEYINPUT71), .ZN(new_n950));
  AOI21_X1  g525(.A(G1384), .B1(new_n950), .B2(new_n504), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n951), .B2(KEYINPUT45), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n949), .B(KEYINPUT111), .C1(new_n951), .C2(KEYINPUT45), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n954), .A2(new_n709), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n935), .B1(new_n957), .B2(new_n936), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n951), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT112), .B1(new_n959), .B2(G2090), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n505), .B2(new_n510), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT112), .ZN(new_n964));
  INV_X1    g539(.A(G2090), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n958), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n948), .B1(new_n956), .B2(new_n967), .ZN(new_n968));
  OAI211_X1 g543(.A(G303), .B(G8), .C1(KEYINPUT114), .C2(KEYINPUT55), .ZN(new_n969));
  NAND2_X1  g544(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n954), .A2(new_n709), .A3(new_n955), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n972), .A2(KEYINPUT113), .A3(new_n960), .A4(new_n966), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n968), .A2(G8), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n975));
  INV_X1    g550(.A(new_n971), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n936), .A2(KEYINPUT50), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n951), .B2(KEYINPUT50), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(new_n965), .A3(new_n934), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G8), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n975), .B(new_n976), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n972), .B2(new_n979), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT117), .B1(new_n983), .B2(new_n971), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n936), .A2(new_n934), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(new_n981), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n572), .B(G1981), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n989), .A2(KEYINPUT115), .A3(new_n988), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT115), .B1(new_n989), .B2(new_n988), .ZN(new_n991));
  OAI221_X1 g566(.A(new_n987), .B1(new_n988), .B2(new_n989), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n987), .ZN(new_n993));
  INV_X1    g568(.A(G1976), .ZN(new_n994));
  NOR2_X1   g569(.A1(G288), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT52), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(G288), .B2(new_n994), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n987), .B(new_n997), .C1(new_n994), .C2(G288), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n992), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n974), .A2(new_n982), .A3(new_n984), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1966), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n843), .A2(new_n961), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n935), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT45), .B(new_n961), .C1(new_n505), .C2(new_n510), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(KEYINPUT118), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n951), .B2(KEYINPUT45), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1001), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G2084), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n963), .A2(new_n1010), .A3(new_n958), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n981), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n609), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n947), .B1(new_n1000), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n968), .A2(G8), .A3(new_n973), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n976), .ZN(new_n1016));
  AND4_X1   g591(.A1(KEYINPUT63), .A2(new_n999), .A3(new_n609), .A4(new_n1012), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n974), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(G168), .A2(new_n981), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1009), .A2(KEYINPUT124), .A3(new_n1011), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT124), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n1024));
  OAI21_X1  g599(.A(G8), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1020), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1012), .A2(KEYINPUT51), .A3(new_n1020), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1023), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AND4_X1   g604(.A1(new_n974), .A2(new_n982), .A3(new_n984), .A4(new_n999), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT58), .B(G1341), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n986), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n934), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n1003), .B2(new_n962), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1034), .B2(new_n939), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT123), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n548), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT59), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  OAI22_X1  g613(.A1(new_n952), .A2(G1996), .B1(new_n986), .B2(new_n1031), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT59), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1039), .A2(new_n1036), .A3(new_n1040), .A4(new_n548), .ZN(new_n1041));
  INV_X1    g616(.A(G1348), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n959), .A2(new_n1042), .B1(new_n809), .B2(new_n986), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n618), .A2(KEYINPUT60), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1038), .A2(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT61), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1956), .B1(new_n978), .B2(new_n934), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT56), .B(G2072), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n949), .B(new_n1048), .C1(new_n951), .C2(KEYINPUT45), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT121), .B1(new_n864), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(G299), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(KEYINPUT57), .B2(new_n1052), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1047), .A2(new_n1050), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1057), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1002), .A2(new_n957), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n962), .B2(new_n957), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n759), .B1(new_n1061), .B2(new_n935), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1059), .B1(new_n1062), .B2(new_n1049), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1046), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1043), .A2(new_n618), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1043), .A2(new_n618), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT60), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1057), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1062), .A2(new_n1059), .A3(new_n1049), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(KEYINPUT61), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1045), .A2(new_n1064), .A3(new_n1067), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1069), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1072), .A2(KEYINPUT122), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(KEYINPUT122), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(G2078), .B1(new_n954), .B2(new_n955), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(KEYINPUT53), .ZN(new_n1077));
  INV_X1    g652(.A(G1961), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n1078), .B2(new_n959), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n782), .A2(KEYINPUT53), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(new_n936), .B2(KEYINPUT45), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1004), .A2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT125), .ZN(new_n1083));
  XNOR2_X1  g658(.A(G301), .B(KEYINPUT54), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n959), .A2(new_n1078), .ZN(new_n1086));
  OR3_X1    g661(.A1(new_n1006), .A2(new_n1008), .A3(new_n1080), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1086), .B(new_n1087), .C1(new_n1076), .C2(KEYINPUT53), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1079), .A2(new_n1085), .B1(new_n1088), .B2(new_n1084), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1029), .A2(new_n1030), .A3(new_n1075), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n992), .A2(new_n994), .A3(new_n703), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(G1981), .B2(new_n572), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n993), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1095));
  INV_X1    g670(.A(new_n974), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1094), .A2(new_n1095), .B1(new_n1096), .B2(new_n999), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1019), .A2(new_n1090), .A3(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1088), .A2(G171), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1030), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1029), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(KEYINPUT62), .B(new_n1023), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n946), .B1(new_n1098), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n937), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(G1996), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(KEYINPUT46), .ZN(new_n1108));
  XOR2_X1   g683(.A(new_n1108), .B(KEYINPUT126), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(KEYINPUT46), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT127), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1106), .B1(new_n938), .B2(new_n768), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(new_n1113), .B(KEYINPUT47), .Z(new_n1114));
  NAND2_X1  g689(.A1(new_n726), .A2(new_n728), .ZN(new_n1115));
  OAI22_X1  g690(.A1(new_n941), .A2(new_n1115), .B1(G2067), .B2(new_n807), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n937), .ZN(new_n1117));
  INV_X1    g692(.A(G1986), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n715), .A2(new_n1118), .A3(new_n937), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n944), .A2(new_n937), .B1(KEYINPUT48), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(KEYINPUT48), .B2(new_n1120), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1114), .A2(new_n1117), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1105), .A2(new_n1123), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g699(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1126));
  AND2_X1   g700(.A1(new_n852), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g701(.A1(new_n929), .A2(new_n1127), .ZN(G225));
  INV_X1    g702(.A(G225), .ZN(G308));
endmodule


