//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n462), .A2(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(KEYINPUT68), .A3(G101), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n467), .A2(G137), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  AND3_X1   g055(.A1(new_n463), .A2(new_n465), .A3(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n467), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND4_X1  g062(.A1(new_n463), .A2(new_n465), .A3(G126), .A4(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n466), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT3), .B(G2104), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n496), .A2(new_n497), .A3(G138), .A4(new_n466), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n495), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n502), .A2(new_n504), .B1(new_n501), .B2(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(G543), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n508), .A2(new_n514), .ZN(G166));
  AND2_X1   g090(.A1(new_n509), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G51), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n505), .A2(G89), .A3(new_n509), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n517), .A2(new_n518), .A3(new_n519), .A4(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n524));
  NAND2_X1  g099(.A1(G77), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n502), .A2(new_n504), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n501), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G64), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G651), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n526), .A2(G90), .A3(new_n527), .A4(new_n509), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n509), .A2(G52), .A3(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n524), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n505), .A2(G64), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n507), .B1(new_n537), .B2(new_n525), .ZN(new_n538));
  NOR3_X1   g113(.A1(new_n538), .A2(new_n534), .A3(KEYINPUT70), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND3_X1  g116(.A1(new_n505), .A2(G81), .A3(new_n509), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT71), .B(G43), .Z(new_n543));
  NAND2_X1  g118(.A1(new_n516), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n542), .B(new_n544), .C1(new_n545), .C2(new_n507), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  AND2_X1   g128(.A1(new_n505), .A2(new_n509), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT6), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n555), .A2(new_n557), .A3(G53), .A4(G543), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n509), .A2(new_n560), .A3(G53), .A4(G543), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n554), .A2(G91), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n503), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT69), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n564));
  OAI211_X1 g139(.A(G65), .B(new_n527), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(KEYINPUT72), .B1(new_n567), .B2(G651), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n569));
  AOI211_X1 g144(.A(new_n569), .B(new_n507), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n562), .B1(new_n568), .B2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G166), .ZN(G303));
  NAND4_X1  g147(.A1(new_n526), .A2(G87), .A3(new_n527), .A4(new_n509), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n509), .A2(G49), .A3(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(G74), .B1(new_n526), .B2(new_n527), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(new_n507), .ZN(G288));
  NAND2_X1  g151(.A1(new_n516), .A2(G48), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n505), .A2(G86), .A3(new_n509), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n526), .A2(G61), .A3(new_n527), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n507), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n579), .A2(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n507), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n510), .A2(new_n586), .B1(new_n587), .B2(new_n513), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n528), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G54), .B2(new_n516), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n505), .A2(G92), .A3(new_n509), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n505), .A2(KEYINPUT10), .A3(G92), .A4(new_n509), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G321));
  XOR2_X1   g178(.A(G321), .B(KEYINPUT73), .Z(G284));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n559), .A2(new_n561), .ZN(new_n606));
  INV_X1    g181(.A(G91), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n510), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n569), .B1(new_n609), .B2(new_n507), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n567), .A2(KEYINPUT72), .A3(G651), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G868), .ZN(G297));
  OAI21_X1  g188(.A(new_n605), .B1(new_n612), .B2(G868), .ZN(G280));
  AND2_X1   g189(.A1(new_n594), .A2(new_n599), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT74), .B(G559), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n615), .B1(G860), .B2(new_n617), .ZN(G148));
  NAND2_X1  g193(.A1(new_n546), .A2(new_n601), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n600), .A2(new_n616), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n601), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g197(.A1(new_n481), .A2(G123), .B1(new_n467), .B2(G135), .ZN(new_n623));
  NOR3_X1   g198(.A1(new_n466), .A2(KEYINPUT76), .A3(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT76), .B1(new_n466), .B2(G111), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n625), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n623), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n496), .A2(new_n472), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XOR2_X1   g205(.A(KEYINPUT75), .B(G2100), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT77), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT78), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT17), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n657), .B(KEYINPUT79), .Z(new_n660));
  OAI21_X1  g235(.A(new_n659), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n653), .A2(new_n657), .A3(new_n654), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT80), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT81), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n676), .A2(new_n674), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n675), .B1(KEYINPUT20), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n672), .A2(new_n676), .A3(new_n674), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n678), .B(new_n679), .C1(KEYINPUT20), .C2(new_n677), .ZN(new_n680));
  XOR2_X1   g255(.A(G1981), .B(G1986), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT82), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G229));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G26), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n481), .A2(G128), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n467), .A2(G140), .ZN(new_n692));
  OR2_X1    g267(.A1(G104), .A2(G2105), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n693), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n690), .B1(new_n696), .B2(new_n689), .ZN(new_n697));
  MUX2_X1   g272(.A(new_n690), .B(new_n697), .S(KEYINPUT28), .Z(new_n698));
  INV_X1    g273(.A(G2067), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G16), .A2(G21), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G168), .B2(G16), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G1966), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n495), .A2(new_n498), .ZN(new_n705));
  INV_X1    g280(.A(new_n493), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n689), .A2(G27), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G2078), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n703), .A2(new_n704), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n710), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n713), .A2(G2078), .B1(new_n702), .B2(G1966), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n700), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n689), .A2(G35), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G162), .B2(new_n689), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT29), .Z(new_n718));
  INV_X1    g293(.A(G2090), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G28), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n721), .A2(KEYINPUT30), .ZN(new_n722));
  AOI21_X1  g297(.A(G29), .B1(new_n721), .B2(KEYINPUT30), .ZN(new_n723));
  OR2_X1    g298(.A1(KEYINPUT31), .A2(G11), .ZN(new_n724));
  NAND2_X1  g299(.A1(KEYINPUT31), .A2(G11), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n722), .A2(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n627), .B2(new_n689), .ZN(new_n727));
  OR2_X1    g302(.A1(G29), .A2(G33), .ZN(new_n728));
  INV_X1    g303(.A(G103), .ZN(new_n729));
  OR3_X1    g304(.A1(new_n469), .A2(KEYINPUT25), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(KEYINPUT25), .B1(new_n469), .B2(new_n729), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n467), .A2(G139), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n496), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n732), .B(new_n733), .C1(new_n466), .C2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n728), .B1(new_n735), .B2(new_n689), .ZN(new_n736));
  INV_X1    g311(.A(G2072), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n727), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n689), .B1(KEYINPUT24), .B2(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(KEYINPUT24), .B2(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n479), .B2(G29), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n736), .A2(new_n737), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n720), .A2(new_n738), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G16), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G5), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G171), .B2(new_n746), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n748), .A2(G1961), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  NOR2_X1   g325(.A1(G29), .A2(G32), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n481), .A2(G129), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n467), .A2(G141), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT26), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n472), .A2(G105), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n752), .A2(new_n753), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  OR3_X1    g332(.A1(new_n757), .A2(KEYINPUT90), .A3(new_n689), .ZN(new_n758));
  OAI21_X1  g333(.A(KEYINPUT90), .B1(new_n757), .B2(new_n689), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n751), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI22_X1  g335(.A1(new_n718), .A2(new_n719), .B1(new_n750), .B2(new_n760), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n715), .A2(new_n745), .A3(new_n749), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n746), .A2(G19), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n547), .B2(new_n746), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G1341), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n746), .A2(G20), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT92), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT23), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n612), .B2(new_n746), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT93), .B(G1956), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n746), .A2(G4), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n615), .B2(new_n746), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(G1348), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(G1348), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n765), .A2(new_n771), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n748), .A2(G1961), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n760), .A2(new_n750), .B1(new_n742), .B2(new_n741), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(KEYINPUT91), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(KEYINPUT91), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n762), .B(new_n777), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G22), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G166), .B2(G16), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT88), .B(G1971), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n746), .A2(G6), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n579), .A2(new_n582), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n746), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT32), .B(G1981), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT85), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n790), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G23), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT86), .ZN(new_n795));
  NAND2_X1  g370(.A1(G288), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n797), .A2(KEYINPUT86), .A3(new_n573), .A4(new_n574), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n794), .B1(new_n799), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT87), .B(KEYINPUT33), .ZN(new_n801));
  INV_X1    g376(.A(G1976), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n800), .A2(new_n803), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n787), .A2(new_n793), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT34), .ZN(new_n807));
  OR2_X1    g382(.A1(G25), .A2(G29), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n481), .A2(G119), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n467), .A2(G131), .ZN(new_n810));
  OR2_X1    g385(.A1(G95), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n808), .B1(new_n813), .B2(new_n689), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT35), .B(G1991), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT83), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT89), .B1(new_n814), .B2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n746), .A2(G24), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n589), .B2(new_n746), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT84), .Z(new_n821));
  AOI211_X1 g396(.A(new_n817), .B(new_n818), .C1(new_n821), .C2(G1986), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n806), .A2(KEYINPUT34), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n821), .A2(G1986), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n807), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n783), .A2(new_n827), .A3(new_n828), .ZN(G311));
  INV_X1    g404(.A(G311), .ZN(G150));
  NAND2_X1  g405(.A1(new_n615), .A2(G559), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT39), .Z(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT96), .B(G55), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n513), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n554), .B2(G93), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n526), .A2(G67), .A3(new_n527), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n837));
  NAND2_X1  g412(.A1(G80), .A2(G543), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G651), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n837), .B1(new_n836), .B2(new_n838), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n835), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n547), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n836), .A2(new_n838), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT95), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n845), .A2(G651), .A3(new_n839), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n846), .A2(new_n546), .A3(new_n835), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(G860), .B1(new_n832), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n832), .B2(new_n850), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT97), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n842), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n856), .ZN(G145));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n488), .A2(new_n858), .A3(new_n492), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n488), .B2(new_n492), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n705), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n695), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n735), .ZN(new_n863));
  INV_X1    g438(.A(new_n757), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n481), .A2(G130), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n467), .A2(G142), .ZN(new_n869));
  OR2_X1    g444(.A1(G106), .A2(G2105), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n870), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n813), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n630), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n867), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n877), .B(new_n630), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n866), .A3(new_n865), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n627), .B(new_n479), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n486), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n880), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT102), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n880), .A2(new_n882), .A3(new_n888), .A4(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n867), .A2(new_n879), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n885), .B1(new_n891), .B2(KEYINPUT101), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n880), .A2(new_n882), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(G37), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g472(.A(new_n848), .B(new_n620), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n615), .A2(G299), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n612), .A2(new_n600), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n615), .A2(G299), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n612), .A2(new_n600), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n904), .A3(KEYINPUT41), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n898), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n900), .A2(new_n901), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n908), .B2(new_n898), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n799), .A2(new_n589), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n799), .A2(new_n589), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(G166), .B(new_n789), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(G305), .B(G166), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n913), .B2(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n911), .A2(new_n912), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n911), .B2(new_n912), .ZN(new_n923));
  OAI21_X1  g498(.A(G868), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n842), .A2(new_n601), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(G295));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n925), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n531), .A2(new_n524), .A3(new_n535), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT70), .B1(new_n538), .B2(new_n534), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n929), .A2(new_n930), .A3(G168), .ZN(new_n931));
  AOI21_X1  g506(.A(G168), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n842), .A2(new_n547), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n546), .B1(new_n846), .B2(new_n835), .ZN(new_n934));
  OAI22_X1  g509(.A1(new_n931), .A2(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(G286), .B1(new_n536), .B2(new_n539), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n929), .A2(new_n930), .A3(G168), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n936), .A2(new_n843), .A3(new_n847), .A4(new_n937), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n902), .A2(new_n905), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n935), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n848), .B(KEYINPUT103), .C1(new_n931), .C2(new_n932), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n939), .B1(new_n943), .B2(new_n908), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n928), .B1(new_n944), .B2(new_n921), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n907), .B1(new_n941), .B2(new_n942), .ZN(new_n946));
  NOR4_X1   g521(.A1(new_n946), .A2(new_n939), .A3(new_n920), .A4(KEYINPUT105), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n945), .A2(new_n947), .A3(G37), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n920), .B(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(new_n939), .B2(new_n946), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT43), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n943), .A2(new_n908), .ZN(new_n953));
  INV_X1    g528(.A(new_n939), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n921), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G37), .B1(new_n955), .B2(KEYINPUT105), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n902), .A2(new_n905), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n941), .A2(new_n957), .A3(new_n942), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n958), .A2(KEYINPUT106), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n908), .A2(new_n938), .A3(new_n935), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n958), .B2(KEYINPUT106), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n950), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n947), .ZN(new_n963));
  AND4_X1   g538(.A1(KEYINPUT43), .A2(new_n956), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT44), .B1(new_n952), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n948), .B2(new_n951), .ZN(new_n968));
  AND4_X1   g543(.A1(new_n967), .A2(new_n956), .A3(new_n962), .A4(new_n963), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n965), .A2(new_n970), .ZN(G397));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT45), .B1(new_n861), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n471), .A2(new_n473), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n496), .A2(G137), .A3(new_n466), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G40), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n973), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n695), .B(new_n699), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT108), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n982), .B2(new_n864), .ZN(new_n983));
  INV_X1    g558(.A(new_n982), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(G1996), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n980), .A2(G1996), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(KEYINPUT107), .A3(new_n864), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n988));
  INV_X1    g563(.A(new_n986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n988), .B1(new_n989), .B2(new_n757), .ZN(new_n990));
  INV_X1    g565(.A(new_n980), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n813), .A2(new_n815), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n813), .A2(new_n815), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n985), .A2(new_n987), .A3(new_n990), .A4(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n589), .B(G1986), .Z(new_n996));
  AOI21_X1  g571(.A(new_n995), .B1(new_n991), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT109), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n999));
  AOI21_X1  g574(.A(G1384), .B1(new_n705), .B2(new_n706), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n979), .B1(new_n1000), .B2(KEYINPUT45), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT110), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n861), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G164), .B2(G1384), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .A4(new_n979), .ZN(new_n1007));
  AOI21_X1  g582(.A(G1971), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n707), .A2(new_n972), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n979), .B1(new_n1009), .B2(KEYINPUT50), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n861), .B2(new_n972), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT111), .B(G2090), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(G8), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G166), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT55), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n861), .A2(new_n1011), .A3(new_n972), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n979), .B1(new_n1000), .B2(new_n1011), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1021), .A2(new_n1022), .A3(new_n1013), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1018), .B(G8), .C1(new_n1008), .C2(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n979), .A2(new_n861), .A3(new_n972), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n802), .B1(new_n796), .B2(new_n798), .ZN(new_n1027));
  OAI211_X1 g602(.A(G8), .B(new_n1026), .C1(new_n1027), .C2(KEYINPUT112), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1029), .B(new_n802), .C1(new_n796), .C2(new_n798), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT52), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n799), .A2(G1976), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1029), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT113), .B(G1976), .Z(new_n1034));
  NAND2_X1  g609(.A1(G288), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT114), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n1038));
  AOI211_X1 g613(.A(new_n1038), .B(KEYINPUT52), .C1(G288), .C2(new_n1034), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n493), .A2(KEYINPUT99), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n488), .A2(new_n858), .A3(new_n492), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1041), .A2(new_n1042), .B1(new_n495), .B2(new_n498), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(G1384), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1016), .B1(new_n1044), .B2(new_n979), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1027), .A2(KEYINPUT112), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1033), .A2(new_n1040), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT49), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT115), .B(G1981), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n789), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n789), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1048), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n789), .A2(new_n1049), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(KEYINPUT49), .C1(new_n1051), .C2(new_n789), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n1045), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1031), .A2(new_n1047), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1031), .A2(new_n1047), .A3(new_n1056), .A4(KEYINPUT118), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1025), .A2(KEYINPUT126), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1020), .A4(new_n1024), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT126), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G299), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n562), .B(KEYINPUT57), .C1(new_n568), .C2(new_n570), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1956), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n474), .A2(G40), .A3(new_n478), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n1009), .B2(new_n1005), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(new_n1003), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1069), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1069), .A2(new_n1071), .A3(new_n1075), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(new_n600), .ZN(new_n1078));
  INV_X1    g653(.A(G1348), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT120), .B1(new_n1026), .B2(G2067), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1044), .A2(new_n1082), .A3(new_n699), .A4(new_n979), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1076), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1080), .A2(KEYINPUT60), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(KEYINPUT124), .A3(new_n600), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT60), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1086), .A2(KEYINPUT124), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n600), .B1(new_n1086), .B2(KEYINPUT124), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT61), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1069), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1069), .A2(new_n1071), .A3(new_n1075), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(KEYINPUT61), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1101));
  XOR2_X1   g676(.A(new_n1101), .B(KEYINPUT123), .Z(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT121), .B(G1996), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1073), .A2(new_n1003), .A3(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1026), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n546), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1103), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1109), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1111), .B(new_n1102), .C1(new_n1112), .C2(new_n546), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1095), .A2(new_n1100), .A3(new_n1110), .A4(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1085), .B1(new_n1093), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1002), .A2(new_n711), .A3(new_n1007), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1072), .B1(new_n1009), .B2(KEYINPUT50), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n861), .A2(new_n1011), .A3(new_n972), .ZN(new_n1121));
  AOI21_X1  g696(.A(G1961), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n478), .A2(G40), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1005), .B1(new_n1043), .B2(G1384), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1118), .A2(G2078), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1127), .A2(new_n1128), .A3(new_n1003), .A4(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1119), .A2(new_n1123), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1116), .B1(new_n1131), .B2(G171), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT127), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n979), .B1(new_n1009), .B2(new_n1005), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1129), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1134), .A2(new_n973), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1119), .A2(G301), .A3(new_n1123), .A4(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1132), .A2(new_n1133), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT51), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n704), .B1(new_n1134), .B2(new_n973), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1120), .A2(new_n742), .A3(new_n1121), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1140), .B(G8), .C1(new_n1143), .C2(G286), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1145));
  AND4_X1   g720(.A1(new_n742), .A2(new_n1121), .A3(new_n979), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1072), .B1(new_n1000), .B2(KEYINPUT45), .ZN(new_n1147));
  AOI21_X1  g722(.A(G1966), .B1(new_n1128), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(G8), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(G286), .A2(G8), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(KEYINPUT51), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1143), .A2(G8), .A3(G286), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1144), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1119), .A2(G301), .A3(new_n1123), .A4(new_n1130), .ZN(new_n1154));
  AOI211_X1 g729(.A(new_n1122), .B(new_n1136), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(G301), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1153), .B1(new_n1156), .B2(new_n1116), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1130), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1122), .B(new_n1158), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1138), .B(KEYINPUT54), .C1(new_n1159), .C2(G301), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT127), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1115), .A2(new_n1139), .A3(new_n1157), .A4(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1144), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1163), .A2(KEYINPUT62), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1155), .A2(G301), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(KEYINPUT62), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1065), .B1(new_n1162), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1143), .A2(G8), .A3(G168), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1169), .B1(new_n1062), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(G8), .B1(new_n1008), .B2(new_n1023), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n1019), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1170), .A2(new_n1169), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1173), .A2(new_n1024), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT119), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT116), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1057), .A2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1031), .A2(new_n1047), .A3(new_n1056), .A4(KEYINPUT116), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1173), .A2(new_n1024), .A3(new_n1174), .ZN(new_n1182));
  OAI21_X1  g757(.A(KEYINPUT119), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1171), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1024), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1178), .A2(new_n1185), .A3(new_n1179), .ZN(new_n1186));
  NOR2_X1   g761(.A1(G288), .A2(G1976), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1056), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1045), .B1(new_n1188), .B2(new_n1050), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(KEYINPUT117), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT117), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1186), .A2(new_n1192), .A3(new_n1189), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1184), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n998), .B1(new_n1168), .B2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n985), .A2(new_n987), .A3(new_n990), .A4(new_n992), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n696), .A2(new_n699), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n980), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AND2_X1   g774(.A1(new_n986), .A2(KEYINPUT46), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n986), .A2(KEYINPUT46), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n983), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT47), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n980), .A2(G1986), .A3(G290), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT48), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n995), .A2(new_n1205), .ZN(new_n1206));
  NOR3_X1   g781(.A1(new_n1199), .A2(new_n1203), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1196), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  AND4_X1   g783(.A1(G319), .A2(new_n687), .A3(new_n650), .A4(new_n667), .ZN(new_n1210));
  OAI211_X1 g784(.A(new_n896), .B(new_n1210), .C1(new_n968), .C2(new_n969), .ZN(G225));
  INV_X1    g785(.A(G225), .ZN(G308));
endmodule


