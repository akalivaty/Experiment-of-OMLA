//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G58), .ZN(new_n208));
  INV_X1    g0008(.A(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G116), .B2(G270), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT65), .B(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n204), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G20), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NAND2_X1  g0027(.A1(new_n202), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n225), .A2(G13), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT64), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT0), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n227), .A2(new_n233), .A3(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G264), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT66), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n231), .A2(new_n256), .A3(KEYINPUT68), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G20), .B2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G159), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n208), .A2(new_n221), .ZN(new_n262));
  OAI21_X1  g0062(.A(G20), .B1(new_n262), .B2(new_n201), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n256), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(new_n231), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT7), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n270), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT75), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT75), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n269), .A2(new_n274), .A3(new_n270), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n271), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(KEYINPUT16), .B(new_n265), .C1(new_n276), .C2(new_n221), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n230), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT16), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n281), .A2(new_n282), .A3(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT7), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n221), .B1(new_n284), .B2(new_n272), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n280), .B1(new_n285), .B2(new_n264), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n277), .A2(new_n279), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G13), .A3(G20), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n279), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n291), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT69), .ZN(new_n296));
  INV_X1    g0096(.A(new_n291), .ZN(new_n297));
  OR3_X1    g0097(.A1(new_n297), .A2(new_n279), .A3(KEYINPUT69), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n290), .A2(G20), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n293), .B1(new_n300), .B2(new_n288), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n287), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G41), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G1), .A3(G13), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n290), .B1(G41), .B2(G45), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n305), .A2(G232), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT76), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n215), .A2(G1698), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n309), .B1(G223), .B2(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G87), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G274), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n306), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n308), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G169), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n318), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n303), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n322), .B(KEYINPUT18), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G190), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n308), .A2(new_n314), .A3(new_n326), .A4(new_n317), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n287), .A2(new_n328), .A3(new_n302), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT17), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n257), .A2(new_n259), .ZN(new_n335));
  INV_X1    g0135(.A(G150), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n231), .A2(G33), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n335), .A2(new_n336), .B1(new_n337), .B2(new_n288), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n231), .B1(new_n201), .B2(new_n214), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n279), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n297), .A2(new_n214), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n340), .B(new_n341), .C1(new_n214), .C2(new_n300), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT9), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(KEYINPUT67), .A2(G223), .ZN(new_n345));
  NOR2_X1   g0145(.A1(KEYINPUT67), .A2(G223), .ZN(new_n346));
  OAI21_X1  g0146(.A(G1698), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT3), .B(G33), .ZN(new_n348));
  INV_X1    g0148(.A(G1698), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G222), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n351), .B(new_n313), .C1(G77), .C2(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n305), .A2(new_n306), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n352), .B(new_n317), .C1(new_n215), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G200), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n342), .A2(new_n343), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n354), .A2(new_n326), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n344), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(KEYINPUT10), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(KEYINPUT10), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(new_n354), .A2(G179), .ZN(new_n362));
  INV_X1    g0162(.A(G169), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n354), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n342), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n289), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n337), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT70), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n291), .B(new_n370), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n371), .A2(new_n299), .A3(new_n294), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n279), .A2(new_n369), .B1(new_n372), .B2(G77), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n291), .B(KEYINPUT70), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n216), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n349), .A2(G232), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n348), .B(new_n378), .C1(new_n222), .C2(new_n349), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n379), .B(new_n313), .C1(G107), .C2(new_n348), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(new_n317), .C1(new_n217), .C2(new_n353), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(new_n326), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(G200), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n377), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n366), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n333), .A2(new_n334), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT13), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n209), .A2(G1698), .ZN(new_n389));
  OAI221_X1 g0189(.A(new_n389), .B1(G226), .B2(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G97), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n316), .B1(new_n392), .B2(new_n313), .ZN(new_n393));
  INV_X1    g0193(.A(G238), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n353), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n388), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n305), .B1(new_n390), .B2(new_n391), .ZN(new_n398));
  NOR4_X1   g0198(.A1(new_n398), .A2(KEYINPUT13), .A3(new_n395), .A4(new_n316), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT72), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n392), .A2(new_n313), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(new_n396), .A3(new_n317), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(new_n400), .A3(KEYINPUT13), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(G190), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n231), .A2(G68), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n337), .A2(new_n216), .ZN(new_n408));
  AOI211_X1 g0208(.A(new_n407), .B(new_n408), .C1(G50), .C2(new_n260), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT11), .B1(new_n409), .B2(new_n294), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT11), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n335), .A2(new_n214), .B1(new_n231), .B2(G68), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(new_n279), .C1(new_n412), .C2(new_n408), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n297), .A2(KEYINPUT12), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT12), .ZN(new_n417));
  OAI21_X1  g0217(.A(G68), .B1(new_n372), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n374), .A2(KEYINPUT12), .A3(new_n221), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n414), .A2(new_n416), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n406), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(G200), .B1(new_n397), .B2(new_n399), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT71), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(KEYINPUT71), .B(G200), .C1(new_n397), .C2(new_n399), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT73), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n403), .A2(KEYINPUT13), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n393), .A2(new_n388), .A3(new_n396), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(KEYINPUT72), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n404), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n420), .B1(new_n432), .B2(G190), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT73), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n425), .A2(new_n426), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n428), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n320), .B1(new_n431), .B2(new_n404), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT74), .B(KEYINPUT14), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n429), .A2(new_n430), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n440), .B1(new_n441), .B2(G169), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT74), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT14), .ZN(new_n445));
  OAI211_X1 g0245(.A(G169), .B(new_n445), .C1(new_n397), .C2(new_n399), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n439), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n420), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n381), .A2(G179), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n381), .A2(new_n363), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n376), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n437), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n387), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT85), .ZN(new_n454));
  AND2_X1   g0254(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n455));
  NOR2_X1   g0255(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n455), .A2(new_n456), .A3(new_n391), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n457), .B2(G20), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n210), .A2(new_n204), .A3(new_n205), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n460));
  OAI211_X1 g0260(.A(KEYINPUT85), .B(new_n231), .C1(new_n460), .C2(new_n391), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n348), .A2(new_n231), .A3(G68), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n460), .B1(new_n204), .B2(new_n337), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n465), .A2(new_n279), .B1(new_n374), .B2(new_n368), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n313), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n469), .A2(G250), .B1(G274), .B2(new_n468), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n394), .A2(new_n349), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n217), .A2(G1698), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n472), .C1(new_n281), .C2(new_n282), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G116), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n313), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n470), .A2(new_n476), .A3(G190), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n294), .B(new_n291), .C1(G1), .C2(new_n256), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G87), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n466), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n470), .A2(new_n476), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G200), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(G179), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n478), .A2(new_n368), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT86), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n466), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n482), .A2(new_n363), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n481), .A2(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g0289(.A(G97), .B(G107), .ZN(new_n490));
  NOR2_X1   g0290(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n491), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n204), .A2(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G97), .A2(G107), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n493), .A2(new_n206), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G20), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT79), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n260), .A2(G77), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n284), .A2(new_n272), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G107), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n231), .B1(new_n492), .B2(new_n496), .ZN(new_n504));
  INV_X1    g0304(.A(new_n500), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT79), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(new_n279), .B1(new_n204), .B2(new_n297), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n479), .A2(G97), .ZN(new_n509));
  OAI211_X1 g0309(.A(G244), .B(new_n349), .C1(new_n281), .C2(new_n282), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT80), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(G250), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT81), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n348), .A2(G244), .A3(new_n349), .A4(new_n512), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n514), .A2(new_n517), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n515), .A2(new_n516), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n313), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g0322(.A(KEYINPUT5), .B(G41), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(G274), .A3(new_n468), .ZN(new_n524));
  AND2_X1   g0324(.A1(KEYINPUT5), .A2(G41), .ZN(new_n525));
  NOR2_X1   g0325(.A1(KEYINPUT5), .A2(G41), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n468), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(G257), .A3(new_n305), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT82), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT82), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n527), .A2(new_n530), .A3(G257), .A4(new_n305), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n522), .A2(new_n524), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n508), .A2(new_n509), .B1(new_n363), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT83), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n534), .B2(G179), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n516), .A2(new_n515), .B1(new_n510), .B2(new_n513), .ZN(new_n538));
  INV_X1    g0338(.A(new_n521), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n538), .A2(new_n539), .A3(new_n518), .A4(new_n519), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n532), .B1(new_n540), .B2(new_n313), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n541), .A2(KEYINPUT83), .A3(new_n320), .A4(new_n524), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n535), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n534), .A2(G200), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n541), .A2(G190), .A3(new_n524), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n508), .A2(new_n545), .A3(new_n546), .A4(new_n509), .ZN(new_n547));
  INV_X1    g0347(.A(G116), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n290), .B2(G33), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n371), .A2(new_n294), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n374), .A2(new_n548), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n278), .A2(new_n230), .B1(G20), .B2(new_n548), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n519), .B(new_n231), .C1(G33), .C2(new_n204), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n552), .A2(KEYINPUT20), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT20), .B1(new_n552), .B2(new_n553), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n550), .B(new_n551), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G264), .A2(G1698), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n348), .B(new_n557), .C1(new_n223), .C2(G1698), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n281), .A2(new_n282), .ZN(new_n559));
  INV_X1    g0359(.A(G303), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(new_n313), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n527), .A2(G270), .A3(new_n305), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT87), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT87), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n527), .A2(new_n565), .A3(G270), .A4(new_n305), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n562), .A2(new_n564), .A3(new_n524), .A4(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n556), .A2(new_n567), .A3(G169), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n567), .A2(new_n320), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n556), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n556), .A2(new_n567), .A3(KEYINPUT21), .A4(G169), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n567), .A2(G200), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n326), .B2(new_n567), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(new_n556), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n489), .A2(new_n544), .A3(new_n547), .A4(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n527), .A2(G264), .A3(new_n305), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n211), .A2(new_n349), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n223), .A2(G1698), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n281), .C2(new_n282), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G33), .A2(G294), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n305), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n524), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n581), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT90), .B1(new_n588), .B2(new_n363), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n584), .A2(new_n585), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n580), .B(new_n524), .C1(new_n590), .C2(new_n305), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT90), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(G169), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT91), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n591), .B2(new_n320), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n581), .A2(new_n586), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n597), .A2(KEYINPUT91), .A3(G179), .A4(new_n524), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT89), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n231), .B(G87), .C1(new_n281), .C2(new_n282), .ZN(new_n602));
  NOR2_X1   g0402(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n348), .A2(new_n231), .A3(G87), .A4(new_n603), .ZN(new_n606));
  NAND2_X1  g0406(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n231), .A2(G107), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT23), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT24), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT24), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n608), .A2(new_n614), .A3(new_n609), .A4(new_n611), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n279), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n478), .A2(new_n205), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n610), .A2(new_n290), .A3(G13), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n619), .B(KEYINPUT25), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n601), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n294), .B1(new_n613), .B2(new_n615), .ZN(new_n623));
  INV_X1    g0423(.A(new_n621), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n623), .A2(KEYINPUT89), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n600), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT92), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n588), .A2(G190), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n591), .A2(G200), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n617), .A2(new_n621), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n626), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n617), .A2(new_n601), .A3(new_n621), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT89), .B1(new_n623), .B2(new_n624), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n632), .A2(new_n633), .B1(new_n594), .B2(new_n599), .ZN(new_n634));
  INV_X1    g0434(.A(new_n630), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT92), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n579), .B1(new_n631), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n453), .A2(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n451), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n437), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n331), .B1(new_n640), .B2(new_n448), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(new_n323), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n361), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n365), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n387), .A2(new_n452), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n489), .A2(KEYINPUT26), .A3(new_n535), .A4(new_n543), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT93), .B1(new_n475), .B2(new_n313), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT93), .ZN(new_n649));
  AOI211_X1 g0449(.A(new_n649), .B(new_n305), .C1(new_n473), .C2(new_n474), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n470), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G200), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n481), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n617), .A2(new_n621), .B1(new_n594), .B2(new_n599), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n630), .B(new_n547), .C1(new_n655), .C2(new_n574), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n656), .B2(new_n544), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n647), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n651), .A2(new_n363), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n487), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n645), .B1(new_n646), .B2(new_n662), .ZN(G369));
  INV_X1    g0463(.A(G13), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G20), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n290), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n556), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n578), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n574), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n672), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  INV_X1    g0476(.A(new_n671), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n632), .B2(new_n633), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n636), .B2(new_n631), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n626), .A2(new_n677), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n636), .A2(new_n631), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n674), .A2(new_n671), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n682), .A2(new_n683), .B1(new_n655), .B2(new_n677), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n234), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n459), .A2(G116), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G1), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n228), .B2(new_n688), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n660), .B(new_n653), .C1(new_n634), .C2(new_n574), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n544), .A2(new_n630), .A3(new_n547), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT98), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n653), .A2(new_n660), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n626), .B2(new_n674), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT98), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n544), .A2(new_n630), .A3(new_n547), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n660), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT26), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n487), .A2(new_n488), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n466), .A2(new_n483), .A3(new_n477), .A4(new_n480), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n706), .B2(new_n544), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n653), .A2(KEYINPUT26), .A3(new_n535), .A4(new_n543), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n702), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n696), .A2(new_n701), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n693), .B1(new_n710), .B2(new_n677), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n661), .A2(new_n677), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT97), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n671), .B1(new_n658), .B2(new_n660), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT97), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n711), .B1(new_n717), .B2(new_n693), .ZN(new_n718));
  AND4_X1   g0518(.A1(new_n489), .A2(new_n544), .A3(new_n547), .A4(new_n578), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n634), .A2(new_n635), .A3(KEYINPUT92), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n627), .B1(new_n626), .B2(new_n630), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n719), .B(new_n677), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n651), .A2(new_n320), .A3(new_n567), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n591), .A3(new_n534), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT95), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n723), .A2(new_n726), .A3(new_n591), .A4(new_n534), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n567), .A2(new_n320), .A3(new_n482), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT94), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n728), .A2(new_n597), .A3(new_n541), .A4(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n597), .A3(new_n541), .ZN(new_n732));
  INV_X1    g0532(.A(new_n730), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n725), .A2(new_n727), .A3(new_n731), .A4(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(new_n671), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n734), .A2(new_n731), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n677), .B1(new_n738), .B2(new_n724), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n739), .B2(new_n736), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n722), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT96), .B1(new_n741), .B2(G330), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT96), .ZN(new_n743));
  INV_X1    g0543(.A(G330), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n743), .B(new_n744), .C1(new_n722), .C2(new_n740), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n718), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n692), .B1(new_n747), .B2(G1), .ZN(G364));
  NAND2_X1  g0548(.A1(new_n665), .A2(G45), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n688), .A2(G1), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n676), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G330), .B2(new_n675), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n231), .A2(new_n326), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n324), .A2(G179), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n231), .A2(G190), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n320), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G87), .A2(new_n757), .B1(new_n761), .B2(G77), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n754), .A2(new_n759), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n208), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n758), .A2(new_n755), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT99), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n764), .B1(G107), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n758), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n770), .A2(KEYINPUT32), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(KEYINPUT32), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n320), .A2(new_n324), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n754), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n772), .B(new_n773), .C1(new_n214), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n231), .B1(new_n769), .B2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n204), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n776), .A2(new_n559), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n774), .A2(new_n758), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n768), .B(new_n779), .C1(new_n221), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n780), .ZN(new_n782));
  INV_X1    g0582(.A(G317), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT33), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(KEYINPUT33), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n770), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G329), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n786), .B(new_n788), .C1(new_n560), .C2(new_n756), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n348), .B(new_n789), .C1(G311), .C2(new_n761), .ZN(new_n790));
  INV_X1    g0590(.A(new_n775), .ZN(new_n791));
  INV_X1    g0591(.A(new_n777), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n791), .A2(G326), .B1(new_n792), .B2(G294), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT100), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n790), .B(new_n794), .C1(new_n795), .C2(new_n766), .ZN(new_n796));
  INV_X1    g0596(.A(G322), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n763), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n781), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n230), .B1(G20), .B2(new_n363), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n800), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n686), .A2(new_n348), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n229), .A2(new_n467), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n805), .B(new_n806), .C1(new_n251), .C2(new_n467), .ZN(new_n807));
  INV_X1    g0607(.A(G355), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n348), .A2(new_n234), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(G116), .B2(new_n234), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n799), .A2(new_n800), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n803), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n811), .B(new_n751), .C1(new_n675), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n753), .A2(new_n813), .ZN(G396));
  OR2_X1    g0614(.A1(new_n451), .A2(KEYINPUT102), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n451), .A2(KEYINPUT102), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n385), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n671), .B(new_n818), .C1(new_n658), .C2(new_n660), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n376), .A2(new_n671), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n817), .A2(new_n821), .B1(new_n639), .B2(new_n671), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n820), .B1(new_n717), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(new_n746), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n746), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n750), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G294), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n763), .A2(new_n828), .B1(new_n770), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n767), .B2(G87), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n757), .A2(G107), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n559), .B1(new_n780), .B2(new_n795), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n778), .B(new_n833), .C1(G116), .C2(new_n761), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n791), .A2(G303), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n831), .A2(new_n832), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n763), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G143), .A2(new_n837), .B1(new_n782), .B2(G150), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n839), .B2(new_n775), .C1(new_n771), .C2(new_n760), .ZN(new_n840));
  XNOR2_X1  g0640(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n840), .B(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n348), .B1(new_n756), .B2(new_n214), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G58), .B2(new_n792), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n844), .B1(new_n845), .B2(new_n770), .C1(new_n221), .C2(new_n766), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n836), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n800), .A2(new_n801), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n847), .A2(new_n800), .B1(new_n216), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n751), .B(new_n849), .C1(new_n823), .C2(new_n802), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n827), .A2(new_n850), .ZN(G384));
  INV_X1    g0651(.A(KEYINPUT104), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n269), .A2(new_n274), .A3(new_n270), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n274), .B1(new_n269), .B2(new_n270), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n284), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n264), .B1(new_n855), .B2(G68), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n294), .B1(new_n856), .B2(KEYINPUT16), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n265), .B1(new_n276), .B2(new_n221), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n280), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n301), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n321), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n852), .B(new_n329), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n277), .A2(new_n279), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n856), .A2(KEYINPUT16), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n302), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n669), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n865), .A2(new_n321), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n852), .B1(new_n869), .B2(new_n329), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT105), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n303), .A2(new_n866), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n322), .A2(new_n873), .A3(new_n329), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT105), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n877), .B(KEYINPUT37), .C1(new_n868), .C2(new_n870), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n872), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n332), .A2(new_n867), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n332), .A2(new_n873), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n874), .B(KEYINPUT37), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n447), .A2(KEYINPUT103), .A3(new_n420), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT103), .ZN(new_n888));
  INV_X1    g0688(.A(new_n446), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n438), .A2(new_n442), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n888), .B1(new_n890), .B2(new_n421), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n421), .A2(new_n677), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n428), .B2(new_n436), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  AND4_X1   g0695(.A1(new_n434), .A2(new_n435), .A3(new_n406), .A4(new_n421), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n434), .B1(new_n433), .B2(new_n435), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n890), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n893), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n822), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n735), .B(new_n671), .C1(KEYINPUT106), .C2(KEYINPUT31), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n735), .A2(new_n671), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT106), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n903), .A3(new_n736), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n722), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n886), .A2(KEYINPUT40), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n900), .A2(new_n905), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n879), .A2(new_n880), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n882), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n908), .B1(new_n910), .B2(new_n881), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n907), .B1(new_n911), .B2(KEYINPUT40), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n453), .A2(new_n905), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n912), .B(new_n913), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(G330), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n715), .B1(new_n661), .B2(new_n677), .ZN(new_n916));
  AOI211_X1 g0716(.A(KEYINPUT97), .B(new_n671), .C1(new_n658), .C2(new_n660), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n693), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n711), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n646), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n920), .A2(new_n644), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n915), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n815), .A2(new_n816), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n923), .A2(new_n671), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n714), .B2(new_n817), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n895), .A2(new_n899), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n910), .A2(new_n881), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n928), .A2(new_n929), .B1(new_n323), .B2(new_n669), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n886), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n910), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n892), .A2(new_n671), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n922), .B(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n290), .B2(new_n665), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n548), .B1(new_n497), .B2(KEYINPUT35), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n939), .B(new_n232), .C1(KEYINPUT35), .C2(new_n497), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT36), .ZN(new_n941));
  OAI21_X1  g0741(.A(G77), .B1(new_n208), .B2(new_n221), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n228), .A2(new_n942), .B1(G50), .B2(new_n221), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(G1), .A3(new_n664), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n938), .A2(new_n941), .A3(new_n944), .ZN(G367));
  AOI22_X1  g0745(.A1(G58), .A2(new_n757), .B1(new_n782), .B2(G159), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n839), .B2(new_n770), .C1(new_n336), .C2(new_n763), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n777), .A2(new_n221), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n348), .B1(new_n765), .B2(new_n216), .C1(new_n214), .C2(new_n760), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(G143), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n775), .ZN(new_n952));
  INV_X1    g0752(.A(new_n765), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n791), .A2(G311), .B1(new_n953), .B2(G97), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n795), .B2(new_n760), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n757), .A2(KEYINPUT46), .A3(G116), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT46), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n756), .B2(new_n548), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n956), .B(new_n958), .C1(new_n205), .C2(new_n777), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n559), .B1(new_n770), .B2(new_n783), .C1(new_n560), .C2(new_n763), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n955), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n828), .B2(new_n780), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n952), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT115), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT47), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n750), .B1(new_n965), .B2(new_n800), .ZN(new_n966));
  INV_X1    g0766(.A(new_n805), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n804), .B1(new_n234), .B2(new_n368), .C1(new_n247), .C2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n466), .A2(new_n480), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n671), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n653), .A2(new_n660), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n660), .B2(new_n970), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n966), .B(new_n968), .C1(new_n812), .C2(new_n972), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT109), .Z(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT107), .B1(new_n544), .B2(new_n677), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT107), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n535), .A2(new_n543), .A3(new_n978), .A4(new_n671), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n508), .A2(new_n509), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n544), .B(new_n547), .C1(new_n981), .C2(new_n677), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n682), .A2(new_n683), .ZN(new_n985));
  OAI21_X1  g0785(.A(KEYINPUT42), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n983), .A2(new_n634), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n671), .B1(new_n988), .B2(new_n544), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT108), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n989), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT108), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(new_n992), .A3(new_n986), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n983), .A2(new_n682), .A3(new_n683), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n990), .B(new_n993), .C1(KEYINPUT42), .C2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n976), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n681), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n996), .A3(new_n976), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n998), .A2(new_n999), .A3(new_n983), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1000), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n1002), .A2(new_n997), .B1(new_n681), .B2(new_n984), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n749), .A2(G1), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT114), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n684), .A2(new_n983), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT44), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n684), .A2(new_n983), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(KEYINPUT111), .B(KEYINPUT112), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT45), .Z(new_n1011));
  XNOR2_X1  g0811(.A(new_n1009), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n999), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1008), .A2(new_n681), .A3(new_n1012), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n679), .A2(new_n680), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n674), .B2(new_n671), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n985), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT113), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n1020), .A3(new_n676), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n676), .A2(new_n1020), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n676), .A2(new_n1020), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1018), .A2(new_n985), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n718), .A2(new_n1025), .A3(new_n746), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n747), .B1(new_n1016), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(KEYINPUT110), .B(KEYINPUT41), .Z(new_n1028));
  XNOR2_X1  g0828(.A(new_n687), .B(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1006), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n973), .B1(new_n1004), .B2(new_n1031), .ZN(G387));
  NAND2_X1  g0832(.A1(new_n1026), .A2(new_n687), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT118), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT118), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n747), .C2(new_n1025), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1025), .A2(new_n1006), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G311), .A2(new_n782), .B1(new_n837), .B2(G317), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n560), .B2(new_n760), .C1(new_n797), .C2(new_n775), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT117), .Z(new_n1040));
  AOI22_X1  g0840(.A1(new_n1040), .A2(KEYINPUT48), .B1(G283), .B2(new_n792), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(KEYINPUT48), .B2(new_n1040), .C1(new_n828), .C2(new_n756), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT49), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n787), .A2(G326), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n348), .B1(new_n953), .B2(G116), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n214), .A2(new_n763), .B1(new_n780), .B2(new_n288), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n767), .B2(G97), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n348), .B1(new_n770), .B2(new_n336), .C1(new_n221), .C2(new_n760), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n777), .A2(new_n368), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n756), .A2(new_n216), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1050), .B(new_n1054), .C1(new_n771), .C2(new_n775), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1048), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n288), .A2(G50), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT50), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n221), .A2(new_n216), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n689), .ZN(new_n1060));
  AOI211_X1 g0860(.A(G45), .B(new_n1059), .C1(new_n1060), .C2(KEYINPUT116), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1058), .B(new_n1061), .C1(KEYINPUT116), .C2(new_n1060), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n805), .C1(new_n243), .C2(new_n467), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(G107), .B2(new_n234), .C1(new_n689), .C2(new_n809), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1056), .A2(new_n800), .B1(new_n804), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1017), .A2(new_n803), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n751), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1036), .A2(new_n1037), .A3(new_n1067), .ZN(G393));
  AOI21_X1  g0868(.A(new_n688), .B1(new_n1016), .B2(new_n1026), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1016), .B2(new_n1026), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT119), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1016), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1014), .A2(KEYINPUT119), .A3(new_n1015), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1072), .A2(new_n1006), .A3(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n804), .B1(new_n204), .B2(new_n234), .C1(new_n254), .C2(new_n967), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G68), .A2(new_n757), .B1(new_n761), .B2(new_n289), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n214), .B2(new_n780), .C1(new_n951), .C2(new_n770), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n777), .A2(new_n216), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1077), .A2(new_n559), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n210), .B2(new_n766), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n775), .A2(new_n336), .B1(new_n763), .B2(new_n771), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT51), .Z(new_n1082));
  NOR2_X1   g0882(.A1(new_n756), .A2(new_n795), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n559), .B1(new_n777), .B2(new_n548), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n780), .A2(new_n560), .B1(new_n760), .B2(new_n828), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(G322), .C2(new_n787), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n775), .A2(new_n783), .B1(new_n763), .B2(new_n829), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT52), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(new_n205), .C2(new_n766), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1080), .A2(new_n1082), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n750), .B1(new_n1090), .B2(new_n800), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1075), .B(new_n1091), .C1(new_n983), .C2(new_n812), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1070), .A2(new_n1074), .A3(new_n1092), .ZN(G390));
  NAND2_X1  g0893(.A1(new_n932), .A2(new_n933), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n801), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n559), .B1(new_n780), .B2(new_n205), .C1(new_n210), .C2(new_n756), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1078), .B(new_n1096), .C1(G294), .C2(new_n787), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n791), .A2(G283), .B1(new_n761), .B2(G97), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n221), .C2(new_n766), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G116), .B2(new_n837), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n765), .A2(new_n214), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT54), .B(G143), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n348), .B1(new_n760), .B2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(G159), .C2(new_n792), .ZN(new_n1104));
  INV_X1    g0904(.A(G125), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n770), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n756), .A2(new_n336), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT53), .ZN(new_n1108));
  INV_X1    g0908(.A(G128), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n775), .C1(new_n845), .C2(new_n763), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1106), .B(new_n1110), .C1(G137), .C2(new_n782), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n800), .B1(new_n1100), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n848), .A2(new_n288), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1095), .A2(new_n751), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n934), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n926), .B1(new_n819), .B2(new_n924), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n932), .A2(new_n933), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n886), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n710), .A2(new_n677), .A3(new_n817), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n924), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n927), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1118), .A2(new_n1121), .A3(new_n934), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n823), .B(new_n926), .C1(new_n742), .C2(new_n745), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1117), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n905), .A2(G330), .A3(new_n823), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1125), .A2(new_n927), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1115), .B1(new_n925), .B2(new_n927), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n880), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT38), .B1(new_n879), .B2(new_n880), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1128), .A2(new_n1129), .A3(new_n931), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT39), .B1(new_n881), .B2(new_n885), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1127), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1115), .B(new_n886), .C1(new_n1133), .C2(new_n927), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1126), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1006), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1114), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n453), .A2(G330), .A3(new_n905), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n920), .A2(new_n1139), .A3(new_n644), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1125), .A2(new_n927), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1123), .A2(new_n1133), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n823), .B1(new_n742), .B2(new_n745), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1126), .B1(new_n1143), .B2(new_n927), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1142), .B1(new_n1144), .B2(new_n925), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1140), .B(new_n1145), .C1(new_n1124), .C2(new_n1135), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1146), .A2(new_n687), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1136), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1138), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(G378));
  OAI211_X1 g0951(.A(G330), .B(new_n907), .C1(new_n911), .C2(KEYINPUT40), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n936), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n935), .A3(new_n930), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n366), .B(KEYINPUT55), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n342), .A2(new_n866), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT56), .Z(new_n1158));
  XNOR2_X1  g0958(.A(new_n1156), .B(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1154), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1159), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1155), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1152), .B1(new_n935), .B2(new_n930), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1160), .A2(new_n1164), .B1(new_n1146), .B2(new_n1140), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n688), .B1(new_n1165), .B2(KEYINPUT57), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1160), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1146), .A2(new_n1140), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1166), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1159), .A2(new_n801), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n848), .A2(new_n214), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n763), .A2(new_n1109), .B1(new_n777), .B2(new_n336), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n761), .A2(G137), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n845), .B2(new_n780), .C1(new_n756), .C2(new_n1102), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(G125), .C2(new_n791), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT59), .ZN(new_n1179));
  AOI21_X1  g0979(.A(G41), .B1(new_n787), .B2(G124), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G33), .B1(new_n953), .B2(G159), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n214), .B1(new_n281), .B2(G41), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G116), .A2(new_n791), .B1(new_n782), .B2(G97), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n208), .B2(new_n765), .C1(new_n795), .C2(new_n770), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n763), .A2(new_n205), .B1(new_n760), .B2(new_n368), .ZN(new_n1186));
  OR4_X1    g0986(.A1(G41), .A2(new_n1186), .A3(new_n948), .A4(new_n1053), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1185), .A2(new_n1187), .A3(new_n348), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT58), .Z(new_n1189));
  NAND3_X1  g0989(.A1(new_n1182), .A2(new_n1183), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n750), .B1(new_n1190), .B2(new_n800), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1173), .A2(new_n1174), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1167), .B2(new_n1006), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1172), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT120), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1167), .A2(new_n1006), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1192), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1166), .B2(new_n1171), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT120), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1196), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(G375));
  NAND3_X1  g1003(.A1(new_n453), .A2(G330), .A3(new_n905), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n645), .B(new_n1204), .C1(new_n718), .C2(new_n646), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1125), .A2(new_n927), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n738), .A2(new_n724), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n671), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT31), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n637), .A2(new_n677), .B1(new_n1209), .B2(new_n737), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n743), .B1(new_n1210), .B2(new_n744), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n741), .A2(KEYINPUT96), .A3(G330), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n822), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1206), .B1(new_n1213), .B2(new_n926), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n925), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1205), .A2(new_n1216), .A3(new_n1142), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1148), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(new_n1029), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT121), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1145), .A2(new_n1006), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n775), .A2(new_n845), .B1(new_n770), .B2(new_n1109), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n348), .B1(new_n765), .B2(new_n208), .C1(new_n839), .C2(new_n763), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(G159), .C2(new_n757), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n760), .A2(new_n336), .B1(new_n777), .B2(new_n214), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT123), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(new_n780), .C2(new_n1102), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n559), .B1(new_n795), .B2(new_n763), .C1(new_n766), .C2(new_n216), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n756), .A2(new_n204), .B1(new_n770), .B2(new_n560), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT122), .Z(new_n1230));
  OAI22_X1  g1030(.A1(new_n775), .A2(new_n828), .B1(new_n760), .B2(new_n205), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1052), .B(new_n1231), .C1(G116), .C2(new_n782), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1227), .B1(new_n1228), .B2(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1234), .A2(new_n800), .B1(new_n221), .B2(new_n848), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n751), .B(new_n1235), .C1(new_n926), .C2(new_n802), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1221), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1220), .A2(new_n1238), .ZN(G381));
  OR2_X1    g1039(.A1(G387), .A2(G390), .ZN(new_n1240));
  INV_X1    g1040(.A(G396), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1036), .A2(new_n1241), .A3(new_n1037), .A4(new_n1067), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G381), .A2(G384), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1202), .A2(new_n1150), .A3(new_n1243), .A4(new_n1244), .ZN(G407));
  NAND3_X1  g1045(.A1(new_n1196), .A2(new_n1150), .A3(new_n1201), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n670), .A2(G213), .ZN(new_n1247));
  OR3_X1    g1047(.A1(new_n1246), .A2(KEYINPUT124), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT124), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1248), .A2(G213), .A3(G407), .A4(new_n1249), .ZN(G409));
  NAND3_X1  g1050(.A1(new_n1167), .A2(new_n1168), .A3(new_n1030), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT125), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT125), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1167), .A2(new_n1168), .A3(new_n1253), .A4(new_n1030), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1252), .A2(new_n1150), .A3(new_n1194), .A4(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1247), .B(new_n1255), .C1(new_n1199), .C2(new_n1150), .ZN(new_n1256));
  INV_X1    g1056(.A(G384), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT60), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1217), .B2(new_n1148), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1145), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT60), .B1(new_n1260), .B2(new_n1205), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1259), .A2(new_n688), .A3(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1257), .B1(new_n1262), .B2(new_n1237), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1218), .A2(KEYINPUT60), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1261), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n687), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(G384), .A3(new_n1238), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT62), .B1(new_n1256), .B2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n670), .A2(G213), .A3(G2897), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1263), .A2(new_n1267), .A3(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1263), .B2(new_n1267), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT61), .B1(new_n1256), .B2(new_n1273), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1255), .A2(new_n1247), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1195), .A2(G378), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1268), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1269), .A2(new_n1274), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G393), .A2(G396), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1281), .A2(new_n1242), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(G387), .A2(G390), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1240), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1242), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(new_n1240), .A3(new_n1283), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1256), .B2(new_n1268), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1256), .A2(KEYINPUT126), .A3(new_n1273), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT126), .B1(new_n1256), .B2(new_n1273), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1291), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1275), .A2(new_n1276), .A3(KEYINPUT63), .A4(new_n1278), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(new_n1289), .A3(new_n1296), .ZN(new_n1297));
  OAI22_X1  g1097(.A1(new_n1280), .A2(new_n1289), .B1(new_n1294), .B2(new_n1297), .ZN(G405));
  NAND2_X1  g1098(.A1(new_n1278), .A2(KEYINPUT127), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1288), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1285), .A2(new_n1299), .A3(new_n1287), .ZN(new_n1302));
  AND4_X1   g1102(.A1(new_n1246), .A2(new_n1301), .A3(new_n1276), .A4(new_n1302), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n1301), .A2(new_n1302), .B1(new_n1246), .B2(new_n1276), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(G402));
endmodule


