//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n202), .B1(new_n210), .B2(KEYINPUT66), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n211), .B1(KEYINPUT66), .B2(new_n210), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT67), .Z(new_n213));
  AND2_X1   g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n213), .A2(G20), .A3(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G1), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n222));
  XNOR2_X1  g0022(.A(new_n221), .B(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n224), .B1(new_n203), .B2(new_n225), .C1(new_n207), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n219), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n215), .B(new_n223), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT68), .Z(new_n234));
  NOR2_X1   g0034(.A1(new_n232), .A2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT69), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT2), .B(G226), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n239), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT79), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n253), .A2(KEYINPUT79), .A3(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n217), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT7), .ZN(new_n261));
  XOR2_X1   g0061(.A(KEYINPUT80), .B(KEYINPUT7), .Z(new_n262));
  NAND4_X1  g0062(.A1(new_n262), .A2(new_n258), .A3(new_n217), .A4(new_n259), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(G68), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G58), .ZN(new_n265));
  INV_X1    g0065(.A(G68), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(G20), .B1(new_n267), .B2(new_n201), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G159), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n264), .A2(KEYINPUT16), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT16), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n262), .B1(G20), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n254), .A2(new_n256), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n266), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n274), .B1(new_n279), .B2(new_n271), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G1), .A2(G13), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n273), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT72), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(new_n217), .B2(G1), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n216), .A2(KEYINPUT72), .A3(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n216), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n283), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n291), .A2(new_n294), .B1(new_n293), .B2(new_n290), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n284), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT70), .B1(new_n297), .B2(new_n282), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT70), .ZN(new_n299));
  NAND2_X1  g0099(.A1(G33), .A2(G41), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n214), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n216), .B1(G41), .B2(G45), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n298), .A2(new_n301), .A3(new_n303), .A4(G274), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n298), .A2(new_n301), .A3(G232), .A4(new_n302), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT71), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n297), .A2(new_n307), .A3(new_n282), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT71), .B1(new_n214), .B2(new_n300), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OR2_X1    g0110(.A1(G223), .A2(G1698), .ZN(new_n311));
  INV_X1    g0111(.A(G226), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G1698), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n258), .B2(new_n259), .ZN(new_n315));
  INV_X1    g0115(.A(G87), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n255), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n310), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n306), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G169), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n306), .A2(new_n318), .A3(G179), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n296), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT18), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n284), .A2(new_n295), .B1(new_n321), .B2(new_n320), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT18), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n306), .A2(new_n318), .A3(G190), .ZN(new_n328));
  INV_X1    g0128(.A(G200), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n306), .B2(new_n318), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(new_n284), .A3(new_n295), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT17), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n331), .A2(new_n284), .A3(KEYINPUT17), .A4(new_n295), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n324), .A2(new_n327), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n289), .A2(new_n202), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n338), .A2(new_n294), .B1(new_n202), .B2(new_n293), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n217), .A2(G33), .ZN(new_n340));
  INV_X1    g0140(.A(G150), .ZN(new_n341));
  INV_X1    g0141(.A(new_n269), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n290), .A2(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n217), .B1(new_n201), .B2(new_n202), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n283), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT9), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT75), .ZN(new_n349));
  NOR2_X1   g0149(.A1(G222), .A2(G1698), .ZN(new_n350));
  INV_X1    g0150(.A(G1698), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(G223), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n275), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n310), .B(new_n353), .C1(G77), .C2(new_n275), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n298), .A2(new_n301), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(G226), .A3(new_n302), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n304), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G190), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n339), .A2(KEYINPUT9), .A3(new_n345), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT76), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(G200), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n359), .A2(new_n360), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n349), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT10), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n357), .A2(G179), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n357), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n346), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n365), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n298), .A2(new_n301), .A3(G238), .A4(new_n302), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n304), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(G33), .A2(G97), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(G226), .A2(G1698), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n241), .B2(G1698), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n375), .B1(new_n377), .B2(new_n275), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n307), .B1(new_n297), .B2(new_n282), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n214), .A2(KEYINPUT71), .A3(new_n300), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n378), .A2(KEYINPUT77), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT77), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n241), .A2(G1698), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(G226), .B2(G1698), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n374), .B1(new_n385), .B2(new_n277), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n386), .B2(new_n310), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n373), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT13), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT77), .B1(new_n378), .B2(new_n381), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n386), .A2(new_n310), .A3(new_n383), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT13), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(new_n373), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G200), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n293), .A2(new_n266), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n397), .B(KEYINPUT12), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n294), .A2(G68), .A3(new_n288), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT78), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n342), .A2(new_n202), .B1(new_n217), .B2(G68), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n340), .A2(new_n203), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n283), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT11), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n400), .B2(new_n401), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n389), .A2(G190), .A3(new_n394), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n396), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n408), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n392), .A2(new_n393), .A3(new_n373), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n393), .B1(new_n392), .B2(new_n373), .ZN(new_n414));
  OAI21_X1  g0214(.A(G169), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n389), .A2(G179), .A3(new_n394), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(G169), .C1(new_n413), .C2(new_n414), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n411), .B1(new_n412), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n275), .A2(G238), .A3(G1698), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n275), .A2(G232), .A3(new_n351), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n422), .B(new_n423), .C1(new_n207), .C2(new_n275), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n310), .ZN(new_n425));
  INV_X1    g0225(.A(G179), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n355), .A2(G244), .A3(new_n302), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n304), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n293), .A2(new_n203), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT73), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n290), .A2(new_n342), .B1(new_n217), .B2(new_n203), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n340), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n283), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n294), .A2(G77), .A3(new_n288), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n430), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n425), .A2(new_n304), .A3(new_n427), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n428), .B(new_n436), .C1(new_n437), .C2(G169), .ZN(new_n438));
  INV_X1    g0238(.A(new_n436), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n425), .A2(G190), .A3(new_n304), .A4(new_n427), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(new_n437), .C2(new_n329), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(new_n442), .B(KEYINPUT74), .ZN(new_n443));
  AND4_X1   g0243(.A1(new_n337), .A2(new_n371), .A3(new_n421), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n283), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n216), .A2(G33), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n292), .A4(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n292), .A2(new_n448), .A3(new_n282), .A4(new_n281), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n451), .A3(G107), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n292), .A2(G107), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT25), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT22), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(new_n217), .A3(G87), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n277), .A2(KEYINPUT84), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT84), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n316), .A2(KEYINPUT22), .A3(G20), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n459), .B1(new_n275), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  AOI211_X1 g0262(.A(G20), .B(new_n316), .C1(new_n258), .C2(new_n259), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(new_n456), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT23), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n217), .B2(G107), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G116), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n466), .A2(new_n467), .B1(new_n469), .B2(new_n217), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT85), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n446), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT85), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT84), .B1(new_n277), .B2(new_n457), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n275), .A2(new_n459), .A3(new_n460), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n258), .A2(new_n259), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(new_n217), .A3(G87), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n477), .B1(KEYINPUT22), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n470), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n474), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n464), .A2(KEYINPUT85), .A3(new_n470), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(KEYINPUT24), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n455), .B1(new_n473), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT87), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n216), .B(G45), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n355), .A2(new_n486), .A3(G264), .A4(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n298), .A3(G264), .A4(new_n301), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT87), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n253), .A2(KEYINPUT79), .A3(G33), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n275), .B2(new_n257), .ZN(new_n494));
  INV_X1    g0294(.A(G250), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n351), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(G257), .B2(new_n351), .ZN(new_n497));
  INV_X1    g0297(.A(G294), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n494), .A2(new_n497), .B1(new_n255), .B2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n490), .A2(new_n492), .B1(new_n499), .B2(new_n310), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n216), .A2(G45), .ZN(new_n501));
  INV_X1    g0301(.A(new_n488), .ZN(new_n502));
  NAND2_X1  g0302(.A1(KEYINPUT5), .A2(G41), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n504), .A2(G274), .A3(new_n298), .A4(new_n301), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n329), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n500), .A2(new_n505), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n506), .B1(new_n508), .B2(G190), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n485), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT86), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n473), .A2(new_n484), .ZN(new_n512));
  INV_X1    g0312(.A(new_n455), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI211_X1 g0314(.A(KEYINPUT86), .B(new_n455), .C1(new_n473), .C2(new_n484), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n367), .B1(new_n500), .B2(new_n505), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n426), .B2(new_n507), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n510), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n225), .A2(G1698), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n522), .B1(new_n494), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n254), .A2(new_n256), .A3(G250), .A4(G1698), .ZN(new_n526));
  AND2_X1   g0326(.A1(KEYINPUT4), .A2(G244), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n254), .A2(new_n256), .A3(new_n527), .A4(new_n351), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G283), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n381), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n489), .A2(new_n298), .A3(G257), .A4(new_n301), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n505), .A2(new_n533), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n532), .A2(new_n358), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n207), .B1(new_n276), .B2(new_n278), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n269), .A2(G77), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT6), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n538), .A2(new_n206), .A3(G107), .ZN(new_n539));
  XNOR2_X1  g0339(.A(G97), .B(G107), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n537), .B1(new_n541), .B2(new_n217), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n283), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n449), .A2(new_n451), .A3(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n293), .A2(new_n206), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n535), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT82), .B1(new_n532), .B2(new_n534), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT4), .B1(new_n478), .B2(new_n523), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n310), .B1(new_n550), .B2(new_n530), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT82), .ZN(new_n552));
  INV_X1    g0352(.A(new_n534), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n554), .A3(G200), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n551), .A2(new_n553), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n367), .B1(new_n543), .B2(new_n546), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n532), .A2(new_n534), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n426), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n548), .A2(new_n555), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT83), .ZN(new_n561));
  AOI211_X1 g0361(.A(G20), .B(new_n266), .C1(new_n258), .C2(new_n259), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT19), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G97), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n340), .A2(new_n564), .ZN(new_n565));
  OAI22_X1  g0365(.A1(new_n375), .A2(G20), .B1(new_n208), .B2(G87), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n561), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n478), .A2(new_n217), .A3(G68), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G97), .A2(G107), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(new_n316), .B1(new_n374), .B2(new_n217), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n571), .A2(new_n563), .B1(new_n340), .B2(new_n564), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n569), .A2(KEYINPUT83), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n568), .A2(new_n283), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n432), .A2(new_n293), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n449), .A2(new_n451), .A3(G87), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n225), .A2(G1698), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(G238), .B2(G1698), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n259), .B2(new_n258), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n310), .B1(new_n580), .B2(new_n469), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n501), .A2(new_n495), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n501), .A2(G274), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n355), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n329), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n581), .A2(new_n584), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n585), .B1(G190), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n432), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n449), .A2(new_n451), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n574), .A2(new_n589), .A3(new_n575), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n581), .A2(new_n426), .A3(new_n584), .ZN(new_n591));
  AOI21_X1  g0391(.A(G169), .B1(new_n581), .B2(new_n584), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n577), .A2(new_n587), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n560), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n226), .A2(G1698), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(G257), .B2(G1698), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n478), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G303), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n275), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n381), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n489), .A2(new_n298), .A3(G270), .A4(new_n301), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n505), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(G116), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n281), .A2(new_n282), .B1(G20), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n529), .B(new_n217), .C1(G33), .C2(new_n206), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(KEYINPUT20), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT20), .B1(new_n609), .B2(new_n610), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n293), .A2(new_n608), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n450), .B2(new_n608), .ZN(new_n616));
  OAI21_X1  g0416(.A(G169), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n596), .B1(new_n607), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(G200), .B1(new_n604), .B2(new_n606), .ZN(new_n619));
  INV_X1    g0419(.A(new_n616), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n613), .B2(new_n612), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n598), .B1(new_n259), .B2(new_n258), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n310), .B1(new_n623), .B2(new_n602), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(G190), .A3(new_n505), .A4(new_n605), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n619), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n505), .A3(new_n605), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n627), .A2(new_n621), .A3(KEYINPUT21), .A4(G169), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n607), .A2(G179), .A3(new_n621), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n618), .A2(new_n626), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NOR4_X1   g0431(.A1(new_n445), .A2(new_n521), .A3(new_n595), .A4(new_n631), .ZN(G372));
  INV_X1    g0432(.A(KEYINPUT89), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n324), .A2(new_n327), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n419), .A2(new_n417), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n418), .B1(new_n395), .B2(G169), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n412), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n411), .B2(new_n438), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n334), .A2(new_n335), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(new_n365), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n633), .B1(new_n641), .B2(new_n370), .ZN(new_n642));
  OAI211_X1 g0442(.A(KEYINPUT89), .B(new_n369), .C1(new_n640), .C2(new_n365), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n482), .A2(KEYINPUT24), .A3(new_n483), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n283), .B1(new_n482), .B2(KEYINPUT24), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n513), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT88), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n648), .A3(new_n519), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n517), .B1(new_n508), .B2(G179), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT88), .B1(new_n485), .B2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n618), .A2(new_n628), .A3(new_n629), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n510), .A2(new_n595), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n577), .A2(new_n587), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n590), .A2(new_n593), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n557), .A2(new_n559), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n656), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n660), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n594), .A2(new_n662), .A3(KEYINPUT26), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n661), .A2(new_n663), .B1(new_n590), .B2(new_n593), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n655), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n444), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n644), .A2(new_n666), .ZN(G369));
  NAND3_X1  g0467(.A1(new_n216), .A2(new_n217), .A3(G13), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT27), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n216), .A3(new_n217), .A4(G13), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  OR3_X1    g0473(.A1(new_n672), .A2(KEYINPUT90), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT90), .B1(new_n672), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n516), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n520), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n516), .A2(new_n519), .A3(new_n676), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n652), .ZN(new_n681));
  INV_X1    g0481(.A(new_n676), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n622), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n631), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n680), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT91), .Z(new_n689));
  AOI21_X1  g0489(.A(new_n676), .B1(new_n649), .B2(new_n651), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n681), .A2(new_n682), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT92), .Z(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n690), .B1(new_n680), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n220), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n212), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT28), .Z(new_n702));
  NAND2_X1  g0502(.A1(new_n665), .A2(new_n682), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n485), .A2(new_n509), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(new_n560), .A3(new_n594), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n647), .A2(KEYINPUT86), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n485), .A2(new_n511), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(new_n709), .A3(new_n519), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n707), .B1(new_n710), .B2(new_n652), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n661), .A2(new_n663), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n658), .ZN(new_n713));
  OAI211_X1 g0513(.A(KEYINPUT29), .B(new_n682), .C1(new_n711), .C2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n705), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  AND4_X1   g0516(.A1(new_n560), .A2(new_n594), .A3(new_n630), .A4(new_n682), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n710), .A2(new_n706), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n607), .A2(G179), .A3(new_n551), .A4(new_n553), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n500), .A2(new_n586), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n497), .B1(new_n259), .B2(new_n258), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n255), .A2(new_n498), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n310), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n491), .A2(KEYINPUT87), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n491), .A2(KEYINPUT87), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n581), .A2(new_n584), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n627), .A2(new_n426), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n731), .A4(new_n558), .ZN(new_n732));
  AOI21_X1  g0532(.A(G179), .B1(new_n581), .B2(new_n584), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n507), .A2(new_n556), .A3(new_n627), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n722), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(KEYINPUT93), .A2(KEYINPUT31), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(new_n676), .A3(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n735), .A2(new_n676), .ZN(new_n738));
  XNOR2_X1  g0538(.A(KEYINPUT93), .B(KEYINPUT31), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n716), .B1(new_n718), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n715), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n702), .B1(new_n743), .B2(new_n216), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT94), .Z(G364));
  INV_X1    g0545(.A(G13), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n216), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n697), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n282), .B1(G20), .B2(new_n367), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G179), .A2(G200), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT95), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n217), .A2(G190), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G159), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT32), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n217), .B1(new_n756), .B2(G190), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n206), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n217), .A2(new_n426), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G190), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n329), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n765), .A2(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n202), .A2(new_n767), .B1(new_n769), .B2(new_n265), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n764), .A2(new_n358), .A3(new_n329), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n764), .A2(new_n358), .A3(G200), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n275), .B1(new_n771), .B2(new_n203), .C1(new_n266), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n217), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G190), .A3(G200), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(new_n358), .A3(G200), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n316), .A2(new_n775), .B1(new_n776), .B2(new_n207), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n763), .A2(new_n770), .A3(new_n773), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G311), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT33), .B(G317), .Z(new_n780));
  OAI221_X1 g0580(.A(new_n277), .B1(new_n771), .B2(new_n779), .C1(new_n772), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n758), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(new_n782), .B2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(new_n762), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G294), .ZN(new_n785));
  INV_X1    g0585(.A(new_n775), .ZN(new_n786));
  INV_X1    g0586(.A(new_n776), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n786), .A2(G303), .B1(new_n787), .B2(G283), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n768), .A2(G322), .B1(new_n766), .B2(G326), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n783), .A2(new_n785), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT96), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n761), .A2(new_n778), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n753), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n752), .ZN(new_n798));
  INV_X1    g0598(.A(G45), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n213), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n696), .A2(new_n478), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n800), .B(new_n801), .C1(new_n799), .C2(new_n248), .ZN(new_n802));
  INV_X1    g0602(.A(G355), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n220), .A2(new_n275), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n802), .B1(G116), .B2(new_n220), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n751), .B(new_n794), .C1(new_n798), .C2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  INV_X1    g0607(.A(new_n797), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n685), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n687), .A2(new_n750), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(G330), .B2(new_n685), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G396));
  NAND3_X1  g0613(.A1(new_n676), .A2(new_n436), .A3(KEYINPUT98), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT98), .B1(new_n676), .B2(new_n436), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n817), .A2(KEYINPUT99), .A3(new_n438), .A4(new_n441), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT99), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n815), .A2(new_n816), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n442), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n665), .A2(new_n682), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n676), .B1(new_n655), .B2(new_n664), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n438), .A2(new_n682), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n818), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n823), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n827), .A2(new_n742), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n750), .B1(new_n827), .B2(new_n742), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n753), .A2(new_n796), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n750), .B1(G77), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n772), .ZN(new_n833));
  INV_X1    g0633(.A(new_n771), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G150), .A2(new_n833), .B1(new_n834), .B2(G159), .ZN(new_n835));
  INV_X1    g0635(.A(G137), .ZN(new_n836));
  INV_X1    g0636(.A(G143), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(new_n836), .B2(new_n767), .C1(new_n837), .C2(new_n769), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT34), .Z(new_n839));
  NOR2_X1   g0639(.A1(new_n776), .A2(new_n266), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n494), .B(new_n840), .C1(G50), .C2(new_n786), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n265), .B2(new_n762), .C1(new_n842), .C2(new_n758), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n316), .A2(new_n776), .B1(new_n775), .B2(new_n207), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n498), .A2(new_n769), .B1(new_n767), .B2(new_n601), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n758), .A2(new_n779), .ZN(new_n846));
  INV_X1    g0646(.A(G283), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n277), .B1(new_n771), .B2(new_n608), .C1(new_n847), .C2(new_n772), .ZN(new_n848));
  OR4_X1    g0648(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n839), .A2(new_n843), .B1(new_n763), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n832), .B1(new_n850), .B2(new_n752), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n826), .B2(new_n796), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT100), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n830), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G384));
  NOR2_X1   g0655(.A1(new_n747), .A2(new_n216), .ZN(new_n856));
  INV_X1    g0656(.A(new_n295), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n266), .B1(new_n260), .B2(KEYINPUT7), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n271), .B1(new_n858), .B2(new_n263), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n446), .B1(new_n859), .B2(KEYINPUT16), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n264), .A2(new_n272), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n274), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n857), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n332), .B1(new_n863), .B2(new_n672), .ZN(new_n864));
  INV_X1    g0664(.A(new_n322), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT103), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n868), .B1(new_n325), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n672), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n296), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n332), .B(new_n872), .C1(new_n323), .C2(KEYINPUT103), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n867), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n863), .A2(new_n672), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n336), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n874), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n323), .A2(new_n872), .A3(new_n332), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n870), .B2(new_n873), .ZN(new_n880));
  INV_X1    g0680(.A(new_n872), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n336), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT40), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT104), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n885), .A2(KEYINPUT31), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n735), .A2(new_n676), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n735), .B2(new_n676), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n718), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n818), .A2(new_n821), .A3(new_n825), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n412), .A2(new_n676), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n637), .A2(new_n410), .A3(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n412), .B(new_n676), .C1(new_n411), .C2(new_n420), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n884), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT105), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n887), .A2(new_n888), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n520), .B2(new_n717), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n637), .A2(new_n410), .A3(new_n892), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n892), .B1(new_n637), .B2(new_n410), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n826), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n898), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n874), .A2(new_n876), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n874), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n890), .A2(new_n895), .A3(KEYINPUT105), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n904), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n897), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n445), .B2(new_n900), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n913), .A2(new_n444), .A3(new_n890), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(G330), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n444), .A2(new_n705), .A3(new_n714), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n644), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n894), .A2(new_n893), .ZN(new_n920));
  INV_X1    g0720(.A(new_n822), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n676), .B(new_n921), .C1(new_n655), .C2(new_n664), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n438), .A2(new_n676), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n909), .B(new_n920), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n877), .B2(new_n883), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n420), .A2(new_n412), .A3(new_n682), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n634), .A2(new_n672), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n924), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n919), .B(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n856), .B1(new_n917), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n933), .B2(new_n917), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n212), .A2(new_n203), .A3(new_n267), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n266), .A2(G50), .ZN(new_n937));
  OAI211_X1 g0737(.A(G1), .B(new_n746), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT101), .Z(new_n939));
  INV_X1    g0739(.A(new_n541), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT35), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(KEYINPUT35), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n282), .A2(new_n217), .A3(new_n608), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT36), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT102), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n935), .A2(new_n947), .ZN(G367));
  NAND2_X1  g0748(.A1(new_n547), .A2(new_n676), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n560), .A2(new_n949), .B1(new_n662), .B2(new_n676), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n680), .A2(new_n693), .A3(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n952), .A2(KEYINPUT42), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n710), .B1(new_n555), .B2(new_n548), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(new_n662), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n952), .A2(KEYINPUT42), .B1(new_n682), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n957), .A2(KEYINPUT106), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(KEYINPUT106), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n577), .A2(new_n682), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n594), .B(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n960), .B1(KEYINPUT43), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n689), .A2(new_n950), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n962), .B(KEYINPUT43), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n958), .B2(new_n959), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n964), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n966), .B1(new_n964), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n688), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n680), .A2(new_n687), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n973), .A2(new_n692), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n743), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n692), .B1(new_n973), .B2(new_n974), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT44), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n694), .A2(new_n979), .A3(new_n951), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(new_n694), .B2(new_n951), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n694), .A2(new_n951), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n694), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n982), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n689), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n978), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n982), .A2(new_n987), .A3(new_n689), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n743), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n697), .B(KEYINPUT41), .Z(new_n993));
  OAI21_X1  g0793(.A(new_n748), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n972), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n801), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n239), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n798), .B1(new_n220), .B2(new_n432), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n750), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n769), .A2(new_n341), .B1(new_n775), .B2(new_n265), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G50), .A2(new_n834), .B1(new_n833), .B2(G159), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n837), .B2(new_n767), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(G137), .C2(new_n782), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n776), .A2(new_n203), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(new_n277), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT108), .Z(new_n1006));
  OAI211_X1 g0806(.A(new_n1003), .B(new_n1006), .C1(new_n266), .C2(new_n762), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n601), .A2(new_n769), .B1(new_n767), .B2(new_n779), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n776), .A2(new_n206), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n494), .B1(new_n847), .B2(new_n771), .C1(new_n498), .C2(new_n772), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G317), .B2(new_n782), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n775), .A2(new_n608), .ZN(new_n1013));
  XOR2_X1   g0813(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(KEYINPUT46), .B2(new_n1013), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n784), .A2(G107), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1010), .A2(new_n1012), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1007), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT47), .Z(new_n1020));
  NOR2_X1   g0820(.A1(new_n1020), .A2(new_n753), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n999), .B(new_n1021), .C1(new_n797), .C2(new_n962), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n995), .A2(new_n1023), .ZN(G387));
  NAND2_X1  g0824(.A1(new_n975), .A2(new_n977), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(new_n748), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n678), .A2(new_n679), .A3(new_n797), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n804), .A2(new_n699), .B1(G107), .B2(new_n220), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n244), .A2(new_n799), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n699), .B(new_n799), .C1(new_n266), .C2(new_n203), .ZN(new_n1030));
  XOR2_X1   g0830(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1031));
  NOR3_X1   g0831(.A1(new_n1031), .A2(G50), .A3(new_n290), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1031), .B1(G50), .B2(new_n290), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n996), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1028), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n798), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n750), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n772), .A2(new_n290), .B1(new_n771), .B2(new_n266), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n494), .B(new_n1039), .C1(new_n782), .C2(G150), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n784), .A2(new_n588), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1009), .B1(G77), .B2(new_n786), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n768), .A2(G50), .B1(new_n766), .B2(G159), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT110), .Z(new_n1045));
  NAND2_X1  g0845(.A1(new_n782), .A2(G326), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n478), .B1(G116), .B2(new_n787), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n762), .A2(new_n847), .B1(new_n498), .B2(new_n775), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G303), .A2(new_n834), .B1(new_n833), .B2(G311), .ZN(new_n1049));
  INV_X1    g0849(.A(G322), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n767), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G317), .B2(new_n768), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT111), .Z(new_n1053));
  INV_X1    g0853(.A(KEYINPUT48), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1048), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n1054), .B2(new_n1053), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT49), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1046), .B(new_n1047), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1045), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1038), .B1(new_n1060), .B2(new_n752), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1026), .B1(new_n1027), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1025), .A2(new_n743), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n697), .B(KEYINPUT112), .Z(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n978), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1062), .A2(new_n1065), .ZN(G393));
  INV_X1    g0866(.A(new_n1064), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n990), .B2(new_n991), .ZN(new_n1068));
  AOI21_X1  g0868(.A(KEYINPUT113), .B1(new_n988), .B2(new_n989), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(new_n991), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n978), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n798), .B1(new_n206), .B2(new_n220), .C1(new_n996), .C2(new_n251), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n762), .A2(new_n203), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n782), .A2(G143), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n786), .A2(G68), .B1(new_n787), .B2(G87), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n290), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1077), .A2(new_n834), .B1(new_n833), .B2(G50), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1075), .A2(new_n478), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n768), .A2(G159), .B1(new_n766), .B2(G150), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT115), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT114), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1074), .B(new_n1079), .C1(new_n1082), .C2(KEYINPUT51), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n784), .A2(G116), .B1(G303), .B2(new_n833), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(KEYINPUT116), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n776), .A2(new_n207), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n277), .B1(new_n771), .B2(new_n498), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1088), .B(new_n1089), .C1(G283), .C2(new_n786), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1050), .B2(new_n758), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n768), .A2(G311), .B1(new_n766), .B2(G317), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT52), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1087), .A2(new_n1091), .A3(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1083), .A2(new_n1084), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n750), .B(new_n1073), .C1(new_n1095), .C2(new_n753), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n797), .B2(new_n950), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1070), .B2(new_n749), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1072), .A2(new_n1098), .ZN(G390));
  NAND2_X1  g0899(.A1(new_n926), .A2(new_n927), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n920), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n923), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1101), .B1(new_n823), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1100), .B1(new_n1103), .B2(new_n929), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n682), .B(new_n822), .C1(new_n711), .C2(new_n713), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n1102), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n920), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n873), .A2(new_n870), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1108), .A2(new_n879), .B1(new_n336), .B2(new_n881), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n908), .B1(new_n1109), .B2(KEYINPUT38), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1110), .A2(new_n928), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n741), .A2(new_n826), .A3(new_n920), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1104), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n923), .B1(new_n824), .B2(new_n822), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n928), .B1(new_n1115), .B2(new_n1101), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1116), .A2(new_n1100), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n716), .B1(new_n889), .B2(new_n718), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n895), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1114), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n444), .A2(new_n1118), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n918), .A2(new_n644), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1113), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n920), .B1(new_n1118), .B2(new_n826), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n920), .B1(new_n741), .B2(new_n826), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n716), .B(new_n891), .C1(new_n718), .C2(new_n740), .ZN(new_n1129));
  OAI21_X1  g0929(.A(KEYINPUT117), .B1(new_n1129), .B2(new_n920), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1128), .A2(new_n1130), .A3(new_n1119), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1115), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1125), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1120), .B1(new_n1122), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1119), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1136), .A2(new_n928), .B1(new_n926), .B2(new_n927), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1110), .A2(new_n928), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n1106), .B2(new_n920), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1135), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1119), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1129), .A2(KEYINPUT117), .A3(new_n920), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1132), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1122), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1140), .A2(new_n1145), .A3(new_n1114), .A4(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1134), .A2(new_n1064), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1140), .A2(new_n749), .A3(new_n1114), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n750), .B1(new_n1077), .B2(new_n831), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n608), .A2(new_n769), .B1(new_n767), .B2(new_n847), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n840), .B(new_n1151), .C1(G87), .C2(new_n786), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n277), .B1(new_n771), .B2(new_n206), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G107), .B2(new_n833), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(new_n498), .C2(new_n758), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n775), .A2(new_n341), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT53), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT54), .B(G143), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n275), .B1(new_n771), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G137), .B2(new_n833), .ZN(new_n1160));
  INV_X1    g0960(.A(G125), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1157), .B(new_n1160), .C1(new_n1161), .C2(new_n758), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n768), .A2(G132), .B1(new_n787), .B2(G50), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n766), .A2(G128), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n762), .C2(new_n759), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n1155), .A2(new_n1074), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1150), .B1(new_n1166), .B2(new_n752), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1100), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n1168), .B2(new_n796), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1148), .A2(new_n1149), .A3(new_n1169), .ZN(G378));
  OAI21_X1  g0970(.A(new_n750), .B1(G50), .B2(new_n831), .ZN(new_n1171));
  INV_X1    g0971(.A(G41), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n494), .A2(new_n1172), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n206), .A2(new_n772), .B1(new_n771), .B2(new_n432), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(G77), .C2(new_n786), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n847), .B2(new_n758), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n762), .A2(new_n266), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n776), .A2(new_n265), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n207), .A2(new_n769), .B1(new_n767), .B2(new_n608), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT118), .Z(new_n1181));
  OR2_X1    g0981(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(KEYINPUT58), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1173), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n255), .B(new_n1172), .C1(new_n776), .C2(new_n759), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT119), .B(G124), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n782), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT120), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n772), .A2(new_n842), .B1(new_n771), .B2(new_n836), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1158), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n786), .B2(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n768), .A2(G128), .B1(new_n766), .B2(G125), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(new_n341), .C2(new_n762), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1188), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1171), .B1(new_n1197), .B2(new_n752), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n346), .A2(new_n871), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n371), .B(new_n1199), .Z(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1200), .B(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1198), .B1(new_n1202), .B2(new_n796), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT121), .Z(new_n1204));
  AND3_X1   g1004(.A1(new_n913), .A2(G330), .A3(new_n932), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n932), .B1(new_n913), .B2(G330), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1202), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n911), .A2(new_n912), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n897), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1208), .A2(G330), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n932), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1201), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1200), .B(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n913), .A2(G330), .A3(new_n932), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n748), .B1(new_n1207), .B2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1204), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1146), .B1(new_n1120), .B2(new_n1133), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1205), .A2(new_n1206), .A3(new_n1202), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1214), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1219), .B(KEYINPUT57), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT122), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n1223), .A3(new_n1064), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT123), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1207), .A2(new_n1216), .B1(new_n1147), .B2(new_n1146), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n1226), .B2(KEYINPUT57), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT57), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(KEYINPUT123), .A3(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1224), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1223), .B1(new_n1222), .B2(new_n1064), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1218), .B1(new_n1231), .B2(new_n1232), .ZN(G375));
  NOR2_X1   g1033(.A1(new_n1133), .A2(new_n1122), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(new_n993), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1143), .A2(new_n1122), .A3(new_n1144), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT124), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT124), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1133), .A2(new_n1238), .A3(new_n1122), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1235), .A2(new_n1237), .A3(new_n1239), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT125), .Z(new_n1241));
  NAND2_X1  g1041(.A1(new_n1101), .A2(new_n795), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n750), .B1(G68), .B2(new_n831), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n847), .A2(new_n769), .B1(new_n767), .B2(new_n498), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1004), .B(new_n1244), .C1(G97), .C2(new_n786), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n782), .A2(G303), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n277), .B1(new_n772), .B2(new_n608), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G107), .B2(new_n834), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1041), .A3(new_n1246), .A4(new_n1248), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n842), .A2(new_n767), .B1(new_n769), .B2(new_n836), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1178), .B(new_n1250), .C1(G159), .C2(new_n786), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n782), .A2(G128), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1190), .A2(new_n833), .B1(new_n834), .B2(G150), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1251), .A2(new_n478), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n762), .A2(new_n202), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1249), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1243), .B1(new_n1256), .B2(new_n752), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1145), .A2(new_n749), .B1(new_n1242), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1241), .A2(new_n1258), .ZN(G381));
  NAND3_X1  g1059(.A1(new_n1062), .A2(new_n812), .A3(new_n1065), .ZN(new_n1260));
  OR4_X1    g1060(.A1(G384), .A2(G390), .A3(G378), .A4(new_n1260), .ZN(new_n1261));
  OR4_X1    g1061(.A1(G387), .A2(new_n1261), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1062(.A(G378), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n673), .A2(G213), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G407), .B(G213), .C1(G375), .C2(new_n1266), .ZN(G409));
  INV_X1    g1067(.A(KEYINPUT127), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G393), .A2(G396), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1260), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1072), .A2(new_n1098), .A3(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1072), .B2(new_n1098), .ZN(new_n1272));
  OAI21_X1  g1072(.A(G387), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1270), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G390), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1022), .B1(new_n972), .B2(new_n994), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1072), .A2(new_n1098), .A3(new_n1270), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1273), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT61), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G378), .B(new_n1218), .C1(new_n1231), .C2(new_n1232), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1218), .B1(new_n993), .B2(new_n1228), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1263), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1265), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1265), .A2(G2897), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT60), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1237), .B(new_n1239), .C1(new_n1234), .C2(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1236), .A2(new_n1288), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(new_n1067), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(G384), .B1(new_n1292), .B2(new_n1258), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1258), .ZN(new_n1294));
  AOI211_X1 g1094(.A(new_n854), .B(new_n1294), .C1(new_n1289), .C2(new_n1291), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1285), .B(new_n1287), .C1(new_n1293), .C2(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1286), .B1(new_n1297), .B2(KEYINPUT126), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(KEYINPUT126), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1296), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1280), .B1(new_n1284), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(new_n1284), .B2(new_n1297), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1297), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n1265), .B(new_n1305), .C1(new_n1281), .C2(new_n1283), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1302), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1279), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1284), .A2(KEYINPUT63), .A3(new_n1297), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1309), .B(new_n1280), .C1(new_n1284), .C2(new_n1300), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1279), .B1(new_n1306), .B2(KEYINPUT63), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1268), .B1(new_n1308), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1301), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1284), .A2(new_n1297), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1314), .A2(new_n1317), .A3(new_n1279), .A4(new_n1309), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1315), .A2(KEYINPUT62), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1319), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1318), .B(KEYINPUT127), .C1(new_n1320), .C2(new_n1279), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1313), .A2(new_n1321), .ZN(G405));
  NAND2_X1  g1122(.A1(G375), .A2(new_n1263), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1281), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(new_n1305), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1325), .B(new_n1279), .ZN(G402));
endmodule


