//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(KEYINPUT64), .A2(G68), .ZN(new_n217));
  NAND2_X1  g0017(.A1(KEYINPUT64), .A2(G68), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT65), .B(G244), .Z(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  AOI21_X1  g0047(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G226), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G41), .ZN(new_n254));
  OAI211_X1 g0054(.A(G1), .B(G13), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n250), .A2(new_n255), .A3(G274), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n252), .A2(KEYINPUT68), .A3(new_n256), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G222), .A2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G223), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n265), .B(new_n248), .C1(G77), .C2(new_n261), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n259), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G190), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(G200), .B2(new_n267), .ZN(new_n270));
  INV_X1    g0070(.A(G13), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n271), .A2(new_n206), .A3(G1), .ZN(new_n272));
  INV_X1    g0072(.A(G50), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n214), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n206), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G150), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n277), .A2(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n206), .B1(new_n201), .B2(new_n273), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n276), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n271), .A2(G1), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT69), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n288), .A2(new_n289), .B1(new_n205), .B2(G20), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n290), .B1(new_n289), .B2(new_n288), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n274), .B(new_n284), .C1(new_n291), .C2(new_n273), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n293), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n270), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n267), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n299), .B(new_n292), .C1(G179), .C2(new_n267), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n219), .A2(new_n206), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n281), .A2(new_n273), .B1(new_n278), .B2(new_n221), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n276), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT11), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  INV_X1    g0107(.A(new_n288), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(G68), .C1(G1), .C2(new_n206), .ZN(new_n309));
  INV_X1    g0109(.A(G68), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT12), .B1(new_n272), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n286), .A2(KEYINPUT12), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n302), .B2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n306), .A2(new_n307), .A3(new_n309), .A4(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n255), .A2(G238), .A3(new_n249), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n256), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT13), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n263), .A2(G232), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n261), .B(new_n319), .C1(G226), .C2(G1698), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G97), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n317), .B(new_n318), .C1(new_n322), .C2(new_n255), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n255), .B1(new_n320), .B2(new_n321), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT13), .B1(new_n324), .B2(new_n316), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT14), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(G169), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n323), .A2(new_n325), .A3(G179), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n327), .B1(new_n326), .B2(G169), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n314), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n326), .A2(G200), .ZN(new_n333));
  INV_X1    g0133(.A(new_n314), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n333), .B(new_n334), .C1(new_n268), .C2(new_n326), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT71), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n277), .B(KEYINPUT70), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n280), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT15), .B(G87), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n253), .A2(G20), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n341), .A2(new_n342), .B1(G20), .B2(G77), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n285), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(G77), .B1(new_n206), .B2(G1), .ZN(new_n345));
  OAI22_X1  g0145(.A1(new_n288), .A2(new_n345), .B1(G77), .B2(new_n287), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G274), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n248), .A2(new_n348), .A3(new_n249), .ZN(new_n349));
  NOR3_X1   g0149(.A1(new_n222), .A2(new_n248), .A3(new_n250), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n261), .A2(G238), .A3(G1698), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n261), .A2(G232), .A3(new_n263), .ZN(new_n352));
  INV_X1    g0152(.A(G107), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n351), .B(new_n352), .C1(new_n353), .C2(new_n261), .ZN(new_n354));
  AOI211_X1 g0154(.A(new_n349), .B(new_n350), .C1(new_n354), .C2(new_n248), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n347), .B1(G190), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G200), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(new_n355), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n355), .A2(G169), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n359), .A2(new_n347), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n301), .A2(new_n337), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n277), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(new_n272), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n291), .B2(new_n366), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT72), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT72), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(G33), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n369), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT7), .B1(new_n374), .B2(G20), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(new_n372), .A3(new_n373), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(new_n206), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(G68), .A3(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(KEYINPUT64), .A2(G68), .ZN(new_n380));
  NOR2_X1   g0180(.A1(KEYINPUT64), .A2(G68), .ZN(new_n381));
  OAI21_X1  g0181(.A(G58), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n202), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G20), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT73), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n206), .B1(new_n382), .B2(new_n202), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(KEYINPUT73), .B1(G159), .B2(new_n280), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n379), .A2(KEYINPUT16), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n276), .ZN(new_n390));
  NOR3_X1   g0190(.A1(new_n261), .A2(new_n377), .A3(G20), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n371), .A2(G33), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n373), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT7), .B1(new_n393), .B2(new_n206), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n219), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n388), .A2(new_n386), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT74), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n390), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(KEYINPUT74), .A3(new_n397), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n368), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n349), .B1(G232), .B2(new_n251), .ZN(new_n402));
  OR2_X1    g0202(.A1(G223), .A2(G1698), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G226), .B2(new_n263), .ZN(new_n404));
  INV_X1    g0204(.A(G87), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n376), .A2(new_n404), .B1(new_n253), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n248), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G169), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n361), .B2(new_n408), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT18), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT74), .ZN(new_n413));
  INV_X1    g0213(.A(G58), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n217), .B2(new_n218), .ZN(new_n415));
  OAI211_X1 g0215(.A(KEYINPUT73), .B(G20), .C1(new_n415), .C2(new_n201), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n280), .A2(G159), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n219), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n377), .B1(new_n261), .B2(G20), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n393), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT73), .B1(new_n383), .B2(G20), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n418), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n413), .B1(new_n424), .B2(KEYINPUT16), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n425), .A2(new_n276), .A3(new_n400), .A4(new_n389), .ZN(new_n426));
  INV_X1    g0226(.A(new_n368), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n410), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n408), .A2(new_n268), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(G200), .B2(new_n408), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n426), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n426), .A2(new_n432), .A3(KEYINPUT17), .A4(new_n427), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n412), .A2(new_n430), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n365), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n205), .B(G45), .C1(new_n254), .C2(KEYINPUT5), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT5), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT76), .B1(new_n442), .B2(G41), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT76), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(new_n254), .A3(KEYINPUT5), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n441), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(new_n248), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G264), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n248), .A2(new_n348), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G250), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n263), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(G257), .B2(new_n263), .ZN(new_n453));
  INV_X1    g0253(.A(G294), .ZN(new_n454));
  OAI22_X1  g0254(.A1(new_n376), .A2(new_n453), .B1(new_n253), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n248), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n448), .A2(new_n450), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G179), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n298), .B2(new_n457), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n405), .A2(KEYINPUT22), .A3(G20), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n261), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT82), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT22), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n369), .A2(new_n372), .A3(new_n206), .A4(new_n373), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n405), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(new_n465), .B2(KEYINPUT81), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT81), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n464), .B2(new_n405), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n462), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n353), .A2(KEYINPUT23), .A3(G20), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT23), .B1(new_n353), .B2(G20), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G116), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n470), .A2(new_n471), .B1(G20), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT24), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n374), .A2(KEYINPUT81), .A3(new_n206), .A4(G87), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(KEYINPUT22), .A3(new_n468), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT82), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n461), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT24), .ZN(new_n480));
  INV_X1    g0280(.A(new_n473), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n285), .B1(new_n474), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT25), .B1(new_n272), .B2(new_n353), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n272), .A2(KEYINPUT25), .A3(new_n353), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n253), .A2(G1), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n272), .A2(new_n276), .A3(new_n487), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n485), .A2(new_n486), .B1(new_n488), .B2(G107), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n459), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n480), .B1(new_n479), .B2(new_n481), .ZN(new_n493));
  AOI211_X1 g0293(.A(KEYINPUT24), .B(new_n473), .C1(new_n476), .C2(new_n478), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n276), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n457), .A2(new_n357), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(G190), .B2(new_n457), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n489), .A3(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n491), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n492), .B1(new_n491), .B2(new_n498), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G238), .A2(G1698), .ZN(new_n502));
  INV_X1    g0302(.A(G244), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(G1698), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n504), .A2(new_n369), .A3(new_n372), .A4(new_n373), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT77), .B1(new_n505), .B2(new_n472), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n503), .A2(G1698), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(G238), .B2(G1698), .ZN(new_n508));
  OAI211_X1 g0308(.A(KEYINPUT77), .B(new_n472), .C1(new_n376), .C2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n248), .B1(new_n506), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G45), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(G1), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n449), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n255), .B(G250), .C1(G1), .C2(new_n512), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT78), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n472), .B1(new_n376), .B2(new_n508), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT77), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n255), .B1(new_n521), .B2(new_n509), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT78), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n522), .A2(new_n523), .A3(new_n516), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n298), .B1(new_n518), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n511), .A2(KEYINPUT78), .A3(new_n517), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n523), .B1(new_n522), .B2(new_n516), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(new_n361), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT19), .B1(new_n342), .B2(G97), .ZN(new_n529));
  INV_X1    g0329(.A(G97), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n405), .A2(new_n530), .A3(new_n353), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT79), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G87), .A2(G97), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT79), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n534), .A3(new_n353), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n206), .B1(new_n321), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n529), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n374), .A2(new_n206), .A3(G68), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n285), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT80), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n341), .A2(new_n287), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NOR4_X1   g0344(.A1(KEYINPUT79), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n534), .B1(new_n533), .B2(new_n353), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n529), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n464), .A2(new_n310), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n276), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n543), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT80), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n488), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n544), .A2(new_n553), .B1(new_n554), .B2(new_n340), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n525), .A2(new_n528), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G200), .B1(new_n518), .B2(new_n524), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n526), .A2(new_n527), .A3(G190), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n554), .A2(new_n405), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n542), .B1(new_n541), .B2(new_n543), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n551), .A2(KEYINPUT80), .A3(new_n552), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n557), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(G116), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G20), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n276), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G33), .A2(G283), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n568), .B(new_n206), .C1(G33), .C2(new_n530), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT20), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  AND4_X1   g0370(.A1(KEYINPUT20), .A2(new_n569), .A3(new_n276), .A4(new_n566), .ZN(new_n571));
  OR2_X1    g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n287), .A2(G116), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n488), .B2(G116), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n298), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  OR2_X1    g0375(.A1(G257), .A2(G1698), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(G264), .B2(new_n263), .ZN(new_n577));
  INV_X1    g0377(.A(G303), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n376), .A2(new_n577), .B1(new_n578), .B2(new_n261), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n248), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n443), .A2(new_n445), .ZN(new_n581));
  OAI211_X1 g0381(.A(G270), .B(new_n255), .C1(new_n581), .C2(new_n441), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n582), .A3(new_n450), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT21), .B1(new_n575), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n574), .B1(new_n570), .B2(new_n571), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n583), .A2(new_n585), .A3(KEYINPUT21), .A4(G169), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n582), .A2(new_n450), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n585), .A2(new_n587), .A3(G179), .A4(new_n580), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n585), .B1(new_n583), .B2(G200), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n268), .B2(new_n583), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n503), .A2(G1698), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT4), .B1(new_n374), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n595));
  AND2_X1   g0395(.A1(KEYINPUT4), .A2(G244), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n392), .A2(new_n373), .A3(new_n596), .A4(new_n263), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n568), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n248), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n447), .A2(G257), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n450), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n298), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n599), .A2(new_n361), .A3(new_n450), .A4(new_n600), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n353), .A2(KEYINPUT6), .A3(G97), .ZN(new_n604));
  XNOR2_X1  g0404(.A(G97), .B(G107), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT6), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n607), .A2(new_n206), .B1(new_n221), .B2(new_n281), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n353), .B1(new_n420), .B2(new_n421), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n608), .B1(KEYINPUT75), .B2(new_n609), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n609), .A2(KEYINPUT75), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n285), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n287), .A2(G97), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n488), .B2(G97), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n602), .B(new_n603), .C1(new_n612), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n601), .A2(G200), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n609), .A2(KEYINPUT75), .ZN(new_n618));
  INV_X1    g0418(.A(new_n608), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n609), .A2(KEYINPUT75), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n276), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n599), .A2(G190), .A3(new_n450), .A4(new_n600), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n617), .A2(new_n622), .A3(new_n614), .A4(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n590), .A2(new_n592), .A3(new_n616), .A4(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n564), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n440), .A2(new_n501), .A3(new_n626), .ZN(G372));
  AND2_X1   g0427(.A1(new_n412), .A2(new_n430), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n435), .A2(new_n436), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n332), .ZN(new_n631));
  INV_X1    g0431(.A(new_n363), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n335), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n628), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n297), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n635), .A2(new_n300), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n522), .A2(new_n516), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n637), .A2(new_n357), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT84), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n560), .A2(new_n561), .ZN(new_n641));
  INV_X1    g0441(.A(new_n559), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI211_X1 g0443(.A(KEYINPUT84), .B(new_n559), .C1(new_n560), .C2(new_n561), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n639), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT85), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT85), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n647), .B(new_n639), .C1(new_n643), .C2(new_n644), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n646), .A2(new_n558), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  INV_X1    g0450(.A(new_n616), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n555), .A2(new_n528), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n637), .A2(G169), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n649), .A2(new_n650), .A3(new_n651), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n495), .A2(new_n489), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT86), .B1(new_n584), .B2(new_n589), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n583), .A2(new_n585), .A3(G169), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT21), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT86), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(new_n586), .A4(new_n588), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n657), .A2(new_n459), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n616), .A2(new_n624), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n498), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n649), .A3(new_n655), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n556), .A2(new_n563), .A3(new_n651), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n655), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n656), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n636), .B1(new_n439), .B2(new_n674), .ZN(G369));
  NAND2_X1  g0475(.A1(new_n590), .A2(new_n592), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n286), .A2(new_n206), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(G213), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n585), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n677), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n658), .A2(new_n663), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n585), .A3(new_n683), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(G330), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n657), .ZN(new_n690));
  INV_X1    g0490(.A(new_n683), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n501), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n657), .A2(new_n459), .A3(new_n683), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n590), .A2(new_n683), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n501), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n657), .A2(new_n459), .A3(new_n691), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n694), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n209), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G1), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n532), .A2(new_n565), .A3(new_n535), .ZN(new_n704));
  OAI22_X1  g0504(.A1(new_n703), .A2(new_n704), .B1(new_n212), .B2(new_n702), .ZN(new_n705));
  XOR2_X1   g0505(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n706));
  XNOR2_X1  g0506(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n587), .A2(G179), .A3(new_n580), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n599), .A2(new_n600), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n448), .A2(new_n456), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n527), .A3(new_n526), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n711), .A2(KEYINPUT30), .A3(new_n527), .A4(new_n526), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n457), .A2(new_n361), .A3(new_n583), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n716), .B(new_n601), .C1(new_n522), .C2(new_n516), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n683), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n491), .A2(new_n498), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT83), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n491), .A2(new_n492), .A3(new_n498), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n626), .A3(new_n724), .A4(new_n691), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT89), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT89), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n501), .A2(new_n727), .A3(new_n626), .A4(new_n691), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n721), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G330), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT29), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n674), .B2(new_n683), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n669), .A2(new_n650), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n648), .A2(new_n558), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n642), .B1(new_n544), .B2(new_n553), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT84), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n562), .A2(new_n640), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n647), .B1(new_n739), .B2(new_n639), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n651), .B(new_n655), .C1(new_n735), .C2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n734), .B1(new_n741), .B2(new_n650), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n666), .B1(new_n491), .B2(new_n590), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n654), .B1(new_n743), .B2(new_n649), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT29), .A3(new_n691), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n731), .B1(new_n733), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n707), .B1(new_n747), .B2(G1), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT90), .Z(G364));
  NOR2_X1   g0549(.A1(new_n271), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n205), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n701), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n689), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n686), .A2(new_n688), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n756), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n214), .B1(G20), .B2(new_n298), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n206), .A2(new_n361), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n767), .A2(new_n268), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G322), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n357), .A2(G190), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n766), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g0572(.A(KEYINPUT33), .B(G317), .Z(new_n773));
  OAI22_X1  g0573(.A1(new_n769), .A2(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT93), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n268), .A2(new_n357), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n766), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n206), .A2(G179), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n771), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n778), .A2(G326), .B1(new_n781), .B2(G283), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G190), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n766), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n779), .A2(new_n783), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G311), .A2(new_n785), .B1(new_n787), .B2(G329), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n268), .A2(G179), .A3(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n206), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n789), .B1(G294), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n776), .A2(new_n779), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n393), .B1(new_n794), .B2(new_n578), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT92), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n775), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n792), .A2(G97), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n310), .B2(new_n772), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT91), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n794), .A2(new_n405), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n777), .A2(new_n273), .B1(new_n784), .B2(new_n221), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n801), .B(new_n802), .C1(G58), .C2(new_n768), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT32), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n787), .B2(G159), .ZN(new_n805));
  INV_X1    g0605(.A(G159), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n786), .A2(KEYINPUT32), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n261), .B1(new_n780), .B2(new_n353), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n805), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n800), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n765), .B1(new_n797), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n700), .A2(new_n393), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G355), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(G116), .B2(new_n209), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n243), .A2(G45), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n700), .A2(new_n374), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n512), .B2(new_n213), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n814), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n761), .A2(new_n764), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n753), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n811), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n755), .A2(new_n758), .B1(new_n763), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  OR2_X1    g0625(.A1(new_n363), .A2(KEYINPUT96), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n363), .A2(KEYINPUT96), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n358), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n673), .A2(new_n691), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n558), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n638), .B1(new_n737), .B2(new_n738), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n647), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n654), .B1(new_n834), .B2(new_n646), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n671), .B1(new_n835), .B2(new_n667), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n683), .B1(new_n836), .B2(new_n656), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n347), .A2(new_n683), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n826), .A2(new_n358), .A3(new_n838), .A4(new_n827), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n632), .A2(new_n683), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n831), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n726), .A2(new_n728), .ZN(new_n843));
  INV_X1    g0643(.A(new_n721), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(G330), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n753), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n846), .B2(new_n842), .ZN(new_n848));
  INV_X1    g0648(.A(new_n772), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G137), .A2(new_n778), .B1(new_n849), .B2(G150), .ZN(new_n850));
  INV_X1    g0650(.A(G143), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n806), .B2(new_n784), .C1(new_n851), .C2(new_n769), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT94), .Z(new_n853));
  AND2_X1   g0653(.A1(new_n853), .A2(KEYINPUT34), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(KEYINPUT34), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n781), .A2(G68), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n273), .B2(new_n794), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT95), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n374), .B1(new_n859), .B2(new_n786), .C1(new_n414), .C2(new_n791), .ZN(new_n860));
  OR4_X1    g0660(.A1(new_n854), .A2(new_n855), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n777), .A2(new_n578), .B1(new_n780), .B2(new_n405), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n261), .B(new_n862), .C1(G311), .C2(new_n787), .ZN(new_n863));
  INV_X1    g0663(.A(new_n794), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G107), .A2(new_n864), .B1(new_n849), .B2(G283), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n768), .A2(G294), .B1(G116), .B2(new_n785), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n863), .A2(new_n798), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n765), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n764), .A2(new_n759), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n754), .B(new_n868), .C1(new_n221), .C2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n841), .B2(new_n760), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n848), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(G384));
  NOR2_X1   g0673(.A1(new_n750), .A2(new_n205), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT40), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT102), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n332), .A2(KEYINPUT99), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT99), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n878), .B(new_n314), .C1(new_n330), .C2(new_n331), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n314), .A2(new_n683), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n335), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n877), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT100), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n330), .A2(new_n331), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n335), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(new_n314), .A3(new_n683), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n882), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n883), .B1(new_n882), .B2(new_n886), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n841), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n876), .B1(new_n729), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n681), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n437), .A2(new_n428), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n428), .A2(new_n410), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n428), .A2(new_n891), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n894), .A3(new_n433), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n893), .A2(new_n894), .A3(new_n897), .A4(new_n433), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n892), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n418), .A2(new_n423), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT16), .B1(new_n902), .B2(new_n379), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n427), .B1(new_n390), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n410), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n433), .A2(new_n905), .A3(KEYINPUT101), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n891), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT101), .B1(new_n433), .B2(new_n905), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n898), .ZN(new_n911));
  INV_X1    g0711(.A(new_n907), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n437), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n901), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n875), .B1(new_n890), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n889), .B1(new_n843), .B2(new_n844), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT38), .ZN(new_n918));
  INV_X1    g0718(.A(new_n898), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n433), .A2(new_n905), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT101), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n906), .A3(new_n907), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n919), .B1(new_n923), .B2(KEYINPUT37), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n437), .A2(new_n912), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n918), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n875), .A3(new_n914), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n876), .A2(KEYINPUT40), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n917), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n916), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT103), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n931), .A2(new_n439), .A3(new_n729), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n931), .B1(new_n439), .B2(new_n729), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(G330), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n828), .A2(new_n683), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n831), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n926), .A2(new_n914), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n887), .A2(new_n888), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT39), .ZN(new_n942));
  AOI221_X4 g0742(.A(new_n918), .B1(new_n437), .B2(new_n912), .C1(new_n910), .C2(new_n898), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n942), .B1(new_n943), .B2(new_n900), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n926), .A2(KEYINPUT39), .A3(new_n914), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n877), .A2(new_n879), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n691), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n944), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n628), .A2(new_n891), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n941), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n733), .A2(new_n440), .A3(new_n746), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n636), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n874), .B1(new_n934), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n934), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n605), .A2(new_n606), .ZN(new_n957));
  INV_X1    g0757(.A(new_n604), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(KEYINPUT35), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(KEYINPUT35), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n960), .A2(G116), .A3(new_n215), .A4(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n415), .A2(new_n212), .A3(new_n221), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n310), .A2(G50), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT98), .Z(new_n967));
  OAI211_X1 g0767(.A(G1), .B(new_n271), .C1(new_n965), .C2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n956), .A2(new_n964), .A3(new_n968), .ZN(G367));
  NOR2_X1   g0769(.A1(new_n739), .A2(new_n691), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n655), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n835), .B2(new_n970), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT104), .Z(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n761), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n768), .A2(G303), .B1(new_n778), .B2(G311), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT111), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n864), .A2(G116), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT46), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n975), .A2(KEYINPUT111), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n780), .A2(new_n530), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G283), .B2(new_n785), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n374), .B1(new_n792), .B2(G107), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G294), .A2(new_n849), .B1(new_n787), .B2(G317), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n778), .A2(G143), .B1(new_n787), .B2(G137), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n273), .B2(new_n784), .C1(new_n279), .C2(new_n769), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n794), .A2(new_n414), .B1(new_n780), .B2(new_n221), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n791), .A2(new_n310), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n261), .B1(new_n772), .B2(new_n806), .ZN(new_n990));
  OR3_X1    g0790(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n980), .A2(new_n985), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT113), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n992), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n764), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n820), .B1(new_n209), .B2(new_n340), .C1(new_n817), .C2(new_n238), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n974), .A2(new_n753), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n683), .B1(new_n612), .B2(new_n615), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n665), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n651), .A2(new_n683), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT105), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT105), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1000), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n696), .A2(new_n1006), .A3(new_n697), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT45), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT44), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1006), .B1(KEYINPUT106), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n698), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1010), .A2(KEYINPUT106), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n694), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1013), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1011), .A2(new_n698), .A3(new_n1016), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1009), .A2(new_n1014), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT110), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n1011), .A2(new_n698), .A3(new_n1016), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1016), .B1(new_n1011), .B2(new_n698), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT110), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1022), .A2(new_n1023), .A3(new_n1015), .A4(new_n1009), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1009), .A2(new_n1014), .A3(new_n1017), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1026), .A2(KEYINPUT107), .A3(new_n694), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n694), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT107), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1025), .A2(new_n1027), .A3(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n692), .B(new_n693), .C1(new_n590), .C2(new_n683), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n689), .A2(KEYINPUT108), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n1032), .A2(new_n696), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1033), .B1(new_n1032), .B2(new_n696), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n733), .A2(new_n746), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n846), .ZN(new_n1039));
  OAI21_X1  g0839(.A(KEYINPUT109), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT109), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n747), .A2(new_n1036), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n747), .B1(new_n1031), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n701), .B(KEYINPUT41), .Z(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n752), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1006), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n616), .B1(new_n1048), .B2(new_n491), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n691), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1006), .A2(new_n501), .A3(new_n695), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(KEYINPUT42), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1051), .A2(KEYINPUT42), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT43), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1053), .A2(new_n1054), .B1(new_n973), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n973), .A2(new_n1055), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1015), .A2(new_n1048), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1058), .B(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n998), .B1(new_n1047), .B2(new_n1060), .ZN(G387));
  OAI21_X1  g0861(.A(new_n701), .B1(new_n747), .B2(new_n1036), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1043), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n692), .A2(new_n693), .A3(new_n761), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n768), .A2(G317), .B1(G303), .B2(new_n785), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G322), .A2(new_n778), .B1(new_n849), .B2(G311), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1068), .A2(KEYINPUT48), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1068), .A2(KEYINPUT48), .ZN(new_n1070));
  INV_X1    g0870(.A(G283), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n791), .A2(new_n1071), .B1(new_n794), .B2(new_n454), .ZN(new_n1072));
  NOR3_X1   g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G116), .A2(new_n781), .B1(new_n787), .B2(G326), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1074), .A2(new_n376), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n769), .A2(new_n273), .B1(new_n794), .B2(new_n221), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n366), .B2(new_n849), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n784), .A2(new_n310), .B1(new_n786), .B2(new_n279), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n981), .B(new_n1080), .C1(G159), .C2(new_n778), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n791), .A2(new_n340), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n376), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n765), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n338), .A2(new_n273), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT50), .Z(new_n1087));
  AOI211_X1 g0887(.A(G45), .B(new_n704), .C1(G68), .C2(G77), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1089), .B(new_n816), .C1(new_n512), .C2(new_n235), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n812), .A2(new_n704), .B1(new_n353), .B2(new_n700), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT114), .Z(new_n1092));
  AOI21_X1  g0892(.A(new_n821), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1085), .A2(new_n754), .A3(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1036), .A2(new_n752), .B1(new_n1065), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1064), .A2(KEYINPUT115), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT115), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1062), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1095), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1096), .A2(new_n1100), .ZN(G393));
  NAND3_X1  g0901(.A1(new_n1025), .A2(new_n752), .A3(new_n1028), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n816), .A2(new_n246), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n821), .B1(G97), .B2(new_n700), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n754), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n219), .A2(new_n864), .B1(new_n781), .B2(G87), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1106), .B(new_n374), .C1(new_n851), .C2(new_n786), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT116), .Z(new_n1108));
  NAND2_X1  g0908(.A1(new_n338), .A2(new_n785), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n791), .A2(new_n221), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G50), .B2(new_n849), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n768), .A2(G159), .B1(new_n778), .B2(G150), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT51), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1109), .B(new_n1111), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n768), .A2(G311), .B1(new_n778), .B2(G317), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT52), .Z(new_n1119));
  OAI221_X1 g0919(.A(new_n393), .B1(new_n780), .B2(new_n353), .C1(new_n791), .C2(new_n565), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n1071), .A2(new_n794), .B1(new_n784), .B2(new_n454), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n772), .A2(new_n578), .B1(new_n786), .B2(new_n770), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1108), .A2(new_n1117), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1105), .B1(new_n765), .B2(new_n1124), .C1(new_n1006), .C2(new_n762), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n701), .B1(new_n1031), .B2(new_n1043), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1127), .A2(new_n1043), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1102), .B(new_n1125), .C1(new_n1126), .C2(new_n1128), .ZN(G390));
  AOI211_X1 g0929(.A(new_n683), .B(new_n829), .C1(new_n742), .C2(new_n744), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT117), .B1(new_n1130), .B2(new_n935), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n745), .A2(new_n691), .A3(new_n830), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT117), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n936), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n940), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n948), .B1(new_n901), .B2(new_n914), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n935), .B1(new_n837), .B2(new_n830), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n947), .B1(new_n1138), .B2(new_n939), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n944), .A2(new_n945), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n841), .ZN(new_n1143));
  NOR4_X1   g0943(.A1(new_n729), .A2(new_n939), .A3(new_n730), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n731), .A2(new_n841), .A3(new_n940), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1137), .A2(new_n1141), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n939), .B1(new_n846), .B2(new_n1143), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1134), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1133), .B1(new_n1132), .B2(new_n936), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1149), .B(new_n1146), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n940), .B1(new_n731), .B2(new_n841), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n937), .B1(new_n1153), .B2(new_n1144), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n952), .B(new_n636), .C1(new_n439), .C2(new_n846), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1148), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1156), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1145), .A2(new_n1147), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1161), .A3(new_n701), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1145), .A2(new_n752), .A3(new_n1147), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT119), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1140), .A2(new_n759), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n754), .B1(new_n277), .B2(new_n869), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n856), .B1(new_n454), .B2(new_n786), .C1(new_n769), .C2(new_n565), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1167), .A2(new_n261), .A3(new_n801), .A4(new_n1110), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n777), .A2(new_n1071), .B1(new_n772), .B2(new_n353), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G97), .B2(new_n785), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT118), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n261), .B1(new_n780), .B2(new_n273), .ZN(new_n1172));
  INV_X1    g0972(.A(G128), .ZN(new_n1173));
  INV_X1    g0973(.A(G125), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n777), .A2(new_n1173), .B1(new_n786), .B2(new_n1174), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1172), .B(new_n1175), .C1(G159), .C2(new_n792), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n864), .A2(G150), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT53), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT54), .B(G143), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n784), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n849), .A2(G137), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n769), .B2(new_n859), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1178), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1168), .A2(new_n1171), .B1(new_n1176), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1165), .B(new_n1166), .C1(new_n765), .C2(new_n1184), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1163), .A2(new_n1164), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1164), .B1(new_n1163), .B2(new_n1185), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1162), .B1(new_n1186), .B2(new_n1187), .ZN(G378));
  AOI21_X1  g0988(.A(new_n754), .B1(new_n273), .B2(new_n869), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n769), .A2(new_n1173), .B1(new_n772), .B2(new_n859), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G125), .A2(new_n778), .B1(new_n785), .B2(G137), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n794), .B2(new_n1179), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(G150), .C2(new_n792), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT59), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n253), .B(new_n254), .C1(new_n780), .C2(new_n806), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G124), .B2(new_n787), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n780), .A2(new_n414), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G283), .B2(new_n787), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n221), .B2(new_n794), .C1(new_n353), .C2(new_n769), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G116), .A2(new_n778), .B1(new_n849), .B2(G97), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n340), .B2(new_n784), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n376), .A2(new_n254), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1202), .A2(new_n1204), .A3(new_n989), .A4(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1205), .B(new_n273), .C1(G33), .C2(G41), .ZN(new_n1209));
  AND4_X1   g1009(.A1(new_n1199), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n292), .A2(new_n891), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n301), .B(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1212), .B(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1189), .B1(new_n765), .B2(new_n1210), .C1(new_n1214), .C2(new_n760), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT120), .ZN(new_n1216));
  OAI21_X1  g1016(.A(G330), .B1(new_n916), .B2(new_n929), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n941), .A2(new_n949), .A3(new_n950), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n951), .B(G330), .C1(new_n916), .C2(new_n929), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1214), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1214), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1219), .A2(new_n1220), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1216), .B1(new_n1225), .B2(new_n752), .ZN(new_n1226));
  AOI221_X4 g1026(.A(new_n1144), .B1(new_n1139), .B2(new_n1140), .C1(new_n1135), .C2(new_n1136), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1146), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1156), .B1(new_n1229), .B2(new_n1155), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1219), .A2(new_n1220), .A3(new_n1223), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1223), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n701), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1161), .A2(new_n1157), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT57), .B1(new_n1235), .B2(new_n1225), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1226), .B1(new_n1234), .B2(new_n1236), .ZN(G375));
  NAND2_X1  g1037(.A1(new_n1155), .A2(new_n752), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT122), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT122), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1155), .A2(new_n1240), .A3(new_n752), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n754), .B1(new_n310), .B2(new_n869), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n786), .A2(new_n1173), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n806), .A2(new_n794), .B1(new_n772), .B2(new_n1179), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(G137), .C2(new_n768), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n778), .A2(KEYINPUT124), .A3(G132), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT124), .B1(new_n778), .B2(G132), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G50), .B2(new_n792), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n376), .B(new_n1200), .C1(G150), .C2(new_n785), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1245), .A2(new_n1246), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n393), .B1(new_n780), .B2(new_n221), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n1251), .B(KEYINPUT123), .Z(new_n1252));
  AOI22_X1  g1052(.A1(new_n768), .A2(G283), .B1(G97), .B2(new_n864), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n778), .A2(G294), .B1(new_n787), .B2(G303), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n353), .A2(new_n784), .B1(new_n772), .B2(new_n565), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1255), .A2(new_n1082), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .A4(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1250), .A2(new_n1257), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1242), .B1(new_n765), .B2(new_n1258), .C1(new_n940), .C2(new_n760), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1239), .A2(new_n1241), .A3(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1152), .A2(new_n1156), .A3(new_n1154), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1045), .B(KEYINPUT121), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1158), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(G381));
  NOR2_X1   g1065(.A1(G393), .A2(G396), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NOR4_X1   g1067(.A1(new_n1267), .A2(G381), .A3(G384), .A4(G390), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1225), .A2(new_n752), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1216), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1235), .A2(new_n1225), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT57), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1273), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n702), .B1(new_n1275), .B2(new_n1235), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1271), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(G387), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1163), .A2(new_n1185), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n702), .B1(new_n1148), .B2(new_n1158), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1280), .B2(new_n1161), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1268), .A2(new_n1277), .A3(new_n1278), .A4(new_n1281), .ZN(G407));
  INV_X1    g1082(.A(G213), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(G343), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1277), .A2(new_n1281), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(G407), .A2(G213), .A3(new_n1285), .ZN(G409));
  INV_X1    g1086(.A(G390), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G387), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n824), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1266), .A2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G390), .B(new_n998), .C1(new_n1047), .C2(new_n1060), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1290), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1290), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT127), .B1(new_n1299), .B2(new_n1292), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1235), .A2(new_n1225), .A3(new_n1263), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1226), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1281), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1187), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1163), .A2(new_n1164), .A3(new_n1185), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n1305), .A2(new_n1306), .B1(new_n1161), .B2(new_n1280), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1304), .B1(G375), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1284), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1262), .A2(KEYINPUT125), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT60), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1262), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1158), .A2(new_n701), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(G384), .A3(new_n1261), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1315), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n872), .B1(new_n1319), .B2(new_n1260), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1308), .A2(new_n1309), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT126), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1308), .A2(KEYINPUT126), .A3(new_n1309), .A4(new_n1322), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT62), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1284), .A2(G2897), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1318), .A2(new_n1320), .A3(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AOI22_X1  g1131(.A1(new_n1277), .A2(G378), .B1(new_n1281), .B2(new_n1303), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1331), .B1(new_n1332), .B2(new_n1284), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT61), .ZN(new_n1334));
  OAI211_X1 g1134(.A(G378), .B(new_n1226), .C1(new_n1236), .C2(new_n1234), .ZN(new_n1335));
  AOI211_X1 g1135(.A(new_n1284), .B(new_n1321), .C1(new_n1335), .C2(new_n1304), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT62), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1333), .B(new_n1334), .C1(new_n1336), .C2(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1301), .B1(new_n1327), .B2(new_n1338), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1340));
  AND3_X1   g1140(.A1(new_n1333), .A2(new_n1334), .A3(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT63), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1325), .A2(new_n1342), .A3(new_n1326), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1336), .A2(KEYINPUT63), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1341), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1339), .A2(new_n1345), .ZN(G405));
  NAND2_X1  g1146(.A1(G375), .A2(new_n1281), .ZN(new_n1347));
  AND2_X1   g1147(.A1(new_n1347), .A2(new_n1335), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1348), .A2(new_n1321), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1348), .A2(new_n1321), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1301), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1351), .ZN(new_n1353));
  OAI22_X1  g1153(.A1(new_n1353), .A2(new_n1349), .B1(new_n1296), .B2(new_n1300), .ZN(new_n1354));
  AND2_X1   g1154(.A1(new_n1352), .A2(new_n1354), .ZN(G402));
endmodule


