//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XOR2_X1   g0002(.A(new_n202), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT65), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  INV_X1    g0007(.A(G226), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n205), .B1(new_n211), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n205), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n219), .B(new_n222), .C1(new_n225), .C2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT66), .ZN(G361));
  XOR2_X1   g0029(.A(G250), .B(G257), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT67), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n213), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G58), .A2(G68), .ZN(new_n249));
  OAI21_X1  g0049(.A(G20), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G159), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(KEYINPUT16), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT7), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n255), .B(new_n224), .C1(new_n259), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G68), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT76), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G33), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(G20), .B1(new_n268), .B2(new_n260), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(new_n255), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n254), .B1(new_n263), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT77), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n247), .B1(new_n269), .B2(new_n255), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n256), .A2(new_n257), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n261), .B1(new_n274), .B2(G33), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT7), .B1(new_n275), .B2(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT77), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(new_n254), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n223), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n250), .A2(new_n252), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n265), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n260), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT7), .B1(new_n287), .B2(new_n224), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT78), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n256), .A2(new_n257), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n266), .A2(new_n258), .A3(new_n267), .ZN(new_n294));
  INV_X1    g0094(.A(new_n292), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT78), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n288), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n285), .B1(new_n297), .B2(new_n247), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT16), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n283), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n280), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G13), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n302), .A2(new_n224), .A3(G1), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n282), .ZN(new_n304));
  INV_X1    g0104(.A(G1), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G20), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT8), .B(G58), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n302), .A2(G1), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G20), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n309), .B1(new_n311), .B2(new_n308), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT79), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G223), .A2(G1698), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n208), .B2(G1698), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n317), .A2(new_n268), .A3(new_n260), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G87), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT80), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n318), .A2(KEYINPUT80), .A3(new_n319), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G190), .ZN(new_n326));
  INV_X1    g0126(.A(G41), .ZN(new_n327));
  OAI211_X1 g0127(.A(G1), .B(G13), .C1(new_n258), .C2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G45), .ZN(new_n329));
  AOI21_X1  g0129(.A(G1), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(G274), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n330), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n328), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n331), .B1(new_n333), .B2(new_n214), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n325), .A2(new_n326), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n328), .B1(new_n320), .B2(new_n321), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n334), .B1(new_n337), .B2(new_n324), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n336), .B1(G200), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n301), .A2(new_n315), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT17), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n314), .B1(new_n280), .B2(new_n300), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  AOI211_X1 g0144(.A(new_n344), .B(new_n334), .C1(new_n337), .C2(new_n324), .ZN(new_n345));
  INV_X1    g0145(.A(G169), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n325), .B2(new_n335), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT18), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n278), .B1(new_n277), .B2(new_n254), .ZN(new_n350));
  AOI211_X1 g0150(.A(KEYINPUT77), .B(new_n253), .C1(new_n273), .C2(new_n276), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n288), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n290), .A2(new_n289), .A3(new_n292), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT78), .B1(new_n294), .B2(new_n295), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n284), .B1(new_n356), .B2(G68), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n282), .B1(new_n357), .B2(KEYINPUT16), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n315), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT18), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n338), .A2(G179), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n346), .B2(new_n338), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n343), .A2(KEYINPUT17), .A3(new_n339), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n342), .A2(new_n349), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n365), .A2(KEYINPUT81), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n260), .A2(new_n286), .ZN(new_n367));
  INV_X1    g0167(.A(G1698), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(G232), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(G238), .A3(G1698), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n287), .A2(G107), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n323), .ZN(new_n373));
  INV_X1    g0173(.A(new_n331), .ZN(new_n374));
  INV_X1    g0174(.A(new_n333), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(G244), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n346), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G20), .A2(G77), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT15), .B(G87), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n224), .A2(G33), .ZN(new_n381));
  INV_X1    g0181(.A(new_n251), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n379), .B1(new_n380), .B2(new_n381), .C1(new_n382), .C2(new_n307), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n311), .A2(KEYINPUT70), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT70), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n303), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G77), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n282), .A2(new_n383), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n282), .B1(new_n384), .B2(new_n386), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n388), .B1(new_n305), .B2(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(KEYINPUT71), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT71), .B1(new_n390), .B2(new_n391), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n378), .B(new_n395), .C1(G179), .C2(new_n377), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n377), .A2(G200), .ZN(new_n397));
  INV_X1    g0197(.A(new_n394), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n392), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n373), .A2(G190), .A3(new_n376), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n397), .A2(new_n399), .A3(new_n389), .A4(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT72), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT10), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n403), .A2(KEYINPUT10), .ZN(new_n405));
  INV_X1    g0205(.A(G150), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n307), .A2(new_n381), .B1(new_n406), .B2(new_n382), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n224), .B1(new_n249), .B2(new_n207), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n282), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n207), .B1(new_n305), .B2(G20), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n304), .A2(new_n410), .B1(new_n207), .B2(new_n303), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT9), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT9), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n409), .A2(new_n414), .A3(new_n411), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n367), .A2(G222), .A3(new_n368), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n367), .A2(G223), .A3(G1698), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n287), .A2(G77), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n323), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n331), .B1(new_n333), .B2(new_n208), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT69), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n331), .B(KEYINPUT69), .C1(new_n333), .C2(new_n208), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n416), .B1(new_n326), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(G200), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n404), .B(new_n405), .C1(new_n427), .C2(new_n429), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n431), .A2(G190), .B1(new_n413), .B2(new_n415), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n432), .A2(new_n403), .A3(KEYINPUT10), .A4(new_n428), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n344), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n426), .A2(new_n346), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n412), .A3(new_n435), .ZN(new_n436));
  AND4_X1   g0236(.A1(new_n402), .A2(new_n430), .A3(new_n433), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n247), .A2(G20), .ZN(new_n438));
  OAI221_X1 g0238(.A(new_n438), .B1(new_n381), .B2(new_n388), .C1(new_n382), .C2(new_n207), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n282), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT11), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n390), .A2(G68), .A3(new_n306), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n387), .A2(new_n247), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n438), .A2(KEYINPUT12), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n444), .A2(new_n445), .B1(new_n310), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n374), .B1(new_n375), .B2(G238), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n260), .A2(new_n286), .A3(G226), .A4(new_n368), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n260), .A2(new_n286), .A3(G232), .A4(G1698), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G97), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n454), .A2(KEYINPUT73), .A3(new_n323), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT73), .B1(new_n454), .B2(new_n323), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n450), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT13), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT13), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n450), .B(new_n459), .C1(new_n455), .C2(new_n456), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT14), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n462), .A3(G169), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n344), .B2(new_n461), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n461), .B2(G169), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n449), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(G200), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT74), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n461), .A2(KEYINPUT74), .A3(G200), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n448), .B1(new_n461), .B2(new_n326), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n437), .A2(new_n466), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n365), .A2(KEYINPUT81), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n366), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n328), .A2(G274), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n329), .A2(G1), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(new_n210), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n479), .A2(new_n480), .B1(new_n328), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT85), .ZN(new_n483));
  OR2_X1    g0283(.A1(KEYINPUT84), .A2(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(KEYINPUT84), .A2(G116), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n258), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(G238), .A2(G1698), .ZN(new_n487));
  INV_X1    g0287(.A(G244), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(G1698), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n486), .B1(new_n275), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n482), .B(new_n483), .C1(new_n490), .C2(new_n328), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n268), .A3(new_n260), .ZN(new_n492));
  INV_X1    g0292(.A(new_n486), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n328), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n481), .A2(new_n328), .ZN(new_n495));
  INV_X1    g0295(.A(new_n480), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n478), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT85), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n491), .A2(new_n498), .A3(G200), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n268), .A2(new_n224), .A3(G68), .A4(new_n260), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT19), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n224), .B1(new_n453), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(G97), .A2(G107), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n209), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n224), .A2(G33), .A3(G97), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n502), .A2(new_n504), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n282), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n387), .A2(new_n380), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n304), .B1(G1), .B2(new_n258), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n510), .B1(G87), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n491), .A2(new_n498), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT87), .B1(new_n514), .B2(G190), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT87), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n516), .B(new_n326), .C1(new_n491), .C2(new_n498), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n499), .B(new_n513), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n508), .B(new_n509), .C1(new_n380), .C2(new_n511), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n519), .A2(KEYINPUT86), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n514), .A2(new_n344), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n491), .A2(new_n498), .A3(new_n346), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(KEYINPUT86), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(G250), .A2(G1698), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n216), .B2(G1698), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(new_n268), .A3(new_n260), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G294), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n328), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g0330(.A(KEYINPUT5), .B(G41), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n480), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n532), .A2(G264), .A3(new_n328), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n531), .A2(new_n328), .A3(G274), .A4(new_n480), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n530), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n536), .A2(G179), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n346), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT23), .B1(new_n224), .B2(G107), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  INV_X1    g0340(.A(G107), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(G20), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n486), .B2(new_n224), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n209), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n268), .A2(new_n224), .A3(new_n260), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n224), .A2(G87), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n545), .B1(new_n287), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n544), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT24), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT24), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n544), .A2(new_n552), .A3(new_n547), .A4(new_n549), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n283), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n303), .A2(new_n541), .ZN(new_n555));
  XOR2_X1   g0355(.A(new_n555), .B(KEYINPUT25), .Z(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n541), .B2(new_n511), .ZN(new_n557));
  OAI22_X1  g0357(.A1(new_n537), .A2(new_n538), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n554), .A2(new_n557), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n530), .A2(new_n533), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n326), .A3(new_n534), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G200), .B2(new_n536), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT89), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n560), .A2(new_n563), .A3(KEYINPUT89), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n559), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n511), .A2(new_n215), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n311), .A2(G97), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n541), .A2(KEYINPUT6), .A3(G97), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n215), .A2(new_n541), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n503), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n573), .B2(KEYINPUT6), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(G20), .B1(G77), .B2(new_n251), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n297), .B2(new_n541), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n569), .B(new_n570), .C1(new_n576), .C2(new_n282), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n532), .A2(G257), .A3(new_n328), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n534), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT83), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(KEYINPUT83), .A3(new_n534), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT4), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n268), .A2(new_n260), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n488), .A2(G1698), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n584), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(KEYINPUT4), .A2(G244), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n260), .A2(new_n286), .A3(new_n589), .A4(new_n368), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n260), .A2(new_n286), .A3(G250), .A4(G1698), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G283), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n328), .B1(new_n588), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n583), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G190), .ZN(new_n597));
  INV_X1    g0397(.A(G200), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT4), .B1(new_n275), .B2(new_n586), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n323), .B1(new_n599), .B2(new_n593), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT82), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n595), .A2(KEYINPUT82), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n583), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n577), .B(new_n597), .C1(new_n598), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n576), .A2(new_n282), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n569), .A2(new_n570), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n600), .A2(new_n581), .A3(new_n582), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n606), .A2(new_n607), .B1(new_n608), .B2(new_n346), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n581), .A2(new_n582), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n595), .A2(KEYINPUT82), .ZN(new_n611));
  AOI211_X1 g0411(.A(new_n601), .B(new_n328), .C1(new_n588), .C2(new_n594), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n610), .B(new_n344), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n605), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n532), .A2(G270), .A3(new_n328), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n616), .B(KEYINPUT88), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n216), .A2(new_n368), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(G264), .B2(new_n368), .ZN(new_n619));
  INV_X1    g0419(.A(G303), .ZN(new_n620));
  OAI22_X1  g0420(.A1(new_n585), .A2(new_n619), .B1(new_n620), .B2(new_n367), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n535), .B1(new_n621), .B2(new_n323), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G200), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n484), .A2(new_n485), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G116), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n305), .B2(G33), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n387), .A2(new_n626), .B1(new_n390), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n592), .B(new_n224), .C1(G33), .C2(new_n215), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n282), .B(new_n630), .C1(new_n625), .C2(new_n224), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT20), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n624), .B(new_n635), .C1(new_n326), .C2(new_n623), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n623), .A2(new_n634), .A3(G169), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n617), .A2(G179), .A3(new_n622), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n634), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n623), .A2(new_n634), .A3(KEYINPUT21), .A4(G169), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n636), .A2(new_n639), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n615), .A2(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n477), .A2(new_n525), .A3(new_n568), .A4(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n436), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n396), .A2(KEYINPUT92), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n396), .A2(KEYINPUT92), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n465), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n650), .B(new_n463), .C1(new_n344), .C2(new_n461), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n474), .A2(new_n649), .B1(new_n651), .B2(new_n449), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n342), .A2(new_n364), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n349), .B(new_n363), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n430), .A2(new_n433), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n646), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT90), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n494), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n482), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n346), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n519), .A3(new_n521), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT91), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n566), .A2(new_n567), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n606), .A2(new_n607), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n608), .A2(new_n326), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G200), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n667), .A2(new_n669), .B1(new_n613), .B2(new_n609), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n639), .A2(new_n558), .A3(new_n641), .A4(new_n642), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n664), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n659), .A2(G200), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n673), .B(new_n513), .C1(new_n515), .C2(new_n517), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n661), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n663), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n675), .B2(new_n614), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n608), .A2(new_n346), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n613), .A2(new_n665), .A3(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n518), .A2(new_n681), .A3(KEYINPUT26), .A4(new_n524), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n477), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n656), .A2(new_n685), .ZN(G369));
  AND3_X1   g0486(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n310), .A2(new_n224), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n310), .A2(new_n691), .A3(new_n224), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT93), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n635), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n688), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n643), .B2(new_n699), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G330), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n558), .A2(new_n698), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT94), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n560), .A2(new_n698), .ZN(new_n708));
  AOI211_X1 g0508(.A(new_n708), .B(new_n559), .C1(new_n566), .C2(new_n567), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n688), .A2(new_n698), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n698), .B(KEYINPUT95), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n558), .ZN(new_n717));
  OR3_X1    g0517(.A1(new_n713), .A2(new_n715), .A3(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n220), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n504), .A2(G116), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n720), .A2(new_n305), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n227), .B2(new_n720), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT28), .Z(new_n725));
  NAND3_X1  g0525(.A1(new_n518), .A2(new_n681), .A3(new_n524), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n678), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n674), .A2(new_n681), .A3(KEYINPUT26), .A4(new_n661), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n661), .B(KEYINPUT91), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n664), .A2(new_n670), .A3(new_n671), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n730), .B1(new_n731), .B2(new_n675), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT29), .B(new_n698), .C1(new_n729), .C2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n716), .B1(new_n677), .B2(new_n683), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(KEYINPUT29), .ZN(new_n735));
  INV_X1    g0535(.A(new_n716), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n644), .A2(new_n525), .A3(new_n568), .A4(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT96), .B1(new_n604), .B2(new_n536), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT96), .ZN(new_n740));
  INV_X1    g0540(.A(new_n536), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n668), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n659), .A2(new_n344), .A3(new_n623), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n640), .A2(new_n596), .A3(new_n514), .A4(new_n561), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT30), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n608), .A2(new_n533), .A3(new_n530), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT30), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(new_n749), .A3(new_n514), .A4(new_n640), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n743), .A2(new_n745), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n738), .B1(new_n751), .B2(new_n698), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n747), .A2(new_n750), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n744), .B1(new_n739), .B2(new_n742), .ZN(new_n754));
  OAI211_X1 g0554(.A(KEYINPUT31), .B(new_n716), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n737), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n735), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n725), .B1(new_n759), .B2(G1), .ZN(G364));
  NAND2_X1  g0560(.A1(new_n702), .A2(new_n703), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT97), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n302), .A2(G20), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT98), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G45), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G1), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n720), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n762), .B(new_n768), .C1(new_n703), .C2(new_n702), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n223), .B1(G20), .B2(new_n346), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n224), .A2(new_n344), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n224), .A2(G179), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(G190), .A3(G200), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n775), .A2(new_n247), .B1(new_n209), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n773), .A2(new_n326), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G190), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G159), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n780), .A2(new_n207), .B1(new_n784), .B2(KEYINPUT32), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n778), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n776), .A2(new_n326), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT99), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G107), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n772), .A2(G190), .A3(new_n598), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n367), .B1(new_n794), .B2(new_n213), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n772), .A2(new_n781), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n795), .B1(G77), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n344), .A2(new_n598), .A3(G190), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n215), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(KEYINPUT32), .B2(new_n784), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n786), .A2(new_n793), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n792), .A2(G283), .ZN(new_n805));
  INV_X1    g0605(.A(new_n794), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n806), .A2(G322), .B1(new_n783), .B2(G329), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n367), .B1(new_n797), .B2(G311), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT33), .B(G317), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n774), .A2(new_n810), .B1(G294), .B2(new_n800), .ZN(new_n811));
  INV_X1    g0611(.A(new_n777), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n779), .A2(G326), .B1(new_n812), .B2(G303), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n805), .A2(new_n809), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n771), .B1(new_n804), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G13), .A2(G33), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G20), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n770), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n220), .A2(G355), .A3(new_n367), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n719), .A2(new_n275), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(G45), .B2(new_n226), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n245), .A2(new_n329), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n820), .B1(G116), .B2(new_n220), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n768), .B(new_n815), .C1(new_n819), .C2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT100), .ZN(new_n826));
  INV_X1    g0626(.A(new_n818), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n701), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n769), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  NAND2_X1  g0630(.A1(new_n771), .A2(new_n817), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n767), .B1(G77), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G294), .ZN(new_n833));
  INV_X1    g0633(.A(G311), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n794), .A2(new_n833), .B1(new_n782), .B2(new_n834), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n367), .B(new_n835), .C1(new_n625), .C2(new_n797), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n792), .A2(G87), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n802), .B1(G107), .B2(new_n812), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n774), .A2(G283), .B1(new_n779), .B2(G303), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n806), .A2(G143), .B1(new_n797), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n775), .B2(new_n406), .C1(new_n842), .C2(new_n780), .ZN(new_n843));
  XNOR2_X1  g0643(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n801), .A2(new_n213), .B1(new_n207), .B2(new_n777), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n585), .B(new_n846), .C1(G132), .C2(new_n783), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n845), .B(new_n847), .C1(new_n247), .C2(new_n791), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n843), .A2(new_n844), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n840), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n832), .B1(new_n850), .B2(new_n770), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n695), .A2(new_n696), .ZN(new_n852));
  INV_X1    g0652(.A(G343), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n647), .A2(new_n395), .A3(new_n648), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n395), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n396), .A2(new_n401), .A3(new_n856), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n857), .A2(KEYINPUT102), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(KEYINPUT102), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n851), .B1(new_n860), .B2(new_n817), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT103), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n734), .B(new_n860), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n864), .A2(new_n757), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n864), .A2(new_n757), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT104), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n865), .B(new_n768), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n863), .B1(new_n868), .B2(new_n870), .ZN(G384));
  NOR2_X1   g0671(.A1(new_n764), .A2(new_n305), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n396), .A2(new_n854), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n734), .B2(new_n860), .ZN(new_n874));
  INV_X1    g0674(.A(new_n339), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n285), .B1(new_n263), .B2(new_n270), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n283), .B1(new_n876), .B2(new_n299), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n314), .B1(new_n280), .B2(new_n877), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n359), .A2(new_n875), .B1(new_n878), .B2(new_n852), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n348), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n359), .A2(new_n362), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n697), .B(KEYINPUT105), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n359), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n882), .A2(new_n884), .A3(new_n885), .A4(new_n340), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n878), .A2(new_n852), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n365), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n887), .B2(new_n889), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n472), .B1(new_n469), .B2(new_n470), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n449), .B(new_n854), .C1(new_n651), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n449), .A2(new_n854), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n466), .A2(new_n474), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n874), .A2(new_n893), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n883), .B1(new_n349), .B2(new_n363), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n891), .A2(new_n892), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT107), .ZN(new_n905));
  AND4_X1   g0705(.A1(new_n905), .A2(new_n887), .A3(KEYINPUT38), .A4(new_n889), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n881), .A2(new_n886), .B1(new_n365), .B2(new_n888), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT38), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT106), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n885), .B1(new_n884), .B2(new_n910), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n911), .A2(new_n882), .A3(new_n340), .A4(new_n884), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n852), .B(KEYINPUT105), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n343), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT37), .B1(new_n914), .B2(KEYINPUT106), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n882), .A2(new_n884), .A3(new_n340), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n365), .A2(new_n914), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n909), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n906), .B1(new_n908), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n904), .B1(new_n921), .B2(new_n903), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n651), .A2(new_n449), .A3(new_n698), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n902), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n477), .B(new_n733), .C1(new_n734), .C2(KEYINPUT29), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n656), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n926), .B(new_n928), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n895), .B2(new_n897), .ZN(new_n931));
  OAI211_X1 g0731(.A(KEYINPUT31), .B(new_n854), .C1(new_n753), .C2(new_n754), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n737), .A2(new_n752), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n931), .A2(KEYINPUT40), .A3(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n933), .B(new_n931), .C1(new_n891), .C2(new_n892), .ZN(new_n935));
  XNOR2_X1  g0735(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n921), .A2(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n477), .A3(new_n933), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n921), .A2(new_n934), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n935), .A2(new_n936), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n477), .A2(new_n933), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n938), .A2(new_n943), .A3(G330), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n872), .B1(new_n929), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n929), .B2(new_n944), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n574), .A2(KEYINPUT35), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n574), .A2(KEYINPUT35), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n947), .A2(G116), .A3(new_n225), .A4(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT36), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n248), .A2(new_n226), .A3(new_n388), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n247), .A2(G50), .ZN(new_n952));
  OAI211_X1 g0752(.A(G1), .B(new_n302), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n946), .A2(new_n950), .A3(new_n953), .ZN(G367));
  NAND2_X1  g0754(.A1(new_n716), .A2(new_n681), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT110), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n670), .B1(new_n736), .B2(new_n577), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n559), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n716), .B1(new_n959), .B2(new_n614), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n698), .A2(new_n513), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n676), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n730), .B2(new_n961), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n715), .A2(new_n958), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT111), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT42), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT111), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n967), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT42), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n960), .B(new_n966), .C1(new_n970), .C2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n956), .A2(new_n957), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n712), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n960), .B1(new_n970), .B2(new_n973), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT43), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n966), .B1(new_n979), .B2(new_n964), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n975), .B(new_n977), .C1(new_n978), .C2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n978), .A2(new_n980), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n982), .A2(new_n974), .B1(new_n712), .B2(new_n976), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n720), .B(KEYINPUT41), .Z(new_n984));
  OAI21_X1  g0784(.A(new_n976), .B1(new_n715), .B2(new_n717), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT44), .Z(new_n986));
  NOR3_X1   g0786(.A1(new_n976), .A2(new_n715), .A3(new_n717), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n713), .ZN(new_n990));
  INV_X1    g0790(.A(new_n714), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n710), .B(new_n991), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(new_n704), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n704), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n758), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n986), .A2(new_n988), .A3(new_n712), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n990), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n984), .B1(new_n998), .B2(new_n759), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n981), .B(new_n983), .C1(new_n999), .C2(new_n766), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n821), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n819), .B1(new_n220), .B2(new_n380), .C1(new_n233), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT112), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n768), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n1003), .B2(new_n1002), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n367), .B1(new_n796), .B2(new_n207), .C1(new_n406), .C2(new_n794), .ZN(new_n1006));
  INV_X1    g0806(.A(G143), .ZN(new_n1007));
  INV_X1    g0807(.A(G159), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n1007), .A2(new_n780), .B1(new_n775), .B2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1006), .B(new_n1009), .C1(G68), .C2(new_n800), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n791), .A2(new_n388), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n777), .A2(new_n213), .B1(new_n782), .B2(new_n842), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1011), .B1(KEYINPUT114), .B2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1010), .B(new_n1013), .C1(KEYINPUT114), .C2(new_n1012), .ZN(new_n1014));
  INV_X1    g0814(.A(G283), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n794), .A2(new_n620), .B1(new_n796), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n585), .B1(new_n780), .B2(new_n834), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(G317), .C2(new_n783), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n626), .B2(new_n777), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n792), .A2(G97), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(KEYINPUT46), .A2(G116), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n775), .A2(new_n833), .B1(new_n777), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G107), .B2(new_n800), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1014), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT47), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1005), .B1(new_n1027), .B2(new_n770), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n963), .B2(new_n827), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1000), .A2(new_n1029), .ZN(G387));
  INV_X1    g0830(.A(new_n995), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n710), .A2(new_n818), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n806), .A2(G317), .B1(new_n797), .B2(G303), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT116), .B(G322), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1033), .B1(new_n775), .B2(new_n834), .C1(new_n780), .C2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n812), .A2(G294), .B1(new_n800), .B2(G283), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT49), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n791), .A2(new_n626), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n275), .B(new_n1044), .C1(G326), .C2(new_n783), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1008), .A2(new_n780), .B1(new_n775), .B2(new_n307), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n777), .A2(new_n388), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n797), .A2(G68), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(KEYINPUT115), .B(G150), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1050), .B1(new_n207), .B2(new_n794), .C1(new_n782), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n380), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n585), .B1(new_n1054), .B2(new_n800), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1049), .A2(new_n1021), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n771), .B1(new_n1046), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n821), .B1(new_n237), .B2(new_n329), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n220), .A2(new_n367), .A3(new_n722), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n307), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1061));
  OAI21_X1  g0861(.A(KEYINPUT50), .B1(new_n307), .B2(G50), .ZN(new_n1062));
  AOI21_X1  g0862(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n721), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1060), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(G107), .B2(new_n220), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n768), .B(new_n1057), .C1(new_n819), .C2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1031), .A2(new_n766), .B1(new_n1032), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n996), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n720), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1031), .A2(new_n759), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(G393));
  NOR2_X1   g0872(.A1(new_n242), .A2(new_n1001), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n819), .B1(new_n220), .B2(new_n215), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n767), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n775), .A2(new_n207), .B1(new_n247), .B2(new_n777), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G77), .B2(new_n800), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n308), .A2(new_n797), .B1(new_n783), .B2(G143), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1077), .A2(new_n275), .A3(new_n837), .A4(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G150), .A2(new_n779), .B1(new_n806), .B2(G159), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT51), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n775), .A2(new_n620), .B1(new_n1015), .B2(new_n777), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n625), .B2(new_n800), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n287), .B1(new_n782), .B2(new_n1034), .C1(new_n833), .C2(new_n796), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n793), .A3(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G317), .A2(new_n779), .B1(new_n806), .B2(G311), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT52), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1079), .A2(new_n1081), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1075), .B1(new_n1089), .B2(new_n770), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n958), .B2(new_n827), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n990), .A2(new_n997), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n766), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n998), .A2(new_n720), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1069), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(G390));
  OAI211_X1 g0898(.A(new_n698), .B(new_n860), .C1(new_n729), .C2(new_n732), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n873), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n898), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n923), .A3(new_n921), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n756), .A2(new_n898), .A3(G330), .A4(new_n860), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n683), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n736), .B(new_n860), .C1(new_n1105), .C2(new_n732), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n1100), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n924), .B1(new_n1107), .B2(new_n898), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1103), .B(new_n1104), .C1(new_n922), .C2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n907), .A2(new_n905), .A3(KEYINPUT38), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n911), .B(new_n916), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n365), .A2(new_n914), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT38), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n890), .A2(KEYINPUT107), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n903), .B(new_n1110), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n893), .A2(KEYINPUT39), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n923), .B1(new_n874), .B2(new_n899), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n923), .B(new_n1110), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1117), .A2(new_n1118), .B1(new_n1120), .B2(new_n1102), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n933), .A2(G330), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n931), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1109), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1124), .A2(new_n1093), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1117), .A2(new_n816), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n367), .B1(new_n783), .B2(G294), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n215), .B2(new_n796), .C1(new_n627), .C2(new_n794), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n812), .A2(G87), .B1(new_n800), .B2(G77), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n775), .B2(new_n541), .C1(new_n1015), .C2(new_n780), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(G68), .C2(new_n792), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n774), .A2(G137), .B1(G159), .B2(new_n800), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n780), .C1(new_n791), .C2(new_n207), .ZN(new_n1134));
  NOR3_X1   g0934(.A1(new_n777), .A2(new_n1051), .A3(KEYINPUT53), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n806), .A2(G132), .B1(new_n783), .B2(G125), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT53), .B1(new_n777), .B2(new_n1051), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT54), .B(G143), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n287), .B1(new_n797), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1136), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1134), .A2(new_n1135), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n770), .B1(new_n1131), .B2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1143), .B(new_n767), .C1(new_n308), .C2(new_n831), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT118), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1125), .B1(new_n1126), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1122), .A2(new_n477), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n927), .A2(new_n656), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT117), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n756), .A2(G330), .A3(new_n860), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1122), .A2(new_n931), .B1(new_n1151), .B2(new_n899), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n898), .B1(new_n1122), .B2(new_n860), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1104), .A2(new_n1100), .A3(new_n1099), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1152), .A2(new_n874), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n927), .A2(new_n1147), .A3(KEYINPUT117), .A4(new_n656), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1150), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1124), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1103), .B1(new_n922), .B2(new_n1108), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1123), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1157), .A2(new_n1109), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1159), .A2(new_n720), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1146), .A2(new_n1164), .ZN(G378));
  INV_X1    g0965(.A(new_n720), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT120), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1155), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1167), .B(new_n1169), .C1(new_n1124), .C2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n655), .A2(new_n436), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n697), .A2(new_n412), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1172), .B(new_n1173), .Z(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n941), .A2(new_n703), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1176), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n937), .B2(G330), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n926), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1176), .B1(new_n941), .B2(new_n703), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n937), .A2(G330), .A3(new_n1178), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1181), .A2(new_n925), .A3(new_n902), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1171), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1167), .B1(new_n1163), .B2(new_n1169), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1166), .B1(new_n1187), .B2(KEYINPUT57), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1169), .B1(new_n1124), .B2(new_n1170), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT120), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(new_n1184), .A3(new_n1171), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT121), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT57), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1193), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT121), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1188), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1184), .A2(new_n766), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n767), .B1(G50), .B2(new_n831), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n794), .A2(new_n1133), .B1(new_n796), .B2(new_n842), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n774), .A2(G132), .B1(new_n812), .B2(new_n1139), .ZN(new_n1201));
  INV_X1    g1001(.A(G125), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(new_n780), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1200), .B(new_n1203), .C1(G150), .C2(new_n800), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n792), .A2(G159), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n258), .A2(new_n327), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT119), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(G124), .B2(new_n783), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n792), .A2(G58), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1048), .B1(G68), .B2(new_n800), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n774), .A2(G97), .B1(new_n779), .B2(G116), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n796), .A2(new_n380), .B1(new_n782), .B2(new_n1015), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n794), .A2(new_n541), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1216), .A2(new_n1217), .A3(new_n275), .A4(G41), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT58), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1210), .B(new_n207), .C1(new_n275), .C2(G41), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1212), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1199), .B1(new_n1224), .B2(new_n770), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1178), .B2(new_n817), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1198), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1197), .A2(new_n1228), .ZN(G375));
  NOR2_X1   g1029(.A1(new_n1169), .A2(new_n1155), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1230), .A2(new_n984), .A3(new_n1157), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT122), .Z(new_n1232));
  NAND2_X1  g1032(.A1(new_n899), .A2(new_n816), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n767), .B1(G68), .B2(new_n831), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n777), .A2(new_n215), .B1(new_n782), .B2(new_n620), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT123), .Z(new_n1236));
  AOI22_X1  g1036(.A1(new_n774), .A2(new_n625), .B1(new_n1054), .B2(new_n800), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n833), .B2(new_n780), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n287), .B1(new_n796), .B2(new_n541), .C1(new_n1015), .C2(new_n794), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1236), .A2(new_n1238), .A3(new_n1011), .A4(new_n1239), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1240), .A2(KEYINPUT124), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(KEYINPUT124), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n779), .A2(G132), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n775), .B2(new_n1138), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G159), .B2(new_n812), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n794), .A2(new_n842), .B1(new_n782), .B2(new_n1133), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G150), .B2(new_n797), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n585), .B1(G50), .B2(new_n800), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1213), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1241), .A2(new_n1242), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1234), .B1(new_n1250), .B2(new_n770), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1155), .A2(new_n766), .B1(new_n1233), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1232), .A2(new_n1252), .ZN(G381));
  NAND3_X1  g1053(.A1(new_n1000), .A2(new_n1097), .A3(new_n1029), .ZN(new_n1254));
  OR2_X1    g1054(.A1(G393), .A2(G396), .ZN(new_n1255));
  OR3_X1    g1055(.A1(new_n1254), .A2(G384), .A3(new_n1255), .ZN(new_n1256));
  OR4_X1    g1056(.A1(G378), .A2(new_n1256), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1057(.A(G378), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n853), .A2(G213), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G407), .B(G213), .C1(G375), .C2(new_n1261), .ZN(G409));
  INV_X1    g1062(.A(new_n1255), .ZN(new_n1263));
  AND2_X1   g1063(.A1(G393), .A2(G396), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1263), .A2(KEYINPUT125), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT125), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1267), .A2(new_n1254), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1097), .B1(new_n1000), .B2(new_n1029), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1266), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1254), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1272), .A2(new_n1265), .A3(new_n1269), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1197), .A2(G378), .A3(new_n1228), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1191), .A2(new_n984), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1258), .B1(new_n1277), .B2(new_n1227), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1259), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1230), .B1(KEYINPUT60), .B2(new_n1158), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1168), .A2(KEYINPUT60), .A3(new_n1170), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n720), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1252), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(G384), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1260), .A2(G2897), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1288), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1280), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT126), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1279), .A2(new_n1259), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT62), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1260), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT62), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1295), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1275), .B1(new_n1294), .B2(new_n1301), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1298), .A2(KEYINPUT63), .A3(new_n1295), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT63), .B1(new_n1298), .B2(new_n1295), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1274), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT126), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1291), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1307), .B(new_n1293), .C1(new_n1308), .C2(new_n1298), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1305), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1302), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(G375), .A2(new_n1258), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1276), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1295), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1295), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1313), .A2(new_n1276), .A3(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1315), .A2(new_n1317), .B1(new_n1275), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1274), .A2(KEYINPUT127), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1315), .A2(KEYINPUT127), .A3(new_n1274), .A4(new_n1317), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(G402));
endmodule


