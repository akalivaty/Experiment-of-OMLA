//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT23), .B1(new_n191), .B2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G128), .ZN(new_n194));
  MUX2_X1   g008(.A(new_n192), .B(KEYINPUT23), .S(new_n194), .Z(new_n195));
  XNOR2_X1  g009(.A(G119), .B(G128), .ZN(new_n196));
  XOR2_X1   g010(.A(KEYINPUT24), .B(G110), .Z(new_n197));
  OAI22_X1  g011(.A1(new_n195), .A2(G110), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT16), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  OR2_X1    g016(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(G146), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n198), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(new_n203), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n205), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n204), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n197), .A2(new_n196), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n195), .A2(G110), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OR2_X1    g028(.A1(new_n214), .A2(KEYINPUT75), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(KEYINPUT75), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n208), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G137), .ZN(new_n218));
  INV_X1    g032(.A(G953), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n219), .A2(G221), .A3(G234), .ZN(new_n220));
  XOR2_X1   g034(.A(new_n218), .B(new_n220), .Z(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n217), .B(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n215), .A2(new_n216), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n207), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n222), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n217), .A2(new_n221), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n188), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n190), .B1(new_n224), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n223), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n189), .A2(G902), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT32), .ZN(new_n238));
  INV_X1    g052(.A(G137), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G134), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT11), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n245), .A3(G131), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT64), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G143), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n252), .A2(new_n254), .A3(new_n205), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n205), .A2(G143), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n257), .B(KEYINPUT1), .C1(new_n251), .C2(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n205), .A2(G143), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n257), .B1(new_n260), .B2(KEYINPUT1), .ZN(new_n261));
  OAI22_X1  g075(.A1(new_n255), .A2(new_n256), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G128), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT64), .B(G143), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n260), .B(new_n266), .C1(new_n267), .C2(new_n205), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n262), .A2(new_n263), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n263), .B1(new_n262), .B2(new_n268), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n250), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n258), .A2(G128), .ZN(new_n274));
  INV_X1    g088(.A(new_n261), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n252), .A2(new_n254), .A3(new_n205), .ZN(new_n276));
  INV_X1    g090(.A(new_n256), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n268), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT68), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n262), .A2(new_n263), .A3(new_n268), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT69), .A3(new_n250), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n193), .A2(G116), .ZN(new_n284));
  INV_X1    g098(.A(G116), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G119), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT2), .B(G113), .Z(new_n290));
  XNOR2_X1  g104(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n260), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n252), .A2(new_n254), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(G146), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT0), .A3(G128), .ZN(new_n295));
  NAND2_X1  g109(.A1(KEYINPUT0), .A2(G128), .ZN(new_n296));
  OR2_X1    g110(.A1(KEYINPUT0), .A2(G128), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n296), .B(new_n297), .C1(new_n255), .C2(new_n256), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(KEYINPUT65), .A2(G131), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n246), .B(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n273), .A2(new_n283), .A3(new_n291), .A4(new_n304), .ZN(new_n305));
  XOR2_X1   g119(.A(KEYINPUT26), .B(G101), .Z(new_n306));
  INV_X1    g120(.A(G237), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(new_n219), .A3(G210), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n306), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n250), .B1(new_n278), .B2(new_n279), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(KEYINPUT30), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n273), .A2(new_n283), .A3(new_n304), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(KEYINPUT30), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n305), .B(new_n311), .C1(new_n316), .C2(new_n291), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT31), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n291), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n315), .A2(KEYINPUT30), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(new_n314), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n322), .A2(KEYINPUT31), .A3(new_n305), .A4(new_n311), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n313), .A2(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n305), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT28), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT72), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n271), .A2(new_n291), .A3(new_n304), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT28), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(new_n331), .A3(KEYINPUT28), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n327), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n311), .B(KEYINPUT71), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n319), .A2(new_n323), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(G472), .A2(G902), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(KEYINPUT73), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n238), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n323), .A2(new_n319), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n334), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n337), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(KEYINPUT32), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G472), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n315), .A2(new_n320), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n305), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT28), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n348), .A2(KEYINPUT29), .A3(new_n311), .A4(new_n330), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT74), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n329), .B1(new_n347), .B2(KEYINPUT28), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT29), .A4(new_n311), .ZN(new_n353));
  AOI21_X1  g167(.A(G902), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n322), .A2(new_n305), .ZN(new_n355));
  INV_X1    g169(.A(new_n311), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n357), .B(new_n358), .C1(new_n334), .C2(new_n333), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n345), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n237), .B1(new_n344), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n354), .A2(new_n359), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G472), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n338), .A3(new_n343), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT76), .A3(new_n237), .ZN(new_n367));
  INV_X1    g181(.A(G221), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT9), .B(G234), .Z(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n188), .ZN(new_n370));
  INV_X1    g184(.A(G469), .ZN(new_n371));
  INV_X1    g185(.A(G104), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(G107), .ZN(new_n373));
  NOR2_X1   g187(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n372), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n376));
  OAI22_X1  g190(.A1(new_n372), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n377));
  INV_X1    g191(.A(G101), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n375), .A2(new_n376), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT4), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n380), .B(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n300), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(G101), .B1(new_n386), .B2(new_n373), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n268), .A2(KEYINPUT78), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n293), .A2(G146), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT78), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n260), .A4(new_n266), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n191), .B1(new_n276), .B2(KEYINPUT1), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(new_n294), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n389), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT10), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n384), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n282), .A2(KEYINPUT10), .A3(new_n389), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n302), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n401), .A2(new_n302), .A3(new_n384), .A4(new_n399), .ZN(new_n403));
  XNOR2_X1  g217(.A(G110), .B(G140), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n219), .A2(G227), .ZN(new_n405));
  XOR2_X1   g219(.A(new_n404), .B(new_n405), .Z(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n388), .A2(new_n262), .A3(new_n268), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n397), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n397), .B2(new_n410), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT12), .B1(new_n413), .B2(new_n303), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n397), .A2(new_n410), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT12), .A3(new_n303), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT79), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n415), .A2(new_n418), .A3(KEYINPUT12), .A4(new_n303), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n403), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n406), .ZN(new_n422));
  AOI211_X1 g236(.A(new_n371), .B(new_n408), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n414), .B2(new_n420), .ZN(new_n425));
  INV_X1    g239(.A(new_n407), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n415), .A2(KEYINPUT80), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n397), .A2(new_n409), .A3(new_n410), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n303), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT12), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n431), .A2(KEYINPUT81), .A3(new_n417), .A4(new_n419), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n425), .A2(new_n426), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n403), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n422), .B1(new_n402), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(G902), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n423), .B1(new_n436), .B2(new_n371), .ZN(new_n437));
  NAND2_X1  g251(.A1(G469), .A2(G902), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n370), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(G475), .A2(G902), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G214), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n442), .A2(G237), .A3(G953), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n443), .B1(new_n293), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n307), .A2(new_n219), .A3(G214), .ZN(new_n446));
  NAND2_X1  g260(.A1(KEYINPUT64), .A2(KEYINPUT85), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n251), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n247), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n443), .A2(new_n251), .A3(new_n447), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT85), .B1(new_n252), .B2(new_n254), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n451), .B(G131), .C1(new_n452), .C2(new_n443), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G125), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G140), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n202), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT19), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n454), .B(new_n204), .C1(G146), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT18), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(KEYINPUT86), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n446), .B1(new_n267), .B2(KEYINPUT85), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(new_n451), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n454), .B2(new_n461), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n457), .A2(G146), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT87), .B1(new_n465), .B2(new_n206), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n206), .A3(KEYINPUT87), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT88), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n461), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n450), .B2(new_n453), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n465), .A2(new_n206), .A3(KEYINPUT87), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(new_n466), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n475));
  NOR4_X1   g289(.A1(new_n472), .A2(new_n474), .A3(new_n475), .A4(new_n463), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n459), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G113), .B(G122), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(new_n372), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n453), .ZN(new_n482));
  AOI21_X1  g296(.A(G131), .B1(new_n462), .B2(new_n451), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n461), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n463), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n485), .A3(new_n469), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n475), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n464), .A2(KEYINPUT88), .A3(new_n469), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n210), .A2(new_n204), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n450), .A2(new_n491), .A3(new_n453), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n482), .A2(KEYINPUT17), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n479), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n441), .B1(new_n481), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT20), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT89), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n479), .B1(new_n489), .B2(new_n459), .ZN(new_n500));
  AOI211_X1 g314(.A(new_n480), .B(new_n494), .C1(new_n487), .C2(new_n488), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n498), .B(new_n440), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT90), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n440), .B1(new_n500), .B2(new_n501), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT20), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n497), .A2(new_n507), .A3(new_n498), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n499), .A2(new_n503), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n494), .B1(new_n487), .B2(new_n488), .ZN(new_n510));
  OR3_X1    g324(.A1(new_n510), .A2(KEYINPUT91), .A3(new_n479), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT91), .B1(new_n510), .B2(new_n479), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n501), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G475), .B1(new_n513), .B2(G902), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n369), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n516), .A2(new_n187), .A3(G953), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n293), .A2(G128), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n519), .B(new_n244), .C1(G128), .C2(new_n251), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G122), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G116), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n285), .A2(G122), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(KEYINPUT92), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n523), .B2(new_n524), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(G107), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n385), .B1(new_n526), .B2(new_n529), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n267), .A2(new_n191), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n533), .B1(new_n534), .B2(KEYINPUT13), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n251), .A2(G128), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n534), .B2(KEYINPUT13), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT13), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n519), .A2(KEYINPUT93), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI221_X4 g354(.A(new_n521), .B1(new_n531), .B2(new_n532), .C1(new_n540), .C2(G134), .ZN(new_n541));
  OAI21_X1  g355(.A(G134), .B1(new_n534), .B2(new_n536), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n520), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n522), .A2(G116), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT14), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n523), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(KEYINPUT95), .B(new_n523), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n548), .B(new_n549), .C1(KEYINPUT14), .C2(new_n524), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G107), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n532), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(KEYINPUT94), .B(new_n385), .C1(new_n526), .C2(new_n529), .ZN(new_n554));
  AND4_X1   g368(.A1(new_n543), .A2(new_n551), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n518), .B1(new_n541), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n540), .A2(G134), .B1(new_n531), .B2(new_n532), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n520), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n551), .A2(new_n543), .A3(new_n553), .A4(new_n554), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n517), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n559), .A2(KEYINPUT96), .A3(new_n560), .A4(new_n517), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n188), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT97), .ZN(new_n565));
  INV_X1    g379(.A(G478), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(KEYINPUT15), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  OR2_X1    g383(.A1(new_n564), .A2(KEYINPUT97), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OR3_X1    g385(.A1(new_n564), .A2(KEYINPUT97), .A3(new_n567), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n515), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n299), .A2(G125), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT83), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n262), .A2(new_n455), .A3(new_n268), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT83), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n299), .A2(new_n578), .A3(G125), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n219), .A2(G224), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT84), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n580), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n320), .A2(new_n383), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT5), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n193), .A3(G116), .ZN(new_n586));
  OAI211_X1 g400(.A(G113), .B(new_n586), .C1(new_n289), .C2(new_n585), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n284), .B(new_n290), .C1(new_n287), .C2(new_n288), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n389), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(G110), .B(G122), .Z(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n591), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n584), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(KEYINPUT6), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT6), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n590), .A2(new_n596), .A3(new_n591), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n583), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n581), .A2(KEYINPUT7), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n580), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n587), .A2(new_n588), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n388), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n589), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n591), .B(KEYINPUT8), .Z(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n575), .A2(new_n577), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n599), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n600), .A2(new_n605), .A3(new_n607), .A4(new_n594), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n598), .A2(new_n188), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G210), .B1(G237), .B2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n598), .A2(new_n188), .A3(new_n608), .A4(new_n610), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(G952), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(G953), .ZN(new_n616));
  NAND2_X1  g430(.A1(G234), .A2(G237), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT21), .B(G898), .Z(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n617), .A2(G902), .A3(G953), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n619), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(G214), .B1(G237), .B2(G902), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT82), .Z(new_n627));
  NAND3_X1  g441(.A1(new_n614), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n439), .A2(new_n574), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n363), .A2(new_n367), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G101), .ZN(G3));
  OAI21_X1  g446(.A(G472), .B1(new_n335), .B2(G902), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n341), .A2(new_n342), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n635), .A2(new_n237), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n636), .A2(new_n439), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n562), .A2(new_n638), .A3(new_n563), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n556), .A2(KEYINPUT33), .A3(new_n561), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n641), .A2(G478), .A3(new_n188), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n564), .A2(new_n643), .A3(new_n566), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n643), .B1(new_n564), .B2(new_n566), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n515), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n626), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n612), .B2(new_n613), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n647), .A2(new_n624), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n637), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  AOI21_X1  g468(.A(new_n624), .B1(new_n571), .B2(new_n572), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n499), .A2(new_n506), .A3(new_n502), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n499), .A2(new_n506), .A3(KEYINPUT99), .A4(new_n502), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n655), .A2(new_n658), .A3(new_n514), .A4(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n637), .A2(new_n649), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT35), .B(G107), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  NOR2_X1   g479(.A1(new_n222), .A2(KEYINPUT36), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n217), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n217), .A2(new_n666), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n234), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n224), .A2(new_n231), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(new_n190), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n630), .A2(new_n635), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  OAI211_X1 g489(.A(new_n649), .B(new_n672), .C1(new_n344), .C2(new_n360), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n619), .B1(new_n623), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n658), .A2(new_n514), .A3(new_n659), .A4(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n573), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n433), .A2(new_n435), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n371), .A3(new_n188), .ZN(new_n685));
  INV_X1    g499(.A(new_n423), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n438), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n370), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n676), .A2(new_n683), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n191), .ZN(G30));
  XNOR2_X1  g505(.A(new_n678), .B(KEYINPUT39), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT102), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n614), .B(new_n697), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n515), .A2(new_n573), .A3(new_n626), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n695), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n672), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n347), .A2(new_n334), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n317), .B1(new_n702), .B2(KEYINPUT103), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n702), .A2(KEYINPUT103), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n188), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G472), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n338), .A2(new_n343), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n700), .A2(new_n701), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n267), .ZN(G45));
  INV_X1    g524(.A(new_n344), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n701), .B1(new_n711), .B2(new_n365), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n515), .A2(new_n646), .A3(new_n679), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n712), .A2(new_n439), .A3(new_n649), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  AOI21_X1  g530(.A(new_n371), .B1(new_n684), .B2(new_n188), .ZN(new_n717));
  AOI211_X1 g531(.A(G469), .B(G902), .C1(new_n433), .C2(new_n435), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n717), .A2(new_n718), .A3(new_n370), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n366), .A2(new_n237), .A3(new_n651), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  INV_X1    g536(.A(new_n361), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n662), .A3(new_n649), .A4(new_n719), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NAND2_X1  g539(.A1(new_n684), .A2(new_n188), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G469), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(new_n688), .A3(new_n685), .A4(new_n649), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n717), .A2(new_n718), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n731), .A3(new_n688), .A4(new_n649), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n712), .A2(new_n574), .A3(new_n625), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  NAND4_X1  g549(.A1(new_n515), .A2(new_n573), .A3(new_n626), .A4(new_n614), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n624), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n317), .B(KEYINPUT31), .ZN(new_n738));
  INV_X1    g552(.A(new_n334), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n351), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n342), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n633), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n737), .A2(new_n742), .A3(new_n237), .A4(new_n719), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  AOI21_X1  g558(.A(G902), .B1(new_n339), .B2(new_n340), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n741), .B(new_n672), .C1(new_n745), .C2(new_n345), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n713), .A2(KEYINPUT105), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n515), .A2(new_n646), .A3(new_n748), .A4(new_n679), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n733), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n751), .B1(new_n733), .B2(new_n750), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n455), .ZN(G27));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n338), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n634), .A2(KEYINPUT107), .A3(new_n238), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n365), .A3(new_n758), .A4(new_n343), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n747), .A2(new_n749), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n612), .A2(new_n626), .A3(new_n613), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n689), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n759), .A2(new_n237), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n366), .A2(new_n762), .A3(new_n237), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT42), .B1(new_n747), .B2(new_n749), .ZN(new_n765));
  AOI22_X1  g579(.A1(KEYINPUT42), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NAND4_X1  g581(.A1(new_n366), .A2(new_n762), .A3(new_n237), .A4(new_n682), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n723), .A2(KEYINPUT108), .A3(new_n682), .A4(new_n762), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  OR2_X1    g587(.A1(new_n635), .A2(new_n701), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT109), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT109), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n646), .A2(new_n514), .A3(new_n509), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT43), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n775), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n761), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n408), .B1(new_n421), .B2(new_n422), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT45), .Z(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(G469), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(KEYINPUT46), .A3(new_n438), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n788), .B(G469), .C1(new_n785), .C2(G902), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n685), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n688), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n791), .A2(new_n692), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n775), .A2(KEYINPUT44), .A3(new_n776), .A4(new_n779), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n782), .A2(new_n783), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  NAND2_X1  g610(.A1(new_n791), .A2(KEYINPUT47), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n790), .A2(new_n798), .A3(new_n688), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n366), .A2(new_n237), .A3(new_n761), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n797), .A2(new_n714), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT110), .B(G140), .Z(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(G42));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  INV_X1    g619(.A(new_n670), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n232), .A2(new_n806), .A3(new_n678), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n687), .A2(new_n688), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n811));
  INV_X1    g625(.A(new_n736), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n810), .A2(new_n811), .A3(new_n707), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT113), .B1(new_n439), .B2(new_n807), .ZN(new_n814));
  AND4_X1   g628(.A1(KEYINPUT113), .A2(new_n687), .A3(new_n688), .A4(new_n807), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n812), .B(new_n707), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT114), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n712), .A2(new_n439), .A3(new_n649), .A4(new_n682), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n819), .B(new_n715), .C1(new_n752), .C2(new_n753), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n805), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n753), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n733), .A2(new_n750), .A3(new_n751), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n690), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n813), .A2(new_n817), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n825), .A3(KEYINPUT52), .A4(new_n715), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n680), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n366), .A2(new_n681), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n760), .A2(new_n742), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n831), .A2(new_n672), .A3(new_n762), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n766), .A2(new_n772), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n647), .B1(new_n681), .B2(new_n515), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n636), .A2(new_n439), .A3(new_n629), .A4(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n631), .A2(new_n673), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n720), .A2(new_n743), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n724), .A3(new_n734), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n833), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n804), .B1(new_n827), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n819), .B1(new_n752), .B2(new_n753), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n805), .B1(new_n813), .B2(new_n817), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n819), .B(KEYINPUT112), .C1(new_n752), .C2(new_n753), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n715), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n821), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n838), .A2(new_n836), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n849), .A2(KEYINPUT53), .A3(new_n833), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n840), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(KEYINPUT115), .A3(KEYINPUT54), .ZN(new_n852));
  INV_X1    g666(.A(new_n719), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n853), .A2(new_n618), .A3(new_n761), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n237), .A2(new_n779), .A3(new_n759), .A4(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n619), .A2(new_n779), .A3(new_n237), .A4(new_n742), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n733), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n707), .A2(new_n232), .A3(new_n236), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(new_n647), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n857), .A2(new_n616), .A3(new_n859), .A4(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n858), .A2(new_n648), .A3(new_n719), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT118), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n864), .A2(new_n698), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n797), .A2(new_n799), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n730), .B(KEYINPUT111), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n688), .B1(new_n869), .B2(KEYINPUT117), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(KEYINPUT117), .B2(new_n869), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(new_n783), .A3(new_n858), .ZN(new_n873));
  OR3_X1    g687(.A1(new_n861), .A2(new_n515), .A3(new_n646), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n865), .A2(KEYINPUT118), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n866), .B(new_n875), .C1(new_n864), .C2(new_n698), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n867), .A2(new_n873), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n779), .A2(new_n854), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n746), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT51), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n876), .A2(new_n873), .A3(new_n874), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n882));
  INV_X1    g696(.A(new_n879), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n867), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n863), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  AOI211_X1 g700(.A(new_n886), .B(new_n840), .C1(new_n847), .C2(new_n850), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT115), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n827), .A2(new_n839), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n731), .B1(new_n719), .B2(new_n649), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n574), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n366), .A2(new_n625), .A3(new_n672), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n720), .B(new_n743), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n660), .A2(KEYINPUT100), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n660), .A2(KEYINPUT100), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n649), .A3(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n898), .A2(new_n361), .A3(new_n853), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n890), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n837), .A2(KEYINPUT116), .A3(new_n724), .A4(new_n734), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n766), .A2(new_n772), .A3(new_n832), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n836), .A2(new_n804), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n889), .A2(new_n804), .B1(new_n905), .B2(new_n847), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n888), .B1(new_n906), .B2(new_n886), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n852), .B(new_n885), .C1(new_n887), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n615), .A2(new_n219), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n869), .B(KEYINPUT49), .Z(new_n911));
  NAND3_X1  g725(.A1(new_n860), .A2(new_n688), .A3(new_n627), .ZN(new_n912));
  OR4_X1    g726(.A1(new_n698), .A2(new_n911), .A3(new_n777), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n910), .A2(new_n913), .ZN(G75));
  NOR2_X1   g728(.A1(new_n219), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n906), .A2(new_n188), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT56), .B1(new_n917), .B2(G210), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n595), .A2(new_n597), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n583), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT55), .Z(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n906), .B2(new_n188), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n821), .B2(new_n846), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT53), .B1(new_n827), .B2(new_n839), .ZN(new_n929));
  OAI211_X1 g743(.A(KEYINPUT120), .B(G902), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n924), .B1(new_n931), .B2(new_n611), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n922), .A2(new_n932), .ZN(G51));
  NAND2_X1  g747(.A1(new_n438), .A2(KEYINPUT57), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n438), .A2(KEYINPUT57), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT54), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n889), .A2(new_n804), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n905), .A2(new_n847), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n886), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n934), .B(new_n935), .C1(new_n936), .C2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n684), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n931), .A2(G469), .A3(new_n785), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n915), .B1(new_n941), .B2(new_n942), .ZN(G54));
  NOR2_X1   g757(.A1(new_n500), .A2(new_n501), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(KEYINPUT58), .A2(G475), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n945), .B1(new_n931), .B2(new_n947), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n944), .B(new_n946), .C1(new_n926), .C2(new_n930), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n915), .ZN(G60));
  XNOR2_X1  g764(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n566), .A2(new_n188), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n936), .B2(new_n939), .ZN(new_n954));
  INV_X1    g768(.A(new_n641), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n916), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n852), .B1(new_n887), .B2(new_n907), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n953), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n958), .B2(new_n955), .ZN(G63));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT60), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n669), .B(new_n962), .C1(new_n928), .C2(new_n929), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n916), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n233), .B1(new_n906), .B2(new_n961), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n965), .A2(KEYINPUT122), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n966), .A2(KEYINPUT122), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n966), .A2(KEYINPUT122), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n937), .A2(new_n938), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n223), .B1(new_n971), .B2(new_n962), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n969), .B(new_n970), .C1(new_n964), .C2(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n968), .A2(new_n973), .ZN(G66));
  INV_X1    g788(.A(G224), .ZN(new_n975));
  OAI21_X1  g789(.A(G953), .B1(new_n621), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n848), .B2(G953), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT123), .Z(new_n978));
  INV_X1    g792(.A(G898), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n919), .B1(new_n979), .B2(G953), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n978), .B(new_n980), .ZN(G69));
  XNOR2_X1  g795(.A(new_n316), .B(KEYINPUT124), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(new_n458), .Z(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n795), .A2(new_n801), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n694), .A2(new_n761), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n986), .A2(new_n363), .A3(new_n367), .A4(new_n834), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT125), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n709), .A2(new_n715), .A3(new_n843), .A4(new_n845), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT62), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n985), .B(new_n988), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n984), .B1(new_n994), .B2(G953), .ZN(new_n995));
  NAND2_X1  g809(.A1(G227), .A2(G900), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(G953), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n677), .A2(G953), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT126), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n782), .A2(new_n783), .A3(new_n794), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n759), .A2(new_n237), .A3(new_n812), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n792), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n843), .A2(new_n715), .A3(new_n845), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n801), .A2(new_n766), .A3(new_n772), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n999), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n983), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n995), .A2(new_n997), .A3(new_n1007), .ZN(new_n1008));
  OAI211_X1 g822(.A(G953), .B(new_n996), .C1(new_n1006), .C2(new_n984), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(new_n357), .A2(new_n317), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n851), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT63), .Z(new_n1014));
  AOI21_X1  g828(.A(new_n915), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1014), .B1(new_n993), .B2(new_n849), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n355), .A3(new_n311), .ZN(new_n1017));
  INV_X1    g831(.A(new_n355), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n1005), .A2(new_n848), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1014), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1018), .B(new_n356), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n1015), .A2(new_n1017), .A3(new_n1021), .ZN(G57));
endmodule


