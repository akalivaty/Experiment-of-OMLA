//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G219), .A2(G218), .A3(G221), .A4(G220), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n454), .A2(new_n448), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT71), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT71), .B(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT72), .A3(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n463), .A2(new_n465), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(G101), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT70), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n468), .A2(new_n483), .A3(KEYINPUT69), .A4(G125), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT69), .B1(new_n486), .B2(G125), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n471), .A2(new_n480), .A3(new_n488), .ZN(G160));
  INV_X1    g064(.A(KEYINPUT73), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n470), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n469), .A2(new_n476), .ZN(new_n493));
  OR2_X1    g068(.A1(new_n476), .A2(G112), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n493), .A2(G124), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n476), .A2(G138), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n486), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n466), .A2(new_n468), .A3(new_n501), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(KEYINPUT4), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n466), .A2(G126), .A3(G2105), .A4(new_n468), .ZN(new_n506));
  OR2_X1    g081(.A1(G102), .A2(G2105), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n507), .B(G2104), .C1(G114), .C2(new_n476), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n505), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT74), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n512), .A2(new_n515), .B1(KEYINPUT6), .B2(new_n511), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(KEYINPUT75), .A3(new_n517), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G88), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n522), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G62), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n527), .A2(G50), .B1(G651), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n526), .A2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n524), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n517), .A2(G63), .ZN(new_n539));
  AND3_X1   g114(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n540));
  OAI21_X1  g115(.A(G651), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT76), .B(G51), .Z(new_n542));
  NAND3_X1  g117(.A1(new_n522), .A2(G543), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT7), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n541), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n538), .A2(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n531), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n527), .A2(G52), .B1(G651), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n521), .A2(G90), .A3(new_n523), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  NAND2_X1  g130(.A1(new_n525), .A2(G81), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n531), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n527), .A2(G43), .B1(G651), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n556), .A2(G860), .A3(new_n560), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(new_n525), .A2(G91), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n522), .A2(G53), .A3(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT9), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n511), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n568), .A3(new_n570), .ZN(G299));
  AND3_X1   g146(.A1(new_n541), .A2(new_n543), .A3(new_n546), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n572), .B(KEYINPUT77), .C1(new_n537), .C2(new_n524), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n574), .B1(new_n538), .B2(new_n547), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G286));
  OAI21_X1  g152(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n578));
  INV_X1    g153(.A(G49), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n522), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G87), .ZN(new_n581));
  OAI221_X1 g156(.A(new_n578), .B1(new_n579), .B2(new_n580), .C1(new_n524), .C2(new_n581), .ZN(G288));
  NAND3_X1  g157(.A1(new_n521), .A2(G86), .A3(new_n523), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(G61), .B1(new_n529), .B2(new_n530), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n511), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n588), .A2(KEYINPUT78), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n516), .A2(G48), .A3(G543), .A4(new_n518), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(new_n588), .B2(KEYINPUT78), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n521), .A2(KEYINPUT79), .A3(new_n523), .A4(G86), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n585), .A2(new_n592), .A3(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(new_n511), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n521), .A2(G85), .A3(new_n523), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n527), .A2(G47), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n597), .A2(KEYINPUT80), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(KEYINPUT80), .B1(new_n597), .B2(new_n598), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G301), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n527), .A2(G54), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(new_n511), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n524), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n521), .A2(KEYINPUT10), .A3(new_n523), .A4(G92), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT81), .Z(new_n613));
  AOI21_X1  g188(.A(new_n603), .B1(new_n613), .B2(new_n602), .ZN(G321));
  XNOR2_X1  g189(.A(G321), .B(KEYINPUT82), .ZN(G284));
  NOR2_X1   g190(.A1(G299), .A2(G868), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n576), .B2(G868), .ZN(G297));
  AOI21_X1  g192(.A(new_n616), .B1(new_n576), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n613), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n556), .A2(new_n560), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n619), .ZN(new_n622));
  MUX2_X1   g197(.A(new_n621), .B(new_n622), .S(G868), .Z(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n473), .A2(new_n486), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(KEYINPUT83), .B2(G2100), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n491), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n493), .A2(G123), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n476), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  AOI22_X1  g212(.A1(new_n627), .A2(new_n632), .B1(new_n637), .B2(G2096), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n631), .B(new_n638), .C1(G2096), .C2(new_n637), .ZN(G156));
  XOR2_X1   g214(.A(KEYINPUT15), .B(G2435), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2438), .ZN(new_n641));
  XOR2_X1   g216(.A(G2427), .B(G2430), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT84), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n641), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT85), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n654), .B(G14), .C1(new_n652), .C2(new_n651), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT86), .ZN(G401));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT17), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n659), .B2(new_n657), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT87), .ZN(new_n665));
  INV_X1    g240(.A(new_n662), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n659), .A3(new_n657), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n659), .A2(new_n662), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n668), .B1(new_n658), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n630), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT88), .B(G2096), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  MUX2_X1   g260(.A(new_n685), .B(new_n684), .S(new_n677), .Z(new_n686));
  NOR2_X1   g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G33), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n491), .A2(G139), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n486), .A2(G127), .ZN(new_n697));
  NAND2_X1  g272(.A1(G115), .A2(G2104), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n476), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(KEYINPUT91), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT25), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(KEYINPUT91), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n696), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n695), .B1(new_n706), .B2(new_n694), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G2072), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(G2072), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G21), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G168), .B2(new_n710), .ZN(new_n712));
  AOI211_X1 g287(.A(new_n708), .B(new_n709), .C1(G1966), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n694), .A2(G32), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n491), .A2(G141), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT26), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n473), .A2(G105), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n719), .B(new_n720), .C1(G129), .C2(new_n493), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n714), .B1(new_n722), .B2(new_n694), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT27), .B(G1996), .Z(new_n724));
  OAI21_X1  g299(.A(new_n713), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n723), .B2(new_n724), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n637), .A2(new_n694), .ZN(new_n727));
  OR2_X1    g302(.A1(KEYINPUT30), .A2(G28), .ZN(new_n728));
  NAND2_X1  g303(.A1(KEYINPUT30), .A2(G28), .ZN(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT31), .B(G11), .Z(new_n731));
  NOR3_X1   g306(.A1(new_n727), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n694), .A2(G27), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G164), .B2(new_n694), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G2078), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(G2078), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n732), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n710), .A2(G5), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G171), .B2(new_n710), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1961), .ZN(new_n740));
  NAND2_X1  g315(.A1(G160), .A2(G29), .ZN(new_n741));
  INV_X1    g316(.A(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n742), .B2(KEYINPUT24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(KEYINPUT24), .B2(new_n742), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2084), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G1966), .B2(new_n712), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n737), .A2(new_n740), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n726), .A2(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT93), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n694), .A2(G35), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G162), .B2(new_n694), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT29), .B(G2090), .Z(new_n753));
  XOR2_X1   g328(.A(new_n752), .B(new_n753), .Z(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT94), .B(KEYINPUT23), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n710), .A2(G20), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT95), .B(G1956), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n758), .B(new_n759), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n694), .A2(G26), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT28), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n491), .A2(G140), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n476), .A2(G116), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n493), .A2(G128), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(G29), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  MUX2_X1   g346(.A(G19), .B(new_n621), .S(G16), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1341), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n754), .A2(new_n760), .A3(new_n771), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n613), .A2(new_n710), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G4), .B2(new_n710), .ZN(new_n776));
  INV_X1    g351(.A(G1348), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n774), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n749), .B2(KEYINPUT93), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n694), .A2(G25), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n491), .A2(G131), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n476), .A2(G107), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n493), .A2(G119), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT89), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n782), .B1(new_n790), .B2(new_n694), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT35), .B(G1991), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n793), .A2(KEYINPUT90), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n710), .A2(G22), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G166), .B2(new_n710), .ZN(new_n796));
  INV_X1    g371(.A(G1971), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(G6), .A2(G16), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G305), .B2(new_n710), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT32), .B(G1981), .Z(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n710), .A2(G23), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n578), .B1(new_n580), .B2(new_n579), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n525), .B2(G87), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n804), .B1(new_n806), .B2(new_n710), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT33), .B(G1976), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n798), .A2(new_n802), .A3(new_n803), .A4(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n710), .A2(G24), .ZN(new_n813));
  INV_X1    g388(.A(G290), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n710), .ZN(new_n815));
  INV_X1    g390(.A(G1986), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n794), .A2(new_n811), .A3(new_n812), .A4(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n750), .A2(new_n781), .A3(new_n820), .A4(new_n821), .ZN(G150));
  INV_X1    g397(.A(G150), .ZN(G311));
  NAND2_X1  g398(.A1(G80), .A2(G543), .ZN(new_n824));
  INV_X1    g399(.A(G67), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n531), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n527), .A2(G55), .B1(G651), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n521), .A2(G93), .A3(new_n523), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n828), .B1(new_n827), .B2(new_n829), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G860), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT37), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n621), .B1(new_n830), .B2(new_n831), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n556), .A2(new_n560), .A3(new_n829), .A4(new_n827), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n613), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT97), .ZN(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n834), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT98), .ZN(G145));
  INV_X1    g421(.A(new_n706), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n509), .A2(KEYINPUT100), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n506), .A2(new_n849), .A3(new_n508), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n852));
  INV_X1    g427(.A(new_n468), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n472), .B2(KEYINPUT3), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n500), .B1(new_n854), .B2(new_n501), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n852), .B1(new_n855), .B2(new_n503), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n857), .A2(KEYINPUT99), .A3(new_n502), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n851), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n768), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n717), .A2(new_n721), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n722), .A2(new_n860), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n847), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n491), .A2(G142), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n476), .A2(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n493), .A2(G130), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT101), .B1(new_n783), .B2(new_n787), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n626), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n783), .A2(KEYINPUT101), .A3(new_n787), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n874), .B1(new_n873), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n871), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  INV_X1    g455(.A(new_n871), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n876), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n861), .A2(new_n862), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n722), .A2(new_n860), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n706), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n865), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n883), .B1(new_n865), .B2(new_n886), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n865), .A2(new_n883), .A3(KEYINPUT102), .A4(new_n886), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G162), .B(new_n637), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(G160), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n888), .A2(new_n894), .ZN(new_n896));
  AOI21_X1  g471(.A(G37), .B1(new_n896), .B2(new_n887), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g474(.A1(new_n832), .A2(new_n602), .ZN(new_n900));
  NAND2_X1  g475(.A1(G290), .A2(G288), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n806), .B(new_n596), .C1(new_n599), .C2(new_n600), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(KEYINPUT104), .A3(new_n902), .ZN(new_n906));
  XNOR2_X1  g481(.A(G303), .B(G305), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n907), .A2(KEYINPUT104), .A3(new_n901), .A4(new_n902), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(KEYINPUT105), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT42), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n837), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n622), .B(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G299), .ZN(new_n922));
  INV_X1    g497(.A(new_n612), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT103), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT103), .B1(G299), .B2(new_n612), .ZN(new_n926));
  NAND2_X1  g501(.A1(G299), .A2(new_n612), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT41), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n925), .A2(new_n926), .A3(new_n930), .A4(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n921), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n921), .A2(new_n928), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n919), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n916), .A3(new_n918), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n900), .B1(new_n938), .B2(new_n602), .ZN(G295));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n940), .B(new_n900), .C1(new_n938), .C2(new_n602), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n602), .B1(new_n935), .B2(new_n937), .ZN(new_n942));
  INV_X1    g517(.A(new_n900), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT106), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n941), .A2(new_n944), .ZN(G331));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n573), .A2(new_n575), .A3(G171), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(G168), .B2(G301), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n573), .A2(new_n575), .A3(new_n948), .A4(G171), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n920), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n837), .A3(new_n951), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n929), .A2(new_n953), .A3(new_n931), .A4(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n954), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n837), .B1(new_n950), .B2(new_n951), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n928), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(new_n913), .A3(new_n914), .ZN(new_n960));
  INV_X1    g535(.A(G37), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(KEYINPUT108), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT108), .B1(new_n960), .B2(new_n961), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n909), .A2(KEYINPUT105), .A3(new_n910), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT105), .B1(new_n909), .B2(new_n910), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n966), .B1(new_n969), .B2(new_n959), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n915), .A2(KEYINPUT109), .A3(new_n958), .A4(new_n955), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n946), .B1(new_n965), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT43), .B1(new_n970), .B2(new_n971), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n960), .A2(new_n961), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n973), .A2(new_n977), .A3(KEYINPUT44), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n965), .A2(new_n974), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n972), .A2(new_n980), .A3(new_n976), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n972), .B2(new_n976), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n978), .B1(new_n984), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n856), .A2(new_n858), .ZN(new_n987));
  INV_X1    g562(.A(new_n850), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n849), .B1(new_n506), .B2(new_n508), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n986), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n471), .A2(new_n480), .A3(new_n488), .A4(G40), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n862), .A2(G1996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n768), .A2(G2067), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n763), .A2(new_n770), .A3(new_n767), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n862), .B2(G1996), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n996), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n788), .B(new_n792), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n996), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n995), .A2(new_n816), .A3(new_n814), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n995), .A2(G1986), .A3(G290), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n1009), .B(KEYINPUT111), .Z(new_n1010));
  NOR2_X1   g585(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n585), .A2(new_n592), .A3(new_n1012), .A4(new_n593), .ZN(new_n1013));
  INV_X1    g588(.A(new_n588), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n583), .A2(new_n1014), .A3(new_n590), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G1981), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT113), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT49), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT113), .B(KEYINPUT49), .C1(new_n1013), .C2(new_n1016), .ZN(new_n1020));
  INV_X1    g595(.A(new_n994), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n859), .A2(new_n1021), .A3(new_n986), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT112), .B(G8), .Z(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1019), .A2(new_n1020), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n806), .A2(G1976), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(G288), .B2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1031), .A2(new_n1022), .A3(new_n1024), .A4(new_n1027), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1026), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G303), .A2(G8), .ZN(new_n1035));
  XOR2_X1   g610(.A(new_n1035), .B(KEYINPUT55), .Z(new_n1036));
  INV_X1    g611(.A(G8), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n986), .B1(new_n505), .B2(new_n509), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n992), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1021), .B(new_n1039), .C1(new_n991), .C2(new_n992), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n797), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n859), .A2(new_n1042), .A3(new_n986), .ZN(new_n1043));
  INV_X1    g618(.A(G2090), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n994), .B1(new_n1038), .B2(KEYINPUT50), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1037), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1034), .A2(new_n1036), .A3(new_n1047), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1026), .A2(G1976), .A3(G288), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1013), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT114), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1049), .A2(KEYINPUT114), .A3(new_n1050), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1048), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(new_n1036), .A3(G8), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1042), .B1(new_n859), .B2(new_n986), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(new_n994), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n857), .A2(KEYINPUT99), .A3(new_n502), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT99), .B1(new_n857), .B2(new_n502), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1384), .B1(new_n1062), .B2(new_n851), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT115), .B(new_n1021), .C1(new_n1063), .C2(new_n1042), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1038), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1042), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1059), .A2(new_n1064), .A3(new_n1044), .A4(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1023), .B1(new_n1067), .B2(new_n1041), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1034), .B(new_n1056), .C1(new_n1068), .C2(new_n1036), .ZN(new_n1069));
  INV_X1    g644(.A(G1966), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT45), .B1(new_n859), .B2(new_n986), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1021), .B1(new_n1038), .B2(new_n992), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G2084), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1043), .A2(new_n1074), .A3(new_n1045), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(new_n576), .A3(new_n1024), .ZN(new_n1077));
  OR3_X1    g652(.A1(new_n1069), .A2(KEYINPUT116), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT63), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT116), .B1(new_n1069), .B2(new_n1077), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1034), .A2(new_n1056), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1083), .B(new_n1084), .C1(new_n1036), .C2(new_n1047), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1054), .B1(new_n1081), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G168), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n994), .B1(new_n1065), .B2(KEYINPUT45), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1966), .B1(new_n993), .B2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1043), .A2(new_n1074), .A3(new_n1045), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1087), .B(new_n1024), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(G168), .A2(new_n1023), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1037), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1091), .B(KEYINPUT51), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1076), .A2(new_n1024), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1092), .A2(KEYINPUT51), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT62), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT118), .ZN(new_n1100));
  INV_X1    g675(.A(G1961), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1043), .A2(new_n1102), .A3(new_n1045), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1040), .B2(G2078), .ZN(new_n1106));
  INV_X1    g681(.A(G2078), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n993), .A2(KEYINPUT53), .A3(new_n1107), .A4(new_n1088), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G171), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1098), .A2(new_n1110), .A3(new_n1069), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1111), .A2(new_n1112), .B1(new_n1114), .B2(KEYINPUT62), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1067), .A2(new_n1041), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1024), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1036), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1110), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1083), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT123), .B1(new_n1121), .B2(new_n1098), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT124), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1098), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1069), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1112), .A3(new_n1120), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1114), .A2(KEYINPUT62), .ZN(new_n1127));
  AND4_X1   g702(.A1(KEYINPUT124), .A2(new_n1122), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1086), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n994), .B1(new_n1063), .B2(KEYINPUT45), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1130), .A2(KEYINPUT53), .A3(new_n1107), .A4(new_n993), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1104), .A2(new_n1106), .A3(new_n1131), .ZN(new_n1132));
  OR3_X1    g707(.A1(new_n1132), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT122), .B1(new_n1132), .B2(G171), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1133), .B(new_n1134), .C1(new_n1120), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1132), .A2(G171), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1137), .B(KEYINPUT54), .C1(G171), .C2(new_n1109), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1136), .A2(new_n1138), .A3(new_n1125), .A4(new_n1114), .ZN(new_n1139));
  XOR2_X1   g714(.A(G299), .B(KEYINPUT57), .Z(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1066), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n994), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(KEYINPUT115), .ZN(new_n1144));
  AOI21_X1  g719(.A(G1956), .B1(new_n1144), .B2(new_n1059), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(G2072), .Z(new_n1147));
  NAND3_X1  g722(.A1(new_n1130), .A2(new_n1039), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1141), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(G1956), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1143), .A2(KEYINPUT115), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(new_n1148), .A3(new_n1140), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1150), .A2(KEYINPUT61), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT120), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1150), .A2(new_n1155), .A3(new_n1158), .A4(KEYINPUT61), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1145), .A2(new_n1149), .A3(new_n1141), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1140), .B1(new_n1154), .B2(new_n1148), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(KEYINPUT58), .B(G1341), .Z(new_n1164));
  NAND2_X1  g739(.A1(new_n1022), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1040), .B2(G1996), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n621), .A2(KEYINPUT119), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT59), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1157), .A2(new_n1159), .A3(new_n1163), .A4(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT121), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n1174), .B2(new_n1160), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1175), .A2(new_n1176), .A3(new_n1157), .A4(new_n1159), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1022), .A2(G2067), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1178), .B1(new_n1179), .B2(new_n777), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(KEYINPUT60), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(new_n612), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(KEYINPUT60), .B2(new_n1180), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1173), .A2(new_n1177), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1180), .A2(new_n923), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1155), .B1(new_n1185), .B2(new_n1162), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1139), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1011), .B1(new_n1129), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n790), .A2(new_n792), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1000), .B1(new_n1003), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n1192), .A2(new_n1193), .A3(new_n996), .ZN(new_n1194));
  INV_X1    g769(.A(G1996), .ZN(new_n1195));
  AOI211_X1 g770(.A(new_n1001), .B(new_n862), .C1(KEYINPUT46), .C2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT46), .B1(new_n995), .B2(new_n1195), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n1198));
  AND2_X1   g773(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1200));
  OAI22_X1  g775(.A1(new_n1196), .A2(new_n996), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT47), .Z(new_n1202));
  XOR2_X1   g777(.A(new_n1007), .B(KEYINPUT48), .Z(new_n1203));
  NOR2_X1   g778(.A1(new_n1006), .A2(new_n1203), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1194), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1188), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n1208));
  INV_X1    g782(.A(KEYINPUT108), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n975), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g784(.A1(new_n972), .A2(new_n1210), .A3(new_n962), .ZN(new_n1211));
  AOI22_X1  g785(.A1(new_n1211), .A2(KEYINPUT43), .B1(new_n976), .B2(new_n974), .ZN(new_n1212));
  NOR3_X1   g786(.A1(G229), .A2(new_n460), .A3(G227), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n896), .A2(new_n887), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n1214), .A2(new_n961), .ZN(new_n1215));
  INV_X1    g789(.A(new_n894), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1216), .B1(new_n890), .B2(new_n891), .ZN(new_n1217));
  OAI211_X1 g791(.A(new_n655), .B(new_n1213), .C1(new_n1215), .C2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g792(.A(new_n1208), .B1(new_n1212), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n1213), .A2(new_n655), .ZN(new_n1220));
  AOI21_X1  g794(.A(new_n1220), .B1(new_n895), .B2(new_n897), .ZN(new_n1221));
  OAI211_X1 g795(.A(new_n1221), .B(KEYINPUT127), .C1(new_n973), .C2(new_n977), .ZN(new_n1222));
  AND2_X1   g796(.A1(new_n1219), .A2(new_n1222), .ZN(G308));
  NAND2_X1  g797(.A1(new_n1219), .A2(new_n1222), .ZN(G225));
endmodule


