//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938;
  AND2_X1   g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(G141gat), .B(G148gat), .Z(new_n203));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT2), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT76), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT76), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G155gat), .B2(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT77), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(KEYINPUT77), .A3(new_n204), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n206), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n203), .A2(new_n205), .ZN(new_n218));
  AND2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT71), .B(KEYINPUT22), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT72), .B(G218gat), .ZN(new_n224));
  INV_X1    g023(.A(G211gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G197gat), .B(G204gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT29), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n222), .B1(new_n233), .B2(KEYINPUT3), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n202), .B1(new_n234), .B2(KEYINPUT81), .ZN(new_n235));
  INV_X1    g034(.A(G22gat), .ZN(new_n236));
  OR2_X1    g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI211_X1 g036(.A(G22gat), .B(new_n202), .C1(new_n234), .C2(KEYINPUT81), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT31), .B(G50gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(new_n217), .B2(new_n221), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n232), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n234), .ZN(new_n250));
  XNOR2_X1  g049(.A(G78gat), .B(G106gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n250), .B(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n235), .A2(new_n236), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n240), .B1(new_n254), .B2(new_n238), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n242), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n253), .B1(new_n255), .B2(new_n242), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G225gat), .A2(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n260));
  INV_X1    g059(.A(G127gat), .ZN(new_n261));
  INV_X1    g060(.A(G134gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G127gat), .A2(G134gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n263), .A2(new_n264), .B1(KEYINPUT70), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G113gat), .B(G120gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n268), .A2(KEYINPUT1), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n266), .B1(KEYINPUT1), .B2(new_n268), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT77), .B1(new_n212), .B2(new_n204), .ZN(new_n272));
  AOI211_X1 g071(.A(new_n214), .B(new_n219), .C1(new_n209), .C2(new_n211), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n218), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n219), .A2(new_n220), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n206), .A2(new_n275), .ZN(new_n276));
  AOI221_X4 g075(.A(new_n260), .B1(new_n270), .B2(new_n271), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n276), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(new_n271), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT4), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n279), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n274), .A2(KEYINPUT3), .A3(new_n276), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n244), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n259), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT39), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT0), .ZN(new_n289));
  XNOR2_X1  g088(.A(G57gat), .B(G85gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT82), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n282), .A2(new_n274), .A3(new_n276), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n279), .B1(new_n217), .B2(new_n221), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n259), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT39), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n285), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT40), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  AND4_X1   g099(.A1(KEYINPUT40), .A2(new_n299), .A3(new_n292), .A4(new_n287), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n295), .A2(new_n260), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n278), .A2(KEYINPUT4), .A3(new_n279), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n297), .A2(KEYINPUT5), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n284), .A2(new_n302), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n281), .A2(KEYINPUT78), .A3(new_n284), .A4(new_n304), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n284), .A2(new_n302), .A3(new_n303), .A4(new_n259), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT5), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(new_n296), .B2(new_n297), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n307), .A2(new_n308), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(new_n292), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n300), .A2(new_n301), .A3(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G8gat), .B(G36gat), .Z(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT75), .ZN(new_n316));
  XNOR2_X1  g115(.A(G64gat), .B(G92gat), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n316), .B(new_n317), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT25), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n321));
  NAND3_X1  g120(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(G183gat), .B2(G190gat), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT23), .ZN(new_n327));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n329), .B1(G169gat), .B2(G176gat), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n324), .ZN(new_n332));
  INV_X1    g131(.A(G183gat), .ZN(new_n333));
  INV_X1    g132(.A(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n332), .A2(KEYINPUT64), .A3(new_n335), .A4(new_n322), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n325), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n323), .B1(KEYINPUT65), .B2(new_n332), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n332), .A2(KEYINPUT65), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AND4_X1   g139(.A1(KEYINPUT25), .A2(new_n327), .A3(new_n328), .A4(new_n330), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n320), .A2(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n326), .A2(KEYINPUT26), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n333), .B2(new_n334), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT26), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(new_n326), .ZN(new_n347));
  OR2_X1    g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT27), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G183gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n333), .A2(KEYINPUT27), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT68), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT68), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n334), .A2(KEYINPUT28), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n333), .A2(KEYINPUT27), .ZN(new_n359));
  AOI21_X1  g158(.A(G190gat), .B1(new_n359), .B2(KEYINPUT66), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT66), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT27), .B1(new_n361), .B2(new_n333), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n348), .B1(new_n358), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT73), .B1(new_n342), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n337), .A2(new_n320), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n340), .A2(new_n341), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n344), .A2(new_n347), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n334), .A2(KEYINPUT28), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n374), .B1(new_n354), .B2(new_n355), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n364), .B1(new_n360), .B2(new_n362), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n371), .A2(new_n372), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n368), .A2(new_n378), .A3(new_n245), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT69), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(KEYINPUT69), .B(new_n373), .C1(new_n375), .C2(new_n376), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n371), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n380), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n248), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n381), .A2(KEYINPUT74), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n378), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n386), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(new_n245), .A3(new_n380), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n248), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT74), .B1(new_n381), .B2(new_n387), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n319), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT30), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n319), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n396), .A2(new_n392), .A3(new_n388), .A4(new_n398), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n393), .A2(new_n319), .A3(new_n394), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n395), .B(new_n399), .C1(new_n400), .C2(KEYINPUT30), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n258), .B1(new_n314), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n393), .A2(new_n394), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT37), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n318), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n390), .A2(new_n391), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n404), .B1(new_n406), .B2(new_n247), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n247), .B1(new_n385), .B2(new_n386), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n381), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT38), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n291), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n307), .A2(new_n308), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n309), .A2(new_n311), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT80), .B1(new_n415), .B2(KEYINPUT6), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418));
  NOR4_X1   g217(.A1(new_n312), .A2(new_n417), .A3(new_n418), .A4(new_n412), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n400), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n291), .B1(new_n309), .B2(new_n311), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT6), .B1(new_n413), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(new_n312), .B2(new_n292), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n411), .A2(new_n420), .A3(new_n421), .A4(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT38), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT37), .B1(new_n393), .B2(new_n394), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n405), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n402), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n413), .A2(new_n422), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT79), .B1(new_n430), .B2(KEYINPUT6), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n414), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n291), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT79), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n423), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n420), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n258), .B1(new_n438), .B2(new_n401), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n385), .A2(new_n279), .ZN(new_n440));
  INV_X1    g239(.A(G227gat), .ZN(new_n441));
  INV_X1    g240(.A(G233gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n383), .A2(new_n371), .A3(new_n384), .A4(new_n282), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XOR2_X1   g246(.A(G15gat), .B(G43gat), .Z(new_n448));
  XNOR2_X1  g247(.A(G71gat), .B(G99gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT34), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n440), .A2(new_n444), .ZN(new_n453));
  INV_X1    g252(.A(new_n443), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI211_X1 g255(.A(KEYINPUT34), .B(new_n443), .C1(new_n440), .C2(new_n444), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n451), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n445), .A2(KEYINPUT32), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n450), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n445), .B2(new_n446), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n455), .B2(new_n457), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n459), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n461), .B1(new_n459), .B2(new_n464), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT36), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n429), .A2(new_n439), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT83), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n465), .B2(new_n466), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n459), .A2(new_n464), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n460), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n459), .A2(new_n461), .A3(new_n464), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(KEYINPUT83), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT35), .B1(new_n420), .B2(new_n424), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n401), .A2(new_n258), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT35), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n401), .B1(new_n436), .B2(new_n420), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n258), .A2(new_n465), .A3(new_n466), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT84), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI211_X1 g284(.A(KEYINPUT84), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n469), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT89), .ZN(new_n488));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT15), .ZN(new_n490));
  NOR2_X1   g289(.A1(G29gat), .A2(G36gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT14), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(G29gat), .ZN(new_n494));
  INV_X1    g293(.A(G36gat), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT85), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR3_X1    g295(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT85), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n490), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(KEYINPUT15), .A3(new_n489), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n501), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT86), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT16), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(G1gat), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(G1gat), .B2(new_n508), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(G8gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n504), .A2(new_n506), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n502), .A2(KEYINPUT17), .B1(KEYINPUT88), .B2(new_n512), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n512), .A2(KEYINPUT88), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n513), .B(new_n514), .C1(new_n517), .C2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT18), .ZN(new_n522));
  INV_X1    g321(.A(new_n512), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n513), .A2(new_n524), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n514), .B(KEYINPUT13), .Z(new_n526));
  AOI22_X1  g325(.A1(new_n521), .A2(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G113gat), .B(G141gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(G197gat), .ZN(new_n529));
  XOR2_X1   g328(.A(KEYINPUT11), .B(G169gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n531), .B(KEYINPUT12), .Z(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n517), .A2(new_n520), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n534), .A2(KEYINPUT18), .A3(new_n514), .A4(new_n513), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n527), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n533), .B1(new_n527), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n488), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n527), .A2(new_n535), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n532), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n527), .A2(new_n533), .A3(new_n535), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT89), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n487), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545));
  INV_X1    g344(.A(G85gat), .ZN(new_n546));
  INV_X1    g345(.A(G92gat), .ZN(new_n547));
  AOI22_X1  g346(.A1(KEYINPUT8), .A2(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT94), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT7), .ZN(new_n550));
  OAI211_X1 g349(.A(G85gat), .B(G92gat), .C1(new_n550), .C2(KEYINPUT93), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(KEYINPUT93), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G99gat), .B(G106gat), .Z(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n554), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT9), .ZN(new_n558));
  XOR2_X1   g357(.A(G57gat), .B(G64gat), .Z(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(KEYINPUT90), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(KEYINPUT90), .B2(new_n559), .ZN(new_n561));
  XNOR2_X1  g360(.A(G71gat), .B(G78gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT91), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n559), .A2(new_n562), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n561), .A2(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n557), .A2(KEYINPUT10), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n557), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(KEYINPUT95), .B2(new_n556), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n557), .B(new_n567), .C1(KEYINPUT95), .C2(new_n556), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT10), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT96), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT96), .A4(new_n573), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n568), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G230gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(new_n442), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n571), .A2(new_n572), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n580), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G120gat), .B(G148gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT97), .ZN(new_n587));
  XNOR2_X1  g386(.A(G176gat), .B(G204gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(new_n584), .A3(new_n589), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n595));
  NOR2_X1   g394(.A1(new_n567), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G127gat), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n512), .B1(new_n567), .B2(KEYINPUT21), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G155gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n507), .A2(new_n557), .B1(KEYINPUT41), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n557), .B1(KEYINPUT17), .B2(new_n502), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(new_n515), .B2(new_n516), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n614), .B(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n610), .A2(KEYINPUT41), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n617), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n594), .A2(new_n609), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n544), .A2(new_n438), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G1gat), .ZN(G1324gat));
  INV_X1    g424(.A(KEYINPUT42), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n544), .A2(new_n401), .A3(new_n623), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT98), .Z(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT16), .B(G8gat), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(G8gat), .ZN(new_n631));
  OR3_X1    g430(.A1(new_n627), .A2(new_n626), .A3(new_n629), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(G1325gat));
  NAND2_X1  g432(.A1(new_n544), .A2(new_n623), .ZN(new_n634));
  OAI21_X1  g433(.A(G15gat), .B1(new_n634), .B2(new_n468), .ZN(new_n635));
  INV_X1    g434(.A(new_n623), .ZN(new_n636));
  INV_X1    g435(.A(new_n476), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n636), .A2(G15gat), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n544), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT99), .ZN(G1326gat));
  INV_X1    g440(.A(new_n258), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n634), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT43), .B(G22gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(G1327gat));
  NOR3_X1   g444(.A1(new_n594), .A2(new_n608), .A3(new_n621), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n544), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n647), .A2(G29gat), .A3(new_n437), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT45), .Z(new_n649));
  NAND3_X1  g448(.A1(new_n487), .A2(KEYINPUT100), .A3(new_n622), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n487), .A2(KEYINPUT100), .A3(KEYINPUT44), .A4(new_n622), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n540), .A2(new_n541), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n594), .A2(new_n608), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT101), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n652), .A2(new_n659), .A3(new_n653), .A4(new_n656), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n658), .A2(new_n438), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n649), .B1(new_n494), .B2(new_n661), .ZN(G1328gat));
  INV_X1    g461(.A(new_n401), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n647), .A2(G36gat), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT46), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n658), .A2(new_n401), .A3(new_n660), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n495), .B2(new_n666), .ZN(G1329gat));
  OAI21_X1  g466(.A(G43gat), .B1(new_n657), .B2(new_n468), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n647), .A2(G43gat), .A3(new_n637), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n670), .A3(KEYINPUT47), .ZN(new_n671));
  INV_X1    g470(.A(new_n468), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n658), .A2(new_n672), .A3(new_n660), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n674));
  AND3_X1   g473(.A1(new_n673), .A2(new_n674), .A3(G43gat), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n674), .B1(new_n673), .B2(G43gat), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n675), .A2(new_n676), .A3(new_n669), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n671), .B1(new_n677), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g477(.A(G50gat), .B1(new_n657), .B2(new_n642), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n647), .A2(G50gat), .A3(new_n642), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n681), .A3(KEYINPUT48), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n658), .A2(new_n258), .A3(new_n660), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n680), .B1(new_n683), .B2(G50gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n682), .B1(new_n684), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g484(.A1(new_n609), .A2(new_n593), .A3(new_n622), .A4(new_n654), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n487), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n438), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g488(.A(new_n663), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n691), .B(KEYINPUT103), .Z(new_n692));
  NOR2_X1   g491(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1333gat));
  NAND3_X1  g493(.A1(new_n687), .A2(G71gat), .A3(new_n672), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT104), .Z(new_n696));
  AND2_X1   g495(.A1(new_n687), .A2(new_n476), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(G71gat), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1334gat));
  NAND2_X1  g499(.A1(new_n687), .A2(new_n258), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g501(.A1(new_n608), .A2(new_n654), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n487), .A2(new_n622), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT51), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n705), .A2(KEYINPUT107), .A3(KEYINPUT51), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n708), .B(new_n709), .C1(KEYINPUT51), .C2(new_n705), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n710), .A2(new_n546), .A3(new_n438), .A4(new_n594), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n593), .A2(new_n608), .A3(new_n654), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n652), .A2(new_n653), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT106), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n652), .A2(new_n715), .A3(new_n653), .A4(new_n712), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n714), .A2(new_n438), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n711), .B1(new_n546), .B2(new_n717), .ZN(G1336gat));
  NAND3_X1  g517(.A1(new_n594), .A2(new_n547), .A3(new_n401), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n710), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722));
  OAI21_X1  g521(.A(G92gat), .B1(new_n713), .B2(new_n663), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n714), .A2(new_n401), .A3(new_n716), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G92gat), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT51), .B1(new_n704), .B2(KEYINPUT108), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n487), .A2(new_n729), .A3(new_n622), .A4(new_n703), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(KEYINPUT109), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n706), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT109), .B1(new_n728), .B2(new_n730), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n720), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n725), .B1(new_n735), .B2(KEYINPUT52), .ZN(new_n736));
  AOI211_X1 g535(.A(KEYINPUT110), .B(new_n722), .C1(new_n727), .C2(new_n734), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n724), .B1(new_n736), .B2(new_n737), .ZN(G1337gat));
  NAND3_X1  g537(.A1(new_n714), .A2(new_n672), .A3(new_n716), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G99gat), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n593), .A2(new_n637), .A3(G99gat), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(KEYINPUT111), .Z(new_n742));
  NAND2_X1  g541(.A1(new_n710), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(G1338gat));
  NOR3_X1   g543(.A1(new_n593), .A2(G106gat), .A3(new_n642), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n710), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n747));
  OAI21_X1  g546(.A(G106gat), .B1(new_n713), .B2(new_n642), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n732), .A2(new_n733), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n714), .A2(new_n258), .A3(new_n716), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n750), .A2(new_n745), .B1(new_n751), .B2(G106gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n752), .B2(new_n747), .ZN(G1339gat));
  INV_X1    g552(.A(new_n580), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n576), .A2(new_n577), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n754), .B(new_n755), .C1(new_n756), .C2(new_n568), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n578), .A2(new_n580), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT54), .B1(new_n578), .B2(new_n580), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n757), .B(new_n590), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n592), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n582), .A2(KEYINPUT54), .A3(new_n758), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n589), .B1(new_n581), .B2(new_n755), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT55), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT113), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n761), .A2(new_n762), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n764), .A2(new_n765), .A3(KEYINPUT55), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .A4(new_n592), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(new_n654), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n514), .B1(new_n534), .B2(new_n513), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n525), .A2(new_n526), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n531), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n541), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n593), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n622), .B1(new_n772), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n767), .A2(new_n771), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n541), .A2(new_n775), .A3(KEYINPUT114), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n622), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n609), .B1(new_n779), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n623), .A2(new_n655), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n437), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n788), .A2(new_n467), .A3(new_n478), .ZN(new_n789));
  AOI21_X1  g588(.A(G113gat), .B1(new_n789), .B2(new_n654), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(new_n478), .A3(new_n476), .ZN(new_n791));
  INV_X1    g590(.A(G113gat), .ZN(new_n792));
  INV_X1    g591(.A(new_n543), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n790), .A2(new_n794), .ZN(G1340gat));
  AOI21_X1  g594(.A(G120gat), .B1(new_n789), .B2(new_n594), .ZN(new_n796));
  INV_X1    g595(.A(G120gat), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n791), .A2(new_n797), .A3(new_n593), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n796), .A2(new_n798), .ZN(G1341gat));
  NAND3_X1  g598(.A1(new_n789), .A2(new_n261), .A3(new_n608), .ZN(new_n800));
  OAI21_X1  g599(.A(G127gat), .B1(new_n791), .B2(new_n609), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1342gat));
  NAND3_X1  g601(.A1(new_n789), .A2(new_n262), .A3(new_n622), .ZN(new_n803));
  OR2_X1    g602(.A1(new_n803), .A2(KEYINPUT56), .ZN(new_n804));
  OAI21_X1  g603(.A(G134gat), .B1(new_n791), .B2(new_n621), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(KEYINPUT56), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(G1343gat));
  NOR3_X1   g606(.A1(new_n672), .A2(new_n401), .A3(new_n437), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n786), .A2(new_n787), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT57), .B1(new_n809), .B2(new_n258), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n642), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n793), .A2(new_n763), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT55), .B1(new_n761), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n815), .B2(new_n761), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n777), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n622), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n609), .B1(new_n819), .B2(new_n785), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n813), .B1(new_n820), .B2(new_n787), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n808), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G141gat), .B1(new_n822), .B2(new_n793), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n468), .A2(new_n258), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n663), .B1(new_n824), .B2(KEYINPUT116), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(KEYINPUT116), .B2(new_n824), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n788), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n793), .A2(G141gat), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT58), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n823), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n654), .B(new_n808), .C1(new_n810), .C2(new_n821), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n832), .A2(G141gat), .B1(new_n828), .B2(new_n829), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(G1344gat));
  INV_X1    g634(.A(G148gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n828), .A2(new_n836), .A3(new_n594), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n808), .A2(new_n594), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n636), .A2(new_n543), .ZN(new_n840));
  INV_X1    g639(.A(new_n763), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n768), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n818), .A2(new_n622), .B1(new_n842), .B2(new_n784), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n840), .B1(new_n843), .B2(new_n609), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n811), .B1(new_n844), .B2(new_n642), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n813), .B1(new_n786), .B2(new_n787), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n839), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n836), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n842), .A2(new_n784), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n817), .A2(new_n543), .A3(new_n841), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n778), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n851), .B1(new_n853), .B2(new_n621), .ZN(new_n854));
  OAI22_X1  g653(.A1(new_n854), .A2(new_n608), .B1(new_n543), .B2(new_n636), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n258), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n846), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n857), .B2(new_n839), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n838), .B1(new_n850), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n822), .A2(new_n593), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(KEYINPUT59), .A3(new_n836), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n837), .B1(new_n859), .B2(new_n861), .ZN(G1345gat));
  NOR3_X1   g661(.A1(new_n822), .A2(new_n207), .A3(new_n609), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT118), .B1(new_n827), .B2(new_n609), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n827), .A2(KEYINPUT118), .A3(new_n609), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(G155gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(G1346gat));
  NAND3_X1  g666(.A1(new_n828), .A2(new_n208), .A3(new_n622), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT119), .B1(new_n822), .B2(new_n621), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G162gat), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n822), .A2(KEYINPUT119), .A3(new_n621), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(G1347gat));
  AOI21_X1  g671(.A(new_n438), .B1(new_n786), .B2(new_n787), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n873), .A2(new_n401), .A3(new_n482), .ZN(new_n874));
  AOI21_X1  g673(.A(G169gat), .B1(new_n874), .B2(new_n654), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n873), .A2(new_n401), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n637), .A2(new_n258), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n543), .A2(G169gat), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n875), .B1(new_n878), .B2(new_n879), .ZN(G1348gat));
  INV_X1    g679(.A(G176gat), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n593), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n876), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT121), .ZN(new_n884));
  AOI211_X1 g683(.A(KEYINPUT120), .B(G176gat), .C1(new_n874), .C2(new_n594), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n874), .A2(new_n594), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n881), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n884), .A2(new_n885), .A3(new_n888), .ZN(G1349gat));
  AND2_X1   g688(.A1(new_n608), .A2(new_n356), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n873), .A2(new_n401), .A3(new_n608), .A4(new_n877), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n874), .A2(new_n890), .B1(new_n891), .B2(G183gat), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT60), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT122), .B1(new_n892), .B2(new_n893), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n892), .B2(KEYINPUT122), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n896), .B1(new_n897), .B2(new_n899), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n874), .A2(new_n334), .A3(new_n622), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n873), .A2(new_n401), .A3(new_n622), .A4(new_n877), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n902), .A2(new_n903), .A3(G190gat), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n903), .B1(new_n902), .B2(G190gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT124), .B(new_n901), .C1(new_n904), .C2(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1351gat));
  NOR2_X1   g709(.A1(new_n672), .A2(new_n663), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n258), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT125), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n873), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(G197gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n915), .A3(new_n654), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT126), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n911), .A2(new_n437), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n856), .B2(new_n846), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n845), .A2(new_n847), .A3(KEYINPUT127), .ZN(new_n921));
  AOI211_X1 g720(.A(new_n793), .B(new_n918), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n917), .B1(new_n915), .B2(new_n922), .ZN(G1352gat));
  INV_X1    g722(.A(G204gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n914), .A2(new_n924), .A3(new_n594), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT62), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n925), .A2(KEYINPUT62), .ZN(new_n927));
  AOI211_X1 g726(.A(new_n593), .B(new_n918), .C1(new_n920), .C2(new_n921), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n926), .B(new_n927), .C1(new_n928), .C2(new_n924), .ZN(G1353gat));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n225), .A3(new_n608), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n918), .A2(new_n609), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n856), .B2(new_n846), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n932), .B2(G211gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G1354gat));
  AOI21_X1  g734(.A(G218gat), .B1(new_n914), .B2(new_n622), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n621), .A2(new_n224), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(G1355gat));
endmodule


