//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1257, new_n1258, new_n1259, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G244), .ZN(new_n215));
  AND2_X1   g0015(.A1(new_n215), .A2(G77), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G107), .A2(G264), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n205), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n208), .B(new_n214), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G68), .B(G77), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT66), .ZN(new_n235));
  XOR2_X1   g0035(.A(G50), .B(G58), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  INV_X1    g0041(.A(G1), .ZN(new_n242));
  NAND3_X1  g0042(.A1(new_n242), .A2(G13), .A3(G20), .ZN(new_n243));
  OR3_X1    g0043(.A1(new_n243), .A2(KEYINPUT12), .A3(G68), .ZN(new_n244));
  OAI21_X1  g0044(.A(KEYINPUT12), .B1(new_n243), .B2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n243), .A2(new_n211), .A3(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n242), .A2(G20), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(G68), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n247), .A2(new_n211), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  INV_X1    g0054(.A(G68), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n254), .A2(G77), .B1(G20), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT71), .ZN(new_n257));
  INV_X1    g0057(.A(G50), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n256), .A2(KEYINPUT71), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n252), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT11), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n246), .B(new_n251), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n263), .A2(new_n264), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT67), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n211), .ZN(new_n271));
  NAND3_X1  g0071(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(G274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n276), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n273), .A2(new_n278), .A3(G238), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G226), .A2(G1698), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(new_n226), .B2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n253), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n281), .A2(new_n285), .B1(G33), .B2(G97), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n271), .A2(new_n268), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n277), .B(new_n279), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT13), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  OAI21_X1  g0091(.A(KEYINPUT14), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(G179), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT14), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(KEYINPUT13), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n288), .A2(KEYINPUT13), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n294), .B(G169), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n292), .A2(new_n293), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT72), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n292), .A2(KEYINPUT72), .A3(new_n298), .A4(new_n293), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n267), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G1698), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n285), .A2(G232), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n285), .A2(G238), .A3(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(G107), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(new_n285), .ZN(new_n308));
  INV_X1    g0108(.A(new_n287), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n211), .B1(new_n269), .B2(new_n268), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n276), .B1(new_n311), .B2(new_n272), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n215), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(new_n277), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n250), .A2(G77), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n248), .A2(new_n317), .B1(G77), .B2(new_n243), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G20), .A2(G77), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT8), .B(G58), .ZN(new_n320));
  INV_X1    g0120(.A(new_n254), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT15), .B(G87), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n319), .B1(new_n320), .B2(new_n260), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n318), .B1(new_n323), .B2(new_n252), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n314), .A2(G200), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT70), .B(G179), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n314), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n324), .B1(new_n314), .B2(new_n291), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n326), .A2(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n252), .ZN(new_n333));
  INV_X1    g0133(.A(G58), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n334), .A2(KEYINPUT8), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n334), .A2(KEYINPUT8), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT68), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT68), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n320), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n339), .A3(new_n254), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n258), .A2(new_n334), .A3(new_n255), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(G20), .B1(G150), .B2(new_n259), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n333), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n250), .A2(G50), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT69), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n250), .A2(KEYINPUT69), .A3(G50), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n249), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G50), .B2(new_n243), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n285), .A2(G222), .A3(new_n304), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n285), .A2(G223), .A3(G1698), .ZN(new_n352));
  INV_X1    g0152(.A(G77), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n351), .B(new_n352), .C1(new_n353), .C2(new_n285), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n309), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n312), .A2(G226), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n277), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n350), .B1(new_n357), .B2(new_n291), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n329), .B2(new_n357), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT10), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(G200), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT9), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n343), .B2(new_n349), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n350), .A2(KEYINPUT9), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n355), .A2(G190), .A3(new_n277), .A4(new_n356), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n360), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n361), .A2(new_n365), .A3(new_n363), .A4(new_n366), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(KEYINPUT10), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n332), .B(new_n359), .C1(new_n368), .C2(new_n370), .ZN(new_n371));
  OR2_X1    g0171(.A1(G223), .A2(G1698), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(G226), .B2(new_n304), .ZN(new_n373));
  AND2_X1   g0173(.A1(KEYINPUT3), .A2(G33), .ZN(new_n374));
  NOR2_X1   g0174(.A1(KEYINPUT3), .A2(G33), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G87), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n373), .A2(new_n376), .B1(new_n253), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n309), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n312), .A2(G232), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n379), .A2(new_n315), .A3(new_n380), .A4(new_n277), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(KEYINPUT76), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n381), .A2(KEYINPUT76), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n379), .A2(new_n277), .A3(new_n380), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n382), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n283), .A2(new_n212), .A3(new_n284), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT74), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n283), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n284), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n392), .A2(new_n391), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(G68), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n334), .A2(new_n255), .ZN(new_n396));
  NOR2_X1   g0196(.A1(G58), .A2(G68), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n259), .A2(G159), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n390), .A2(new_n392), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n400), .B1(new_n405), .B2(G68), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n333), .B1(new_n406), .B2(KEYINPUT16), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n337), .A2(new_n339), .A3(new_n250), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n248), .B1(new_n409), .B2(KEYINPUT75), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT75), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n337), .A2(new_n339), .A3(new_n411), .A4(new_n250), .ZN(new_n412));
  INV_X1    g0212(.A(new_n243), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n337), .A2(new_n339), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n410), .A2(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n387), .A2(KEYINPUT17), .A3(new_n408), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n405), .A2(G68), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n401), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n252), .ZN(new_n419));
  INV_X1    g0219(.A(new_n403), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n395), .B2(new_n401), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n415), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n384), .A2(G169), .ZN(new_n423));
  INV_X1    g0223(.A(G274), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n311), .B2(new_n272), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n378), .A2(new_n309), .B1(new_n425), .B2(new_n276), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(new_n329), .A3(new_n380), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT18), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n422), .A2(new_n431), .A3(new_n428), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT76), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n426), .A2(new_n434), .A3(new_n315), .A4(new_n380), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n381), .A2(KEYINPUT76), .ZN(new_n436));
  AOI21_X1  g0236(.A(G200), .B1(new_n426), .B2(new_n380), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n433), .B1(new_n422), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n416), .A2(new_n430), .A3(new_n432), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n290), .A2(G190), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n267), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n290), .A2(new_n385), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR4_X1   g0244(.A1(new_n303), .A2(new_n371), .A3(new_n440), .A4(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(G257), .B(G1698), .C1(new_n374), .C2(new_n375), .ZN(new_n446));
  OAI211_X1 g0246(.A(G250), .B(new_n304), .C1(new_n374), .C2(new_n375), .ZN(new_n447));
  INV_X1    g0247(.A(G294), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n446), .B(new_n447), .C1(new_n253), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n309), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n275), .A2(G1), .ZN(new_n451));
  OR2_X1    g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  NAND2_X1  g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n273), .A2(G274), .A3(new_n451), .A4(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n453), .ZN(new_n456));
  NOR2_X1   g0256(.A1(KEYINPUT5), .A2(G41), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n451), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n273), .A2(new_n458), .A3(G264), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n450), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT83), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT83), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n450), .A2(new_n462), .A3(new_n455), .A4(new_n459), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(G169), .A3(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n273), .A2(new_n458), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n309), .A2(new_n449), .B1(new_n465), .B2(G264), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(G179), .A3(new_n455), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT82), .B1(new_n212), .B2(G107), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT23), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT23), .ZN(new_n470));
  OAI211_X1 g0270(.A(KEYINPUT82), .B(new_n470), .C1(new_n212), .C2(G107), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n469), .A2(new_n471), .B1(G116), .B2(new_n254), .ZN(new_n472));
  AOI21_X1  g0272(.A(G20), .B1(new_n283), .B2(new_n284), .ZN(new_n473));
  AND2_X1   g0273(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(G87), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n212), .B(G87), .C1(new_n374), .C2(new_n375), .ZN(new_n476));
  NOR2_X1   g0276(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n472), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n480), .A2(KEYINPUT24), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(KEYINPUT24), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n252), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n242), .A2(G33), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT77), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n484), .B(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n248), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT25), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n243), .B2(G107), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n413), .A2(KEYINPUT25), .A3(new_n307), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n487), .A2(G107), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n464), .A2(new_n467), .B1(new_n483), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n483), .A2(new_n491), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n462), .B1(new_n466), .B2(new_n455), .ZN(new_n495));
  INV_X1    g0295(.A(new_n463), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n315), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n460), .A2(new_n385), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n492), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(G250), .B(G1698), .C1(new_n374), .C2(new_n375), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  OAI211_X1 g0302(.A(G244), .B(new_n304), .C1(new_n374), .C2(new_n375), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT4), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n501), .B(new_n502), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  XOR2_X1   g0305(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n506));
  AND2_X1   g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n309), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n273), .A2(new_n458), .A3(G257), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n455), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n508), .A2(new_n328), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(G169), .B1(new_n508), .B2(new_n510), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n393), .A2(G107), .A3(new_n394), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT6), .ZN(new_n515));
  INV_X1    g0315(.A(G97), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n307), .ZN(new_n517));
  NOR2_X1   g0317(.A1(G97), .A2(G107), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n307), .A2(KEYINPUT6), .A3(G97), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n252), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n243), .A2(G97), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n484), .B(KEYINPUT77), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n249), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n528), .B2(new_n516), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n513), .A2(new_n531), .A3(KEYINPUT79), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT79), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n508), .A2(new_n328), .A3(new_n510), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n455), .A2(new_n509), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n503), .A2(new_n506), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n304), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n536), .A2(new_n537), .A3(new_n501), .A4(new_n502), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n535), .B1(new_n538), .B2(new_n309), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n534), .B1(new_n539), .B2(G169), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n529), .B1(new_n523), .B2(new_n252), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n533), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n508), .A2(new_n510), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n541), .B(new_n544), .C1(new_n315), .C2(new_n543), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n532), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n285), .A2(G264), .A3(G1698), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n285), .A2(G257), .A3(new_n304), .ZN(new_n548));
  INV_X1    g0348(.A(G303), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n547), .B(new_n548), .C1(new_n549), .C2(new_n285), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n309), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n273), .A2(new_n458), .A3(G270), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n455), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n527), .A2(G116), .A3(new_n249), .ZN(new_n555));
  INV_X1    g0355(.A(G116), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n413), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n247), .A2(new_n211), .B1(G20), .B2(new_n556), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n502), .B(new_n212), .C1(G33), .C2(new_n516), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT20), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n558), .A2(KEYINPUT20), .A3(new_n559), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n555), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n554), .A2(KEYINPUT21), .A3(G169), .A4(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n562), .A2(G179), .A3(new_n551), .A4(new_n553), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n291), .B1(new_n551), .B2(new_n553), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT21), .B1(new_n566), .B2(new_n562), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n254), .A2(G97), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT19), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n473), .A2(G68), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n212), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT80), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT80), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n575), .A3(new_n212), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n377), .A2(new_n516), .A3(new_n307), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n333), .B1(new_n571), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n322), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(new_n243), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n486), .A2(new_n377), .A3(new_n248), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(G244), .B(G1698), .C1(new_n374), .C2(new_n375), .ZN(new_n584));
  OAI211_X1 g0384(.A(G238), .B(new_n304), .C1(new_n374), .C2(new_n375), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(new_n585), .C1(new_n253), .C2(new_n556), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n309), .ZN(new_n587));
  AOI21_X1  g0387(.A(G250), .B1(new_n242), .B2(G45), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n424), .B2(new_n451), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n273), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(G190), .A3(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n586), .A2(new_n309), .B1(new_n273), .B2(new_n589), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n583), .B(new_n591), .C1(new_n385), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n571), .A2(new_n578), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n252), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n487), .A2(new_n580), .ZN(new_n596));
  INV_X1    g0396(.A(new_n581), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n587), .A2(new_n590), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n291), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n592), .A2(new_n328), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n562), .B1(new_n554), .B2(G200), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n315), .B2(new_n554), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n568), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n445), .A2(new_n500), .A3(new_n546), .A4(new_n606), .ZN(G372));
  INV_X1    g0407(.A(new_n359), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n416), .A2(new_n439), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n301), .A2(new_n302), .ZN(new_n610));
  INV_X1    g0410(.A(new_n267), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n444), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n330), .A2(new_n331), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n609), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n430), .A2(new_n432), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT85), .ZN(new_n620));
  INV_X1    g0420(.A(new_n368), .ZN(new_n621));
  INV_X1    g0421(.A(new_n370), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n619), .A2(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OR3_X1    g0423(.A1(new_n617), .A2(new_n620), .A3(new_n618), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n608), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n464), .A2(new_n467), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n493), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n568), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT84), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n599), .A2(new_n629), .A3(G200), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT84), .B1(new_n592), .B2(new_n385), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n582), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n591), .A2(new_n597), .A3(new_n595), .A4(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n602), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n499), .B2(new_n494), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n546), .A2(new_n628), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n532), .A2(new_n542), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n640), .B2(new_n603), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n630), .A2(new_n631), .A3(new_n583), .A4(new_n591), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n642), .A2(new_n513), .A3(new_n531), .A4(new_n602), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n602), .B1(new_n643), .B2(KEYINPUT26), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n445), .B1(new_n638), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n625), .A2(new_n647), .ZN(G369));
  NAND2_X1  g0448(.A1(new_n566), .A2(new_n562), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT21), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n651), .A2(new_n564), .A3(new_n563), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n242), .A2(new_n212), .A3(G13), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n653), .A2(KEYINPUT86), .A3(KEYINPUT27), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT86), .B1(new_n653), .B2(KEYINPUT27), .ZN(new_n655));
  OAI221_X1 g0455(.A(G213), .B1(KEYINPUT27), .B2(new_n653), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(new_n562), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n605), .A2(new_n651), .A3(new_n564), .A4(new_n563), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n659), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n658), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n500), .B1(new_n494), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n492), .A2(new_n658), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n652), .A2(new_n665), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n500), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n492), .A2(new_n665), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n669), .A2(new_n674), .ZN(G399));
  INV_X1    g0475(.A(new_n206), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n577), .A2(G116), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G1), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n209), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n543), .A2(new_n460), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n592), .A2(new_n329), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n554), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT87), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT87), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n554), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n683), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n539), .A2(new_n466), .A3(new_n592), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n551), .A2(new_n553), .A3(G179), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n692), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n466), .A2(new_n592), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(KEYINPUT30), .A4(new_n539), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n658), .B1(new_n689), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT31), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n606), .A2(new_n500), .A3(new_n546), .A4(new_n665), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n699), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT89), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n637), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n546), .A2(new_n628), .A3(new_n636), .A4(KEYINPUT89), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT79), .B1(new_n513), .B2(new_n531), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n540), .A2(new_n541), .A3(new_n533), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n603), .B(new_n639), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n602), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n643), .B2(KEYINPUT26), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n707), .A2(new_n708), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(KEYINPUT29), .A3(new_n665), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT90), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n715), .A2(KEYINPUT90), .A3(KEYINPUT29), .A4(new_n665), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n658), .B1(new_n645), .B2(new_n637), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  XOR2_X1   g0522(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n705), .B1(new_n720), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n682), .B1(new_n726), .B2(G1), .ZN(G364));
  AND2_X1   g0527(.A1(new_n212), .A2(G13), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n242), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n677), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n664), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(G330), .B2(new_n662), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n285), .A2(new_n206), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n203), .A2(new_n734), .B1(G116), .B2(new_n206), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n376), .A2(new_n206), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT91), .Z(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n275), .B2(new_n210), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n237), .A2(G45), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n735), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT92), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n211), .B1(G20), .B2(new_n291), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n731), .B1(new_n741), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n212), .A2(new_n385), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n329), .A2(new_n315), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT95), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n752), .B(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(KEYINPUT33), .B(G317), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n212), .A2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(G179), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n757), .A2(new_n758), .A3(G200), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT94), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n212), .A2(new_n315), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n329), .A2(new_n385), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n763), .A2(G283), .B1(G322), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n757), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G329), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n764), .A2(new_n758), .A3(G200), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n376), .B1(new_n769), .B2(new_n770), .C1(new_n771), .C2(new_n549), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n768), .A2(G190), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n772), .B1(G294), .B2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n328), .A2(new_n212), .A3(new_n385), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n776), .A2(G190), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n329), .A2(new_n385), .A3(new_n757), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n777), .A2(G326), .B1(new_n779), .B2(G311), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n756), .A2(new_n767), .A3(new_n775), .A4(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n777), .A2(G50), .B1(new_n766), .B2(G58), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(new_n353), .B2(new_n778), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  INV_X1    g0584(.A(new_n774), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n516), .ZN(new_n786));
  INV_X1    g0586(.A(new_n771), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G87), .ZN(new_n788));
  INV_X1    g0588(.A(new_n769), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G159), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n788), .B(new_n285), .C1(KEYINPUT32), .C2(new_n790), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n786), .B(new_n791), .C1(KEYINPUT32), .C2(new_n790), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n763), .A2(G107), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n752), .B(KEYINPUT95), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n792), .B(new_n793), .C1(new_n255), .C2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n781), .B1(new_n784), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n750), .B1(new_n796), .B2(new_n747), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n662), .B2(new_n745), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n733), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  OR2_X1    g0600(.A1(new_n614), .A2(KEYINPUT99), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n326), .A2(new_n327), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n614), .A2(KEYINPUT99), .ZN(new_n803));
  AND3_X1   g0603(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n721), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n665), .A2(new_n324), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n801), .A2(new_n802), .A3(new_n807), .A4(new_n803), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n615), .A2(new_n658), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n805), .B1(new_n721), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n704), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT100), .Z(new_n813));
  AOI21_X1  g0613(.A(new_n731), .B1(new_n811), .B2(new_n704), .ZN(new_n814));
  INV_X1    g0614(.A(new_n810), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n742), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n747), .A2(new_n742), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n763), .A2(G87), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n820), .B2(new_n769), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT97), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n285), .B(new_n786), .C1(G107), .C2(new_n787), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n556), .B2(new_n778), .ZN(new_n824));
  INV_X1    g0624(.A(new_n777), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n825), .A2(new_n549), .B1(new_n448), .B2(new_n765), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n822), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n794), .A2(KEYINPUT96), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT96), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n754), .A2(new_n829), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G283), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n777), .A2(G137), .B1(new_n779), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  INV_X1    g0634(.A(G150), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n834), .B2(new_n765), .C1(new_n794), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n763), .A2(G68), .ZN(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n285), .B1(new_n769), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G50), .B2(new_n787), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n839), .B(new_n842), .C1(new_n334), .C2(new_n785), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n836), .B2(new_n837), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n827), .A2(new_n832), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n747), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n731), .B1(G77), .B2(new_n818), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT98), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n813), .A2(new_n814), .B1(new_n816), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  OR2_X1    g0650(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n851), .A2(G116), .A3(new_n213), .A4(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT36), .Z(new_n854));
  OAI211_X1 g0654(.A(new_n210), .B(G77), .C1(new_n334), .C2(new_n255), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n258), .A2(G68), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n242), .B(G13), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n658), .B1(new_n801), .B2(new_n803), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n721), .B2(new_n804), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n267), .A2(new_n665), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n612), .B2(new_n613), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n303), .A2(new_n444), .A3(new_n861), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n407), .B1(new_n420), .B2(new_n406), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n656), .B1(new_n867), .B2(new_n415), .ZN(new_n868));
  INV_X1    g0668(.A(new_n428), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n869), .A2(new_n656), .B1(new_n867), .B2(new_n415), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n422), .A2(new_n438), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n386), .A2(KEYINPUT76), .A3(new_n381), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n408), .A2(new_n873), .A3(new_n415), .A4(new_n435), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n656), .B(KEYINPUT101), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n422), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n874), .A2(new_n429), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n440), .A2(new_n868), .B1(new_n872), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(KEYINPUT38), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n875), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n866), .A2(new_n883), .B1(new_n618), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n876), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n440), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n874), .A2(new_n429), .A3(new_n876), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n878), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT102), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT102), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n440), .A2(new_n886), .B1(new_n889), .B2(new_n878), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n893), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(new_n895), .A3(new_n882), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n612), .A2(new_n658), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n885), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT104), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n619), .A2(new_n620), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n621), .A2(new_n622), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(new_n624), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n359), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n445), .B1(new_n721), .B2(new_n723), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n720), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT103), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n720), .A2(KEYINPUT103), .A3(new_n909), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n907), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n903), .B(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n896), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n612), .A2(new_n613), .A3(new_n862), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n861), .B1(new_n303), .B2(new_n444), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n815), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n702), .A2(KEYINPUT105), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT105), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n698), .A2(new_n921), .A3(new_n699), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n920), .A2(new_n700), .A3(new_n701), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT40), .B1(new_n916), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT40), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n883), .A2(new_n919), .A3(new_n926), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n445), .A2(new_n923), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT106), .Z(new_n930));
  OAI21_X1  g0730(.A(G330), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n931), .A2(KEYINPUT107), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n928), .A2(new_n930), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(KEYINPUT107), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n915), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n242), .B2(new_n728), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n915), .A2(new_n935), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n858), .B1(new_n937), .B2(new_n938), .ZN(G367));
  OAI21_X1  g0739(.A(new_n546), .B1(new_n541), .B2(new_n665), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n513), .A2(new_n531), .A3(new_n658), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n672), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT42), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n940), .A2(new_n941), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n627), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n665), .B1(new_n948), .B2(new_n640), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n665), .A2(new_n583), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n712), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n635), .B2(new_n950), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n946), .A2(new_n949), .B1(KEYINPUT43), .B2(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n669), .A2(new_n947), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n677), .B(KEYINPUT41), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n711), .A2(new_n713), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n706), .B2(new_n637), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n658), .B1(new_n960), .B2(new_n708), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT90), .B1(new_n961), .B2(KEYINPUT29), .ZN(new_n962));
  INV_X1    g0762(.A(new_n719), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n725), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n965), .A2(new_n663), .A3(new_n672), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n663), .B1(new_n965), .B2(new_n672), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n964), .A2(new_n704), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(KEYINPUT108), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT108), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n726), .A2(new_n972), .A3(new_n969), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n674), .B2(new_n942), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n672), .A2(new_n673), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n947), .A2(new_n976), .A3(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT45), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n947), .B2(new_n976), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n674), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n978), .A2(new_n982), .A3(new_n669), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n669), .B1(new_n978), .B2(new_n982), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n971), .A2(new_n973), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n958), .B1(new_n987), .B2(new_n726), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n957), .B1(new_n988), .B2(new_n730), .ZN(new_n989));
  INV_X1    g0789(.A(new_n731), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n748), .B1(new_n206), .B2(new_n322), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n232), .B2(new_n737), .ZN(new_n992));
  INV_X1    g0792(.A(G137), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n285), .B1(new_n769), .B2(new_n993), .C1(new_n771), .C2(new_n334), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n777), .A2(G143), .B1(new_n779), .B2(G50), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n763), .A2(G77), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(new_n835), .C2(new_n765), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n994), .B(new_n997), .C1(G68), .C2(new_n774), .ZN(new_n998));
  INV_X1    g0798(.A(G159), .ZN(new_n999));
  INV_X1    g0799(.A(new_n831), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n766), .A2(G303), .B1(new_n779), .B2(G283), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n763), .A2(G97), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(new_n820), .C2(new_n825), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n285), .B1(new_n789), .B2(G317), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n771), .A2(new_n556), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(KEYINPUT46), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(KEYINPUT46), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n307), .B2(new_n785), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n1004), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n1000), .B2(new_n448), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1001), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT47), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n990), .B(new_n992), .C1(new_n1013), .C2(new_n747), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT109), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n745), .B2(new_n952), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT110), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n989), .A2(new_n1017), .ZN(G387));
  NAND3_X1  g0818(.A1(new_n666), .A2(new_n667), .A3(new_n746), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n229), .A2(G45), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT111), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n320), .A2(G50), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT50), .Z(new_n1023));
  OAI211_X1 g0823(.A(new_n679), .B(new_n275), .C1(new_n255), .C2(new_n353), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n737), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(G107), .B2(new_n206), .C1(new_n679), .C2(new_n734), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n990), .B1(new_n1026), .B2(new_n748), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n777), .A2(G159), .B1(new_n779), .B2(G68), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1028), .B(new_n1003), .C1(new_n258), .C2(new_n765), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n794), .A2(new_n414), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n376), .B1(new_n789), .B2(G150), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n787), .A2(G77), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n322), .C2(new_n785), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n777), .A2(G322), .B1(new_n766), .B2(G317), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n549), .B2(new_n778), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n831), .B2(G311), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT48), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(KEYINPUT48), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n787), .A2(G294), .B1(new_n774), .B2(G283), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT49), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n763), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(new_n556), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n285), .B(new_n1044), .C1(G326), .C2(new_n789), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1034), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1019), .B(new_n1027), .C1(new_n1046), .C2(new_n846), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT112), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n968), .A2(new_n729), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n718), .A2(new_n719), .B1(new_n722), .B2(new_n724), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n968), .B1(new_n1051), .B2(new_n705), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n972), .B1(new_n726), .B2(new_n969), .ZN(new_n1053));
  NOR4_X1   g0853(.A1(new_n1051), .A2(KEYINPUT108), .A3(new_n705), .A4(new_n968), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n677), .B(new_n1052), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1050), .A2(new_n1055), .ZN(G393));
  OAI22_X1  g0856(.A1(new_n1053), .A2(new_n1054), .B1(new_n984), .B2(new_n985), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(new_n677), .A3(new_n987), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n978), .A2(new_n982), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n669), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(new_n730), .A3(new_n983), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n749), .B1(G97), .B2(new_n676), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n737), .A2(new_n240), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n990), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n777), .A2(G317), .B1(new_n766), .B2(G311), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT114), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT52), .Z(new_n1068));
  AOI21_X1  g0868(.A(new_n285), .B1(new_n787), .B2(G283), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n789), .A2(G322), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(new_n556), .C2(new_n785), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n793), .B1(new_n448), .B2(new_n778), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n831), .C2(G303), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n777), .A2(G150), .B1(new_n766), .B2(G159), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT51), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n785), .A2(new_n353), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n819), .B1(new_n320), .B2(new_n778), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n285), .B1(new_n769), .B2(new_n834), .C1(new_n771), .C2(new_n255), .ZN(new_n1078));
  NOR4_X1   g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n831), .A2(G50), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1068), .A2(new_n1073), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n947), .A2(new_n746), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1082), .A2(KEYINPUT113), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(KEYINPUT113), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1065), .B1(new_n846), .B2(new_n1081), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n1062), .A2(KEYINPUT115), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT115), .B1(new_n1062), .B2(new_n1085), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1058), .A2(new_n1089), .ZN(G390));
  AND2_X1   g0890(.A1(new_n923), .A2(G330), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n445), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT103), .B1(new_n720), .B2(new_n909), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n911), .B(new_n908), .C1(new_n718), .C2(new_n719), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n625), .B(new_n1092), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n899), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n860), .B2(new_n865), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n891), .A2(KEYINPUT102), .B1(KEYINPUT38), .B2(new_n879), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n1099), .B2(new_n895), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n882), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1101), .A2(new_n880), .A3(new_n897), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1098), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT116), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n919), .A2(new_n1104), .A3(G330), .A4(new_n923), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n703), .A2(G330), .A3(new_n810), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n865), .A2(new_n1106), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n715), .A2(new_n665), .A3(new_n804), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n859), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n917), .A2(new_n918), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n899), .B1(new_n1099), .B2(new_n895), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1103), .A2(new_n1108), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n898), .A2(new_n900), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1117), .A2(new_n1098), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1091), .A2(new_n919), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n1104), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1116), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1091), .A2(new_n810), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n865), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n865), .A2(new_n1106), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n860), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1096), .A2(new_n1121), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1120), .B1(new_n1103), .B2(new_n1115), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n860), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1116), .C1(new_n1095), .C2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1129), .A2(new_n1134), .A3(new_n677), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n743), .B1(new_n898), .B2(new_n900), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n990), .B1(new_n414), .B2(new_n817), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1076), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n789), .A2(G294), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1138), .A2(new_n376), .A3(new_n788), .A4(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n777), .A2(G283), .B1(new_n779), .B2(G97), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1141), .B(new_n839), .C1(new_n556), .C2(new_n765), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(new_n831), .C2(G107), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT54), .B(G143), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n1000), .A2(new_n993), .B1(new_n778), .B2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT117), .Z(new_n1146));
  NOR2_X1   g0946(.A1(new_n771), .A2(new_n835), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT53), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n376), .B1(new_n789), .B2(G125), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(new_n999), .C2(new_n785), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1043), .A2(new_n258), .B1(new_n840), .B2(new_n765), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G128), .C2(new_n777), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1143), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1137), .B1(new_n1153), .B2(new_n846), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1136), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n1121), .B2(new_n730), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1135), .A2(new_n1156), .ZN(G378));
  INV_X1    g0957(.A(G330), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n925), .B2(new_n927), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n905), .A2(new_n359), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n350), .A2(new_n656), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1161), .B(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n885), .A2(new_n901), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(new_n885), .B2(new_n901), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1160), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1166), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1100), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n805), .A2(new_n1110), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(new_n883), .A3(new_n1112), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n618), .A2(new_n884), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1171), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n1159), .A3(new_n1167), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1170), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1171), .A2(new_n742), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n731), .B1(G50), .B2(new_n818), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT121), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n789), .A2(G283), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n285), .A2(G41), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1032), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n763), .A2(G58), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n307), .B2(new_n765), .C1(new_n556), .C2(new_n825), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G68), .C2(new_n774), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n754), .A2(G97), .B1(new_n580), .B2(new_n779), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT119), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1188), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1194));
  OR2_X1    g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G50), .B(new_n1184), .C1(new_n253), .C2(new_n274), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT118), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n777), .A2(G125), .B1(new_n766), .B2(G128), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n785), .A2(new_n835), .B1(new_n1144), .B2(new_n771), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G137), .B2(new_n779), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1199), .B(new_n1201), .C1(new_n794), .C2(new_n840), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n789), .C2(G124), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1043), .B2(new_n999), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n1202), .B2(KEYINPUT59), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1198), .B1(new_n1203), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1195), .A2(new_n1196), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1182), .B1(new_n1208), .B2(new_n747), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1179), .A2(new_n730), .B1(new_n1180), .B2(new_n1209), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1177), .A2(new_n1159), .A3(new_n1167), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1159), .B1(new_n1177), .B2(new_n1167), .ZN(new_n1212));
  OAI21_X1  g1012(.A(KEYINPUT57), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1095), .B1(new_n1121), .B2(new_n1128), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n677), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1108), .A2(new_n1103), .A3(new_n1115), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1216), .A2(new_n1130), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1096), .B1(new_n1217), .B2(new_n1133), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT57), .B1(new_n1218), .B2(new_n1179), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1210), .B1(new_n1215), .B2(new_n1219), .ZN(G375));
  NAND3_X1  g1020(.A1(new_n914), .A2(new_n1092), .A3(new_n1128), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n958), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1095), .A2(new_n1133), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n865), .A2(new_n742), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n731), .B1(G68), .B2(new_n818), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1000), .A2(new_n556), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n777), .A2(G294), .B1(new_n766), .B2(G283), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n376), .B1(new_n769), .B2(new_n549), .C1(new_n771), .C2(new_n516), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n580), .B2(new_n774), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n779), .A2(G107), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1230), .A3(new_n996), .A4(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1000), .A2(new_n1144), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n376), .B1(new_n789), .B2(G128), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n999), .B2(new_n771), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G50), .B2(new_n774), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n779), .A2(G150), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n777), .A2(G132), .B1(new_n766), .B2(G137), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1236), .A2(new_n1186), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1227), .A2(new_n1232), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1226), .B1(new_n1240), .B2(new_n747), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1128), .A2(new_n730), .B1(new_n1225), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1224), .A2(new_n1242), .ZN(G381));
  NAND3_X1  g1043(.A1(new_n1050), .A2(new_n799), .A3(new_n1055), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n849), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT122), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n678), .B1(new_n1248), .B2(new_n986), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1088), .B1(new_n1249), .B2(new_n1057), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n989), .A2(new_n1250), .A3(new_n1017), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1217), .A2(new_n729), .B1(new_n1136), .B2(new_n1154), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n678), .B1(new_n1221), .B2(new_n1217), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(new_n1253), .B2(new_n1129), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n1242), .A3(new_n1224), .ZN(new_n1255));
  OR4_X1    g1055(.A1(G375), .A2(new_n1247), .A3(new_n1251), .A4(new_n1255), .ZN(G407));
  NAND2_X1  g1056(.A1(new_n657), .A2(G213), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(G375), .A2(G378), .A3(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT123), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(G407), .A2(G213), .A3(new_n1259), .ZN(G409));
  AOI21_X1  g1060(.A(new_n799), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1244), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT127), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n989), .B2(new_n1017), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1265), .B2(new_n1250), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1264), .B(G390), .C1(new_n989), .C2(new_n1017), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT126), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1245), .B2(new_n1261), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1262), .A2(KEYINPUT126), .A3(new_n1244), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1251), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1250), .B1(new_n1017), .B2(new_n989), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n1266), .A2(new_n1267), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G378), .B(new_n1210), .C1(new_n1215), .C2(new_n1219), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1277), .A2(new_n1214), .A3(new_n958), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1180), .A2(new_n1209), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1277), .B2(new_n729), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1254), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1276), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1242), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n677), .B1(new_n1095), .B2(new_n1133), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT60), .B1(new_n1095), .B2(new_n1133), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1095), .A2(KEYINPUT60), .A3(new_n1133), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n849), .B(new_n1283), .C1(new_n1286), .C2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1223), .A2(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1290), .A2(new_n677), .A3(new_n1221), .A4(new_n1287), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G384), .B1(new_n1291), .B2(new_n1242), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1293));
  AND4_X1   g1093(.A1(KEYINPUT63), .A2(new_n1282), .A3(new_n1257), .A4(new_n1293), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1276), .A2(new_n1281), .B1(G213), .B2(new_n657), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT63), .B1(new_n1295), .B2(new_n1293), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1275), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1282), .A2(new_n1257), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n657), .A2(G213), .A3(G2897), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1299), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT124), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1287), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1302), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n849), .B1(new_n1303), .B2(new_n1283), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1291), .A2(G384), .A3(new_n1242), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1299), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1300), .A2(new_n1301), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1301), .B1(new_n1300), .B2(new_n1307), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1298), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT125), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT125), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1312), .B(new_n1298), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1297), .A2(new_n1311), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1273), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1293), .ZN(new_n1316));
  OAI21_X1  g1116(.A(KEYINPUT62), .B1(new_n1298), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1300), .A2(new_n1307), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT61), .B1(new_n1298), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(new_n1298), .A2(KEYINPUT62), .A3(new_n1316), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1315), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1314), .A2(new_n1322), .ZN(G405));
  NAND2_X1  g1123(.A1(G375), .A2(new_n1254), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1276), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1325), .B(new_n1293), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n1315), .ZN(G402));
endmodule


