//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n892, new_n893, new_n895, new_n896, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947;
  OR3_X1    g000(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(G148gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G141gat), .ZN(new_n205));
  INV_X1    g004(.A(G141gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G148gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n202), .A2(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n207), .ZN(new_n209));
  AND2_X1   g008(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n210));
  NOR2_X1   g009(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n209), .A2(new_n212), .B1(G155gat), .B2(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(G155gat), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n208), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G113gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT67), .A3(G120gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(G127gat), .A2(G134gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G127gat), .A2(G134gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G120gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G113gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n218), .A2(G120gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n228), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n220), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n225), .A2(new_n230), .B1(new_n232), .B2(new_n224), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT73), .B1(new_n217), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G141gat), .B(G148gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT72), .B(KEYINPUT2), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n203), .B(new_n216), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n202), .A2(new_n203), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n209), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n230), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n219), .B(new_n220), .C1(new_n223), .C2(new_n222), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT1), .B1(new_n227), .B2(new_n228), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n222), .A2(new_n223), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n241), .A2(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT73), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n240), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT4), .B1(new_n234), .B2(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n240), .A2(new_n245), .A3(KEYINPUT4), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(KEYINPUT75), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n217), .A2(KEYINPUT73), .A3(new_n233), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n246), .B1(new_n240), .B2(new_n245), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n252), .B1(new_n256), .B2(new_n249), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT5), .ZN(new_n259));
  NAND2_X1  g058(.A1(G225gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n217), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n240), .A2(KEYINPUT3), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n245), .A3(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n258), .A2(new_n259), .A3(new_n260), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT76), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n254), .A2(new_n255), .B1(new_n245), .B2(new_n240), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT5), .B1(new_n267), .B2(new_n260), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n268), .A2(KEYINPUT74), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(KEYINPUT74), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n253), .B1(new_n234), .B2(new_n247), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n240), .A2(new_n245), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT4), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n271), .A2(new_n260), .A3(new_n264), .A4(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n269), .A2(new_n270), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n264), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n276), .B1(new_n251), .B2(new_n257), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT76), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n259), .A4(new_n260), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n266), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281));
  INV_X1    g080(.A(G85gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT0), .B(G57gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n283), .B(new_n284), .Z(new_n285));
  NAND2_X1  g084(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n287));
  INV_X1    g086(.A(new_n285), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n266), .A2(new_n275), .A3(new_n288), .A4(new_n279), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT82), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT82), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n286), .A2(new_n292), .A3(new_n287), .A4(new_n289), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n280), .A2(KEYINPUT6), .A3(new_n285), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT38), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G211gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT22), .ZN(new_n301));
  AND2_X1   g100(.A1(KEYINPUT69), .A2(G218gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(KEYINPUT69), .A2(G218gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n300), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G204gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G197gat), .ZN(new_n308));
  INV_X1    g107(.A(G197gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G204gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n311), .A2(new_n301), .A3(G211gat), .ZN(new_n312));
  OAI21_X1  g111(.A(G218gat), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(KEYINPUT69), .A2(G218gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(KEYINPUT69), .A2(G218gat), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT22), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(G211gat), .B1(new_n316), .B2(new_n311), .ZN(new_n317));
  INV_X1    g116(.A(G218gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n305), .A2(KEYINPUT22), .A3(new_n300), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322));
  AND2_X1   g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(KEYINPUT23), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n322), .B1(new_n325), .B2(KEYINPUT65), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n324), .A2(KEYINPUT23), .ZN(new_n327));
  INV_X1    g126(.A(G169gat), .ZN(new_n328));
  INV_X1    g127(.A(G176gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT23), .ZN(new_n330));
  NAND2_X1  g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT65), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n327), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT66), .ZN(new_n335));
  AND2_X1   g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(KEYINPUT24), .ZN(new_n337));
  INV_X1    g136(.A(G183gat), .ZN(new_n338));
  INV_X1    g137(.A(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(KEYINPUT24), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT66), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n337), .A2(new_n340), .A3(new_n341), .A4(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n334), .A3(new_n344), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n324), .A2(KEYINPUT23), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347));
  NAND2_X1  g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n340), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n325), .B(new_n346), .C1(new_n349), .C2(new_n342), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT27), .B(G183gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n339), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT28), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT26), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n331), .A2(new_n357), .ZN(new_n358));
  MUX2_X1   g157(.A(new_n358), .B(new_n357), .S(new_n324), .Z(new_n359));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n354), .A2(new_n360), .A3(new_n339), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n356), .A2(new_n359), .A3(new_n348), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G226gat), .A2(G233gat), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n353), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n353), .B2(new_n362), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n321), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n362), .A3(new_n363), .ZN(new_n370));
  INV_X1    g169(.A(new_n321), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n359), .A2(new_n348), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n356), .A2(new_n361), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n373), .A2(new_n374), .B1(new_n345), .B2(new_n352), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n370), .B(new_n371), .C1(new_n375), .C2(new_n367), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n369), .A2(KEYINPUT70), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n370), .B1(new_n375), .B2(new_n367), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT70), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n379), .A3(new_n321), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT37), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n382), .B1(new_n381), .B2(new_n383), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n296), .B(new_n299), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n388), .A3(new_n376), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n378), .A2(KEYINPUT83), .A3(new_n321), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(KEYINPUT37), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT85), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n299), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n381), .A2(new_n383), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT84), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n394), .B1(new_n396), .B2(new_n384), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT85), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n397), .A2(new_n391), .A3(new_n398), .A4(new_n296), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n299), .B1(new_n377), .B2(new_n380), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n397), .B1(new_n383), .B2(new_n381), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(KEYINPUT38), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n294), .A2(new_n295), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n401), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT30), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n377), .A2(new_n380), .A3(new_n299), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT71), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n401), .A2(new_n409), .A3(KEYINPUT30), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n401), .B2(KEYINPUT30), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n407), .B(new_n408), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n260), .B1(new_n258), .B2(new_n264), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT39), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n267), .A2(new_n260), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n416), .B(KEYINPUT39), .C1(new_n277), .C2(new_n260), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n417), .A3(new_n288), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT40), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n285), .B1(new_n413), .B2(new_n414), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(KEYINPUT40), .A3(new_n417), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n412), .A2(new_n286), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT81), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n421), .A2(KEYINPUT40), .A3(new_n417), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT40), .B1(new_n421), .B2(new_n417), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT81), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n286), .A4(new_n412), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n313), .A2(new_n320), .A3(new_n365), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n430), .A2(KEYINPUT77), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n313), .A2(new_n320), .A3(new_n432), .A4(new_n365), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n261), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n240), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(G228gat), .ZN(new_n436));
  INV_X1    g235(.A(G233gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n262), .A2(new_n365), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n321), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n440), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n217), .B1(new_n430), .B2(new_n261), .ZN(new_n445));
  OAI22_X1  g244(.A1(new_n444), .A2(new_n445), .B1(new_n436), .B2(new_n437), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n435), .A2(KEYINPUT78), .A3(new_n438), .A4(new_n440), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT80), .B1(new_n448), .B2(G22gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(G22gat), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n443), .A2(new_n451), .A3(new_n446), .A4(new_n447), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT79), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n448), .A2(KEYINPUT80), .A3(G22gat), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n450), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G78gat), .B(G106gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT31), .B(G50gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n448), .A2(G22gat), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(new_n460), .A3(new_n452), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n424), .A2(new_n429), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n404), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT68), .ZN(new_n467));
  XNOR2_X1  g266(.A(G15gat), .B(G43gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n468), .B(new_n469), .Z(new_n470));
  NAND2_X1  g269(.A1(G227gat), .A2(G233gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n375), .A2(new_n233), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n353), .A2(new_n362), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n245), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n470), .B1(new_n475), .B2(KEYINPUT33), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n472), .A2(new_n474), .ZN(new_n478));
  INV_X1    g277(.A(new_n471), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT34), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n472), .A2(new_n474), .A3(new_n481), .A4(new_n471), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n475), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n485), .A2(KEYINPUT32), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n476), .A2(new_n480), .A3(new_n482), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n486), .B1(new_n484), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n467), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n290), .A2(new_n295), .ZN(new_n493));
  INV_X1    g292(.A(new_n412), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n448), .A2(KEYINPUT80), .A3(G22gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n496), .A2(new_n449), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n452), .B(KEYINPUT79), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n460), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n464), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n492), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n466), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n294), .A2(new_n295), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(new_n462), .B2(new_n464), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n412), .A2(KEYINPUT35), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n505), .B1(new_n499), .B2(new_n500), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT35), .B1(new_n510), .B2(new_n495), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n503), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G43gat), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT15), .B1(new_n514), .B2(G50gat), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n514), .B2(G50gat), .ZN(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  INV_X1    g316(.A(G36gat), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NOR3_X1   g319(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n521));
  OAI221_X1 g320(.A(new_n516), .B1(new_n517), .B2(new_n518), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  OAI22_X1  g321(.A1(new_n520), .A2(new_n521), .B1(new_n517), .B2(new_n518), .ZN(new_n523));
  XOR2_X1   g322(.A(KEYINPUT87), .B(G50gat), .Z(new_n524));
  OAI21_X1  g323(.A(KEYINPUT88), .B1(new_n524), .B2(G43gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT87), .B(G50gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n527), .A3(new_n514), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n525), .B(new_n528), .C1(new_n514), .C2(G50gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT86), .B(KEYINPUT15), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n523), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n522), .B1(new_n531), .B2(new_n516), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT17), .ZN(new_n533));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534));
  INV_X1    g333(.A(G1gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT16), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(G1gat), .B2(new_n534), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(KEYINPUT90), .Z(new_n541));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n542), .B(new_n522), .C1(new_n531), .C2(new_n516), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT89), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n533), .B(new_n541), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n532), .A2(new_n540), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT18), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n540), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n532), .B(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n548), .B(KEYINPUT13), .ZN(new_n556));
  OR3_X1    g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n547), .A2(KEYINPUT18), .A3(new_n548), .A4(new_n549), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n552), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G113gat), .B(G141gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n309), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT11), .B(G169gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n565), .B(KEYINPUT12), .Z(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n566), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n552), .A2(new_n559), .A3(new_n560), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n543), .B(KEYINPUT89), .ZN(new_n573));
  NAND2_X1  g372(.A1(G99gat), .A2(G106gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT8), .A2(new_n574), .B1(new_n282), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(new_n282), .B2(new_n575), .ZN(new_n578));
  NAND3_X1  g377(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G99gat), .B(G106gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n533), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n573), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n532), .A2(new_n582), .ZN(new_n585));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n586), .B(KEYINPUT94), .Z(new_n587));
  INV_X1    g386(.A(KEYINPUT41), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n572), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n592));
  INV_X1    g391(.A(new_n590), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n593), .B(new_n571), .C1(new_n573), .C2(new_n583), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n587), .A2(new_n588), .ZN(new_n596));
  XOR2_X1   g395(.A(G134gat), .B(G162gat), .Z(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT9), .ZN(new_n601));
  INV_X1    g400(.A(G71gat), .ZN(new_n602));
  INV_X1    g401(.A(G78gat), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT92), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G71gat), .B(G78gat), .Z(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G57gat), .B(G64gat), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n605), .B2(new_n604), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n609), .A2(new_n601), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n607), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G127gat), .B(G155gat), .Z(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n608), .A2(new_n610), .B1(new_n612), .B2(new_n607), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT21), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n540), .A2(new_n621), .A3(new_n338), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n338), .B1(new_n540), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n622), .B2(new_n623), .ZN(new_n628));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n300), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n631), .B1(new_n626), .B2(new_n628), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n619), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n636), .A2(new_n618), .A3(new_n632), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n591), .A2(new_n594), .A3(new_n592), .A4(new_n598), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n580), .A2(new_n581), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n580), .A2(new_n581), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n644), .B(new_n620), .C1(KEYINPUT96), .C2(new_n643), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n643), .A2(KEYINPUT96), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n582), .B1(new_n614), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n644), .A2(KEYINPUT10), .A3(new_n620), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n641), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n645), .A2(new_n648), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n641), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n653), .B(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n600), .A2(new_n638), .A3(new_n639), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT97), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n513), .A2(new_n570), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n493), .B(KEYINPUT98), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n535), .ZN(G1324gat));
  NOR2_X1   g463(.A1(new_n660), .A2(new_n494), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT42), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(new_n539), .B2(new_n665), .ZN(G1325gat));
  NOR2_X1   g468(.A1(new_n660), .A2(new_n506), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(G15gat), .ZN(new_n671));
  INV_X1    g470(.A(new_n492), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n660), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(G15gat), .B2(new_n673), .ZN(G1326gat));
  INV_X1    g473(.A(new_n501), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT43), .B(G22gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  AOI22_X1  g477(.A1(new_n502), .A2(new_n466), .B1(new_n509), .B2(new_n511), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n600), .A2(new_n639), .ZN(new_n680));
  INV_X1    g479(.A(new_n570), .ZN(new_n681));
  INV_X1    g480(.A(new_n657), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n681), .A2(new_n638), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n679), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(new_n517), .A3(new_n661), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT45), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n600), .A2(new_n639), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n513), .B2(new_n689), .ZN(new_n690));
  AOI211_X1 g489(.A(KEYINPUT44), .B(new_n680), .C1(new_n503), .C2(new_n512), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n683), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT99), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT44), .B1(new_n679), .B2(new_n680), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n513), .A2(new_n688), .A3(new_n689), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n697), .A3(new_n683), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n662), .B1(new_n693), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n687), .B1(new_n699), .B2(new_n517), .ZN(G1328gat));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n518), .A3(new_n412), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT46), .Z(new_n702));
  AOI21_X1  g501(.A(new_n494), .B1(new_n693), .B2(new_n698), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n703), .B2(new_n518), .ZN(G1329gat));
  AOI21_X1  g503(.A(new_n672), .B1(new_n693), .B2(new_n698), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT100), .B1(new_n705), .B2(new_n514), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n685), .A2(new_n514), .A3(new_n505), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n697), .B1(new_n696), .B2(new_n683), .ZN(new_n708));
  AOI211_X1 g507(.A(KEYINPUT99), .B(new_n684), .C1(new_n694), .C2(new_n695), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n492), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT100), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(G43gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n706), .A2(new_n707), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G43gat), .B1(new_n692), .B2(new_n672), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(KEYINPUT47), .A3(new_n707), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(G1330gat));
  OAI21_X1  g517(.A(new_n526), .B1(new_n692), .B2(new_n675), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n685), .A2(new_n524), .A3(new_n501), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(KEYINPUT48), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n720), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n501), .B1(new_n708), .B2(new_n709), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(new_n526), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT101), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n724), .A2(new_n725), .A3(KEYINPUT48), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n675), .B1(new_n693), .B2(new_n698), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n720), .B1(new_n727), .B2(new_n524), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT101), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n721), .B1(new_n726), .B2(new_n730), .ZN(G1331gat));
  INV_X1    g530(.A(new_n638), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n679), .A2(new_n732), .A3(new_n689), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n570), .A2(new_n657), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n661), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g537(.A(new_n494), .B(new_n735), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n739), .B(new_n742), .ZN(G1333gat));
  NAND3_X1  g542(.A1(new_n736), .A2(new_n602), .A3(new_n505), .ZN(new_n744));
  OAI21_X1  g543(.A(G71gat), .B1(new_n735), .B2(new_n672), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g546(.A1(new_n735), .A2(new_n675), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT104), .B(G78gat), .Z(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1335gat));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n732), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT105), .Z(new_n752));
  NAND2_X1  g551(.A1(new_n696), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT106), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(G85gat), .A3(new_n661), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n513), .A2(new_n681), .A3(new_n732), .A4(new_n689), .ZN(new_n757));
  OR3_X1    g556(.A1(new_n757), .A2(KEYINPUT107), .A3(KEYINPUT51), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT107), .B(KEYINPUT51), .Z(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n758), .A2(new_n661), .A3(new_n682), .A4(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n756), .B1(new_n282), .B2(new_n761), .ZN(G1336gat));
  NAND3_X1  g561(.A1(new_n412), .A2(new_n575), .A3(new_n682), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT108), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n758), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(G92gat), .B1(new_n753), .B2(new_n494), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n754), .A2(new_n412), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n757), .A2(KEYINPUT109), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n769), .A2(G92gat), .B1(new_n764), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n768), .B1(new_n775), .B2(new_n767), .ZN(G1337gat));
  AND4_X1   g575(.A1(new_n505), .A2(new_n758), .A3(new_n682), .A4(new_n760), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n754), .A2(new_n492), .ZN(new_n778));
  MUX2_X1   g577(.A(new_n777), .B(new_n778), .S(G99gat), .Z(G1338gat));
  NOR2_X1   g578(.A1(new_n675), .A2(G106gat), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n772), .A2(new_n682), .A3(new_n773), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT111), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT110), .B(G106gat), .Z(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n754), .B2(new_n501), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT53), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n758), .A2(new_n682), .A3(new_n760), .A4(new_n780), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n753), .A2(new_n675), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n786), .B(new_n787), .C1(new_n783), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(G1339gat));
  NAND3_X1  g589(.A1(new_n649), .A2(new_n641), .A3(new_n650), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT54), .ZN(new_n792));
  AND2_X1   g591(.A1(KEYINPUT112), .A2(KEYINPUT54), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n651), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n649), .A2(new_n650), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n640), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n796), .A2(new_n797), .A3(KEYINPUT54), .A4(new_n791), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n798), .A3(new_n656), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  INV_X1    g599(.A(new_n656), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n653), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n794), .A2(new_n798), .A3(new_n800), .A4(new_n656), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n570), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n554), .A2(new_n556), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT113), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n548), .B1(new_n547), .B2(new_n549), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n565), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(new_n569), .A3(new_n682), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(KEYINPUT114), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n567), .A2(new_n569), .B1(new_n803), .B2(new_n804), .ZN(new_n814));
  INV_X1    g613(.A(new_n811), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n812), .A2(new_n816), .A3(new_n680), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n689), .A2(new_n569), .A3(new_n805), .A4(new_n810), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n638), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n658), .A2(new_n570), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n821), .A2(new_n507), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n661), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n412), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n681), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n570), .A2(new_n218), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(KEYINPUT115), .Z(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n825), .B2(new_n828), .ZN(G1340gat));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n682), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g630(.A1(new_n824), .A2(new_n638), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g632(.A1(new_n823), .A2(G134gat), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n689), .A2(new_n494), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT116), .Z(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n838));
  OAI21_X1  g637(.A(G134gat), .B1(new_n825), .B2(new_n680), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G1343gat));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n821), .A2(new_n501), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n662), .A2(new_n492), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n494), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n570), .A2(new_n206), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT119), .Z(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n842), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  XOR2_X1   g651(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n843), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n680), .B1(new_n814), .B2(new_n815), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n818), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n732), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI22_X1  g658(.A1(new_n859), .A2(KEYINPUT118), .B1(new_n570), .B2(new_n658), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT57), .B(new_n501), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n846), .B1(new_n855), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n570), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n852), .B1(new_n864), .B2(G141gat), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n865), .B(new_n866), .ZN(G1344gat));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n659), .B2(new_n681), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n680), .A2(KEYINPUT97), .A3(new_n638), .A4(new_n657), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT97), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n658), .A2(new_n872), .ZN(new_n873));
  AND4_X1   g672(.A1(new_n869), .A2(new_n871), .A3(new_n681), .A4(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n858), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT122), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n877), .B(new_n858), .C1(new_n870), .C2(new_n874), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n501), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n501), .B(new_n853), .C1(new_n819), .C2(new_n820), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n682), .B(new_n847), .C1(new_n881), .C2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n868), .B1(new_n884), .B2(G148gat), .ZN(new_n885));
  AOI211_X1 g684(.A(KEYINPUT59), .B(new_n204), .C1(new_n863), .C2(new_n682), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n682), .A2(new_n204), .ZN(new_n887));
  OAI22_X1  g686(.A1(new_n885), .A2(new_n886), .B1(new_n848), .B2(new_n887), .ZN(G1345gat));
  NOR2_X1   g687(.A1(new_n732), .A2(new_n214), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n844), .A2(new_n638), .A3(new_n847), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n863), .A2(new_n889), .B1(new_n890), .B2(new_n214), .ZN(G1346gat));
  NAND4_X1  g690(.A1(new_n844), .A2(new_n215), .A3(new_n836), .A4(new_n845), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n863), .A2(new_n689), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n215), .ZN(G1347gat));
  NAND4_X1  g693(.A1(new_n821), .A2(new_n662), .A3(new_n412), .A4(new_n507), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n681), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(new_n328), .ZN(G1348gat));
  NOR2_X1   g696(.A1(new_n895), .A2(new_n657), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(new_n329), .ZN(G1349gat));
  NOR2_X1   g698(.A1(new_n895), .A2(new_n732), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n354), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n901), .B1(new_n338), .B2(new_n900), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT60), .ZN(G1350gat));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G190gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n895), .A2(new_n680), .ZN(new_n906));
  MUX2_X1   g705(.A(new_n904), .B(new_n905), .S(new_n906), .Z(G1351gat));
  AOI21_X1  g706(.A(new_n883), .B1(new_n879), .B2(new_n880), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n661), .A2(new_n492), .A3(new_n494), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n570), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT123), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n914), .A3(new_n570), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(G197gat), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n821), .A2(new_n501), .A3(new_n909), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(new_n309), .A3(new_n570), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(G1352gat));
  NOR3_X1   g719(.A1(new_n917), .A2(G204gat), .A3(new_n657), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n923), .A2(KEYINPUT62), .A3(new_n924), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n908), .A2(new_n657), .A3(new_n910), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n927), .B(new_n928), .C1(new_n307), .C2(new_n929), .ZN(G1353gat));
  NAND3_X1  g729(.A1(new_n918), .A2(new_n300), .A3(new_n638), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n300), .B1(new_n911), .B2(new_n638), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n932), .A2(KEYINPUT63), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(KEYINPUT63), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1354gat));
  OAI211_X1 g734(.A(KEYINPUT126), .B(new_n909), .C1(new_n881), .C2(new_n883), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n937), .B1(new_n908), .B2(new_n910), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n302), .A2(new_n303), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n936), .A2(new_n938), .A3(new_n939), .A4(new_n689), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n318), .B1(new_n917), .B2(new_n680), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT127), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n940), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1355gat));
endmodule


