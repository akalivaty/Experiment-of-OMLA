//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT4), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G107), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT3), .A3(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  OR3_X1    g014(.A1(new_n197), .A2(KEYINPUT79), .A3(G104), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT79), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n193), .B(G101), .C1(new_n200), .C2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n208), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  INV_X1    g032(.A(new_n204), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(new_n199), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n199), .A2(new_n218), .A3(new_n201), .A4(new_n203), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT4), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n205), .B(new_n217), .C1(new_n220), .C2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n207), .A2(new_n224), .A3(G128), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n210), .B(G146), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n212), .A3(G143), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n197), .A2(G104), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n202), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G101), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n232), .A3(new_n221), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT10), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n221), .A2(new_n232), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n227), .A2(new_n228), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n227), .A2(KEYINPUT67), .A3(new_n228), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(new_n225), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(KEYINPUT10), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n223), .A2(new_n235), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G131), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT66), .ZN(new_n245));
  INV_X1    g059(.A(G134), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT11), .B1(new_n246), .B2(G137), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n248));
  INV_X1    g062(.A(G137), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G134), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n252), .B1(new_n249), .B2(G134), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n246), .A2(KEYINPUT65), .A3(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n245), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n253), .A2(new_n254), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n247), .A2(new_n250), .ZN(new_n258));
  INV_X1    g072(.A(new_n245), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n243), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n261), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n223), .A2(new_n235), .A3(new_n242), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G110), .B(G140), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G227), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n266), .B(new_n268), .Z(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT12), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n233), .B1(new_n236), .B2(new_n241), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(new_n274), .B2(new_n261), .ZN(new_n275));
  NOR2_X1   g089(.A1(KEYINPUT80), .A2(KEYINPUT12), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n269), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n274), .A2(new_n261), .A3(new_n271), .A4(new_n272), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n278), .A2(new_n264), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n270), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n192), .B1(new_n282), .B2(new_n190), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n278), .A2(new_n264), .A3(new_n280), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n269), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n262), .A2(new_n264), .A3(new_n279), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(G469), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n189), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G119), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G116), .ZN(new_n291));
  INV_X1    g105(.A(G116), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G119), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT2), .B(G113), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OR2_X1    g110(.A1(new_n291), .A2(KEYINPUT5), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n291), .A2(new_n293), .A3(KEYINPUT5), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .A4(G113), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(G113), .A3(new_n299), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT81), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n236), .A2(new_n296), .A3(new_n300), .A4(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n294), .A2(new_n295), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n296), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT68), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n296), .A2(KEYINPUT68), .A3(new_n304), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(new_n205), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n220), .A2(new_n222), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G110), .B(G122), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n303), .B(new_n312), .C1(new_n309), .C2(new_n310), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(KEYINPUT6), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n241), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n217), .A2(G125), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n267), .A2(G224), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT82), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT6), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n311), .A2(new_n325), .A3(new_n313), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n316), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(KEYINPUT7), .B(new_n322), .C1(new_n318), .C2(new_n320), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n301), .A2(new_n296), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n236), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n312), .B(KEYINPUT8), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n302), .A2(new_n296), .A3(new_n300), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n330), .B(new_n331), .C1(new_n332), .C2(new_n236), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n322), .A2(KEYINPUT7), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n319), .B(new_n334), .C1(new_n317), .C2(G125), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n328), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(G902), .B1(new_n336), .B2(new_n315), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(G210), .B1(G237), .B2(G902), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n327), .A2(new_n337), .A3(new_n339), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G214), .B1(G237), .B2(G902), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT15), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G478), .ZN(new_n347));
  XNOR2_X1  g161(.A(G128), .B(G143), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(new_n246), .ZN(new_n349));
  INV_X1    g163(.A(G122), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G116), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n292), .A2(G122), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(new_n197), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n352), .A2(KEYINPUT14), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n351), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(KEYINPUT14), .B2(new_n352), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n349), .B(new_n353), .C1(new_n356), .C2(new_n197), .ZN(new_n357));
  INV_X1    g171(.A(G217), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n187), .A2(new_n358), .A3(G953), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n197), .B1(new_n351), .B2(new_n352), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT87), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n353), .ZN(new_n363));
  INV_X1    g177(.A(new_n353), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT87), .B1(new_n364), .B2(new_n360), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  XOR2_X1   g180(.A(KEYINPUT88), .B(KEYINPUT13), .Z(new_n367));
  AOI21_X1  g181(.A(new_n246), .B1(new_n367), .B2(new_n348), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(G128), .A3(new_n210), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n368), .A2(new_n370), .B1(new_n246), .B2(new_n348), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT89), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n366), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n372), .B1(new_n366), .B2(new_n371), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n357), .B(new_n359), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT90), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n366), .A2(new_n371), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT89), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n366), .A2(new_n371), .A3(new_n372), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n357), .A4(new_n359), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n357), .B1(new_n373), .B2(new_n374), .ZN(new_n383));
  INV_X1    g197(.A(new_n359), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n376), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n347), .B1(new_n386), .B2(new_n191), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n191), .A3(new_n347), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G140), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G125), .ZN(new_n392));
  INV_X1    g206(.A(G125), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT76), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G125), .B(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT76), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n399), .A3(new_n212), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT75), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n393), .A2(KEYINPUT75), .A3(G140), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(G146), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT18), .A2(G131), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G237), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n267), .A3(G214), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(KEYINPUT83), .B2(new_n210), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT83), .B(G143), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n410), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n405), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(G237), .A2(G953), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G143), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n210), .A2(KEYINPUT83), .ZN(new_n417));
  OAI211_X1 g231(.A(G214), .B(new_n414), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n410), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n419), .B1(new_n418), .B2(new_n410), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n407), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT85), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n412), .A2(KEYINPUT84), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n420), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n407), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n413), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G113), .B(G122), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n430), .B(new_n195), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n412), .A2(G131), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT17), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n418), .A2(new_n244), .A3(new_n410), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(KEYINPUT16), .B(new_n403), .C1(new_n395), .C2(KEYINPUT75), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT16), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n392), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(new_n212), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n439), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G146), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n412), .A2(KEYINPUT17), .A3(G131), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n436), .A2(new_n440), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n429), .A2(new_n432), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n413), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n427), .B1(new_n426), .B2(new_n407), .ZN(new_n448));
  AOI211_X1 g262(.A(KEYINPUT85), .B(new_n406), .C1(new_n425), .C2(new_n420), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n431), .B1(new_n450), .B2(new_n444), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n191), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G475), .ZN(new_n453));
  INV_X1    g267(.A(G234), .ZN(new_n454));
  OAI211_X1 g268(.A(G952), .B(new_n267), .C1(new_n454), .C2(new_n408), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT91), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(G898), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT92), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n191), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n456), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n433), .A2(new_n435), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n442), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT19), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n397), .A2(new_n399), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n402), .A2(KEYINPUT19), .A3(new_n403), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n465), .B1(new_n469), .B2(G146), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT86), .A4(new_n212), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n432), .B1(new_n429), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n450), .A2(new_n431), .A3(new_n444), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(G475), .A2(G902), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n462), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n476), .ZN(new_n478));
  AOI211_X1 g292(.A(KEYINPUT20), .B(new_n478), .C1(new_n473), .C2(new_n474), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n453), .B(new_n461), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  NOR4_X1   g294(.A1(new_n289), .A2(new_n345), .A3(new_n390), .A4(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n251), .A2(new_n255), .A3(new_n245), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n259), .B1(new_n257), .B2(new_n258), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n217), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n307), .A2(new_n308), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n246), .A2(G137), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n249), .A2(G134), .ZN(new_n488));
  OAI21_X1  g302(.A(G131), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n257), .A2(new_n244), .A3(new_n258), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n241), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT69), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n261), .A2(new_n492), .A3(new_n217), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n485), .A2(new_n486), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT64), .ZN(new_n496));
  INV_X1    g310(.A(new_n206), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n214), .B2(new_n215), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n207), .A2(new_n208), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n209), .A2(new_n216), .A3(KEYINPUT64), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n500), .B(new_n501), .C1(new_n482), .C2(new_n483), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n486), .B1(new_n502), .B2(new_n491), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT28), .B1(new_n495), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n486), .A2(new_n491), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT28), .B1(new_n505), .B2(new_n484), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n509));
  NAND2_X1  g323(.A1(new_n414), .A2(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G101), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n513), .B(KEYINPUT72), .Z(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT31), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT71), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n256), .A2(new_n260), .B1(new_n216), .B2(new_n209), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n491), .B1(new_n519), .B2(new_n492), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n261), .A2(new_n492), .A3(new_n217), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT30), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n502), .A2(new_n523), .A3(new_n491), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n486), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n513), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n494), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n518), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n494), .A2(new_n526), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n502), .A2(new_n523), .A3(new_n491), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n485), .A2(new_n491), .A3(new_n493), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(KEYINPUT30), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT71), .B(new_n529), .C1(new_n532), .C2(new_n486), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n517), .B1(new_n528), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n486), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n490), .A2(new_n489), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n484), .A2(KEYINPUT69), .B1(new_n536), .B2(new_n241), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n523), .B1(new_n537), .B2(new_n493), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n535), .B1(new_n538), .B2(new_n530), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT31), .B1(new_n539), .B2(new_n529), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n516), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(G472), .A2(G902), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n516), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT71), .B1(new_n539), .B2(new_n529), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n525), .A2(new_n518), .A3(new_n527), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT31), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n540), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n542), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n544), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT73), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT29), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n525), .A2(new_n495), .ZN(new_n557));
  OAI221_X1 g371(.A(new_n556), .B1(new_n557), .B2(new_n526), .C1(new_n508), .C2(new_n515), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n531), .A2(new_n535), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n494), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n506), .B1(new_n560), .B2(KEYINPUT28), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n513), .A2(new_n556), .ZN(new_n562));
  AOI21_X1  g376(.A(G902), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G472), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT73), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n541), .A2(new_n566), .A3(new_n553), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n545), .A2(new_n555), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT77), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT22), .B(G137), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G119), .B(G128), .ZN(new_n574));
  INV_X1    g388(.A(G110), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n575), .A2(KEYINPUT24), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(KEYINPUT24), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT74), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT24), .B(G110), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT74), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n574), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT23), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n290), .B2(G128), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n226), .A2(KEYINPUT23), .A3(G119), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n584), .B(new_n585), .C1(G119), .C2(new_n226), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(G110), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n400), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n212), .B1(new_n437), .B2(new_n439), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n578), .A2(new_n581), .A3(new_n574), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(G110), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n442), .B2(new_n440), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n573), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n440), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n591), .B(new_n592), .C1(new_n597), .C2(new_n589), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n442), .B(new_n400), .C1(new_n587), .C2(new_n582), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n599), .A3(new_n572), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(G217), .B1(new_n454), .B2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n191), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n596), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n595), .A2(new_n600), .A3(new_n191), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT25), .B1(new_n605), .B2(KEYINPUT78), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(new_n602), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n481), .A2(new_n568), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  NAND2_X1  g425(.A1(new_n541), .A2(new_n191), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(G472), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n613), .A2(new_n543), .A3(new_n609), .A4(new_n288), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n470), .A2(new_n471), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n442), .A3(new_n463), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n431), .B1(new_n616), .B2(new_n450), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n476), .B1(new_n446), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT20), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n475), .A2(new_n462), .A3(new_n476), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n386), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n385), .A2(KEYINPUT33), .A3(new_n375), .ZN(new_n624));
  INV_X1    g438(.A(G478), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(G902), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n386), .A2(new_n191), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n625), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n621), .A2(new_n453), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT93), .ZN(new_n631));
  INV_X1    g445(.A(new_n344), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n341), .B2(new_n342), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n630), .A2(new_n631), .A3(new_n633), .A4(new_n461), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n627), .A2(new_n629), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n453), .B1(new_n477), .B2(new_n479), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n327), .A2(new_n337), .A3(new_n339), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n339), .B1(new_n327), .B2(new_n337), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n344), .B(new_n461), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT93), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n614), .B1(new_n634), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT34), .B(G104), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(new_n636), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n390), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n461), .B(KEYINPUT94), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n633), .A2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n614), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT35), .B(G107), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NOR2_X1   g465(.A1(new_n289), .A2(new_n345), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n598), .A2(new_n599), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT95), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n603), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n657), .A2(new_n658), .B1(new_n608), .B2(new_n607), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n659), .A2(new_n480), .A3(new_n390), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n652), .A2(new_n543), .A3(new_n613), .A4(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  NAND2_X1  g477(.A1(new_n607), .A2(new_n608), .ZN(new_n664));
  INV_X1    g478(.A(new_n657), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n664), .B1(new_n665), .B2(new_n603), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n288), .A3(new_n633), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n541), .A2(new_n566), .A3(new_n553), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n566), .B1(new_n541), .B2(new_n553), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n543), .A2(new_n544), .B1(new_n564), .B2(G472), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n456), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(new_n459), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n646), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  NAND2_X1  g492(.A1(new_n528), .A2(new_n533), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n514), .B1(new_n494), .B2(new_n559), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n191), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G472), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n545), .A2(new_n555), .A3(new_n567), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT96), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT96), .ZN(new_n685));
  AOI22_X1  g499(.A1(new_n543), .A2(new_n544), .B1(G472), .B2(new_n681), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n670), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n390), .A2(new_n636), .A3(new_n344), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n659), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT97), .Z(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT98), .B(KEYINPUT39), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n675), .B(new_n693), .Z(new_n694));
  NOR2_X1   g508(.A1(new_n289), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT40), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n343), .B(KEYINPUT38), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NOR4_X1   g512(.A1(new_n689), .A2(new_n692), .A3(new_n696), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n210), .ZN(G45));
  OR2_X1    g514(.A1(new_n637), .A2(new_n675), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n667), .B(new_n701), .C1(new_n670), .C2(new_n671), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n212), .ZN(G48));
  NAND2_X1  g517(.A1(KEYINPUT99), .A2(G469), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n279), .B1(new_n262), .B2(new_n264), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n264), .A2(new_n280), .ZN(new_n707));
  AOI211_X1 g521(.A(new_n273), .B(new_n276), .C1(new_n274), .C2(new_n261), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n706), .B1(new_n709), .B2(new_n279), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n705), .B1(new_n710), .B2(G902), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n282), .A2(new_n704), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n711), .A2(new_n712), .A3(new_n188), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n609), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n634), .B2(new_n641), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n568), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NOR3_X1   g532(.A1(new_n714), .A2(new_n648), .A3(new_n646), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT100), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n568), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n720), .B1(new_n568), .B2(new_n719), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n292), .ZN(G18));
  AND3_X1   g538(.A1(new_n660), .A2(new_n633), .A3(new_n713), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n725), .A2(new_n568), .A3(KEYINPUT101), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT101), .B1(new_n725), .B2(new_n568), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT102), .B(G119), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G21));
  INV_X1    g544(.A(new_n713), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n343), .A2(new_n390), .A3(new_n636), .A4(new_n344), .ZN(new_n732));
  INV_X1    g546(.A(new_n647), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(G472), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n541), .B2(new_n191), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n549), .A2(new_n550), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n561), .A2(new_n514), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n552), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n609), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n736), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NAND2_X1  g557(.A1(new_n713), .A2(new_n633), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n701), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT103), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n738), .B1(new_n534), .B2(new_n540), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n612), .A2(G472), .B1(new_n747), .B2(new_n542), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n746), .B1(new_n748), .B2(new_n666), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n736), .A2(new_n739), .A3(KEYINPUT103), .A4(new_n659), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n745), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  OAI21_X1  g566(.A(new_n671), .B1(new_n551), .B2(new_n554), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n638), .A2(new_n639), .A3(new_n189), .A4(new_n632), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n284), .A2(KEYINPUT104), .A3(new_n269), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT104), .B1(new_n284), .B2(new_n269), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n286), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n283), .B1(new_n758), .B2(new_n190), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n701), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n753), .A2(new_n761), .A3(new_n609), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT42), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n740), .B1(new_n670), .B2(new_n671), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n765), .A3(new_n761), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  NOR3_X1   g582(.A1(new_n760), .A2(new_n646), .A3(new_n675), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n568), .A3(new_n609), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  OAI211_X1 g585(.A(KEYINPUT45), .B(new_n286), .C1(new_n756), .C2(new_n757), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n285), .B2(new_n286), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n190), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n192), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n778), .A2(KEYINPUT46), .B1(new_n190), .B2(new_n282), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT105), .B1(new_n778), .B2(KEYINPUT46), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n778), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n188), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n784));
  OR3_X1    g598(.A1(new_n783), .A2(new_n784), .A3(new_n694), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n784), .B1(new_n783), .B2(new_n694), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT43), .B1(new_n645), .B2(KEYINPUT107), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n636), .B1(new_n629), .B2(new_n627), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n787), .B(new_n788), .Z(new_n789));
  NAND2_X1  g603(.A1(new_n613), .A2(new_n543), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n790), .A3(new_n666), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n343), .A2(new_n632), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n791), .B2(new_n792), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n785), .A2(new_n786), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT108), .B(G137), .Z(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(G39));
  INV_X1    g613(.A(new_n568), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n701), .A2(new_n795), .A3(new_n609), .ZN(new_n801));
  INV_X1    g615(.A(new_n783), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT47), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(KEYINPUT47), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n800), .B(new_n801), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  AND2_X1   g620(.A1(new_n698), .A2(new_n788), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n711), .A2(new_n712), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT49), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n609), .A2(new_n188), .A3(new_n344), .ZN(new_n810));
  XOR2_X1   g624(.A(new_n810), .B(KEYINPUT109), .Z(new_n811));
  NAND4_X1  g625(.A1(new_n689), .A2(new_n807), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n789), .A2(new_n673), .A3(new_n741), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n744), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n267), .A2(KEYINPUT116), .A3(G952), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT116), .B1(new_n267), .B2(G952), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n754), .A2(new_n673), .A3(new_n808), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n789), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n753), .A2(new_n609), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(KEYINPUT117), .A3(KEYINPUT48), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n820), .ZN(new_n823));
  XOR2_X1   g637(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n824));
  AOI21_X1  g638(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n689), .A2(new_n609), .A3(new_n818), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n697), .A2(new_n344), .A3(new_n731), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT115), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n813), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT50), .ZN(new_n830));
  OR3_X1    g644(.A1(new_n826), .A2(new_n636), .A3(new_n635), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n747), .A2(new_n542), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n613), .A2(new_n666), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT103), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n748), .A2(new_n746), .A3(new_n666), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n819), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n830), .A2(KEYINPUT51), .A3(new_n831), .A4(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n813), .A2(new_n795), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n803), .A2(new_n804), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n808), .A2(new_n189), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI221_X1 g657(.A(new_n825), .B1(new_n637), .B2(new_n826), .C1(new_n838), .C2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n830), .A2(new_n831), .A3(new_n837), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n803), .B2(new_n804), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n842), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(KEYINPUT114), .B2(new_n841), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n845), .B1(new_n849), .B2(new_n840), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  XOR2_X1   g666(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n853));
  NAND2_X1  g667(.A1(new_n751), .A2(new_n677), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n666), .A2(new_n189), .A3(new_n675), .ZN(new_n855));
  INV_X1    g669(.A(new_n732), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n856), .A3(new_n759), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n684), .B2(new_n687), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n854), .A2(new_n858), .A3(new_n859), .A4(new_n702), .ZN(new_n860));
  INV_X1    g674(.A(new_n857), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n702), .B1(new_n688), .B2(new_n861), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n836), .A2(new_n745), .B1(new_n676), .B2(new_n672), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT52), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n761), .B1(new_n749), .B2(new_n750), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n795), .A2(new_n659), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n390), .A2(new_n636), .A3(new_n675), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n568), .A2(new_n288), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n770), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT110), .ZN(new_n871));
  INV_X1    g685(.A(new_n389), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n387), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n873), .B2(new_n636), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n390), .A2(KEYINPUT110), .A3(new_n453), .A4(new_n621), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n637), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n633), .A3(new_n647), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n610), .B(new_n661), .C1(new_n614), .C2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n715), .A2(new_n568), .B1(new_n734), .B2(new_n741), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n721), .B2(new_n722), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n728), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n882), .A3(new_n767), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n853), .B1(new_n865), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n683), .A2(KEYINPUT96), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n685), .B1(new_n670), .B2(new_n686), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n861), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n702), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n859), .B1(new_n889), .B2(new_n854), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n862), .A2(KEYINPUT52), .A3(new_n863), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n763), .A2(KEYINPUT53), .A3(new_n766), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT113), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n882), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT112), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n870), .B2(new_n878), .ZN(new_n897));
  INV_X1    g711(.A(new_n610), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n661), .B1(new_n877), .B2(new_n614), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n770), .A2(new_n869), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT112), .A4(new_n866), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT113), .B1(new_n881), .B2(new_n728), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n892), .A2(new_n895), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n884), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n865), .A2(new_n883), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT53), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n853), .B2(new_n908), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n911), .B2(KEYINPUT54), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n852), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT118), .ZN(new_n914));
  OR2_X1    g728(.A1(G952), .A2(G953), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n913), .A2(KEYINPUT118), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n812), .B1(new_n916), .B2(new_n917), .ZN(G75));
  NOR2_X1   g732(.A1(new_n267), .A2(G952), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n884), .A2(new_n905), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n191), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT56), .B1(new_n922), .B2(G210), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n316), .A2(new_n326), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n324), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT55), .Z(new_n926));
  OAI21_X1  g740(.A(new_n920), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n921), .B2(new_n191), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n906), .A2(KEYINPUT119), .A3(G902), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n340), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n927), .B1(new_n931), .B2(new_n933), .ZN(G51));
  INV_X1    g748(.A(new_n775), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n929), .A2(new_n935), .A3(new_n930), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n192), .B(KEYINPUT57), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT121), .B1(new_n906), .B2(KEYINPUT54), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT54), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n939), .B(new_n940), .C1(new_n884), .C2(new_n905), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT120), .B1(new_n906), .B2(KEYINPUT54), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n884), .A2(new_n905), .A3(new_n944), .A4(new_n940), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n937), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n710), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n936), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT122), .B1(new_n949), .B2(new_n919), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n943), .B(new_n945), .C1(new_n938), .C2(new_n941), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n710), .B1(new_n952), .B2(new_n937), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n951), .B(new_n920), .C1(new_n953), .C2(new_n936), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n950), .A2(new_n954), .ZN(G54));
  NAND4_X1  g769(.A1(new_n929), .A2(KEYINPUT58), .A3(G475), .A4(new_n930), .ZN(new_n956));
  INV_X1    g770(.A(new_n475), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n956), .A2(KEYINPUT123), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n920), .B1(new_n956), .B2(new_n957), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT123), .B1(new_n956), .B2(new_n957), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(G60));
  AND2_X1   g775(.A1(new_n623), .A2(new_n624), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT59), .Z(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n952), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n912), .A2(new_n965), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n919), .B(new_n967), .C1(new_n963), .C2(new_n968), .ZN(G63));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT60), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n921), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n596), .A2(new_n601), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n920), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n657), .B2(new_n972), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g790(.A(new_n267), .B1(new_n458), .B2(G224), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n882), .A2(new_n900), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT124), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n977), .B1(new_n980), .B2(new_n267), .ZN(new_n981));
  INV_X1    g795(.A(G898), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n924), .B1(new_n982), .B2(G953), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n981), .B(new_n983), .ZN(G69));
  XOR2_X1   g798(.A(new_n532), .B(new_n469), .Z(new_n985));
  NAND4_X1  g799(.A1(new_n764), .A2(new_n695), .A3(new_n794), .A4(new_n876), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n805), .A2(new_n797), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n863), .A2(new_n888), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n699), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n985), .B1(new_n992), .B2(G953), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n993), .A2(KEYINPUT125), .ZN(new_n994));
  INV_X1    g808(.A(new_n988), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n805), .A2(new_n767), .A3(new_n770), .A4(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n785), .A2(new_n856), .A3(new_n820), .A4(new_n786), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n797), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n267), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n267), .A2(G900), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT126), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n985), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n993), .B2(KEYINPUT125), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n994), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(G72));
  OR3_X1    g820(.A1(new_n980), .A2(new_n996), .A3(new_n998), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G472), .A2(G902), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1010), .A2(new_n513), .A3(new_n557), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n557), .A2(new_n526), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n911), .B(new_n1009), .C1(new_n679), .C2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1011), .A2(new_n920), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n992), .A2(new_n979), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n1009), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT127), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n557), .A2(new_n513), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1017), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n1014), .A2(new_n1019), .A3(new_n1020), .ZN(G57));
endmodule


