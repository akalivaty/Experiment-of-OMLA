//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  OAI22_X1  g000(.A1(KEYINPUT68), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(KEYINPUT68), .A2(KEYINPUT26), .ZN(new_n203));
  AOI22_X1  g002(.A1(new_n202), .A2(new_n203), .B1(G169gat), .B2(G176gat), .ZN(new_n204));
  OAI211_X1 g003(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n205));
  AOI22_X1  g004(.A1(new_n204), .A2(new_n205), .B1(G183gat), .B2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT27), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT27), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT28), .A4(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n211), .A2(KEYINPUT28), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n215), .A2(KEYINPUT67), .A3(new_n208), .A4(new_n210), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n209), .A2(KEYINPUT27), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n207), .A2(G183gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT66), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221));
  AOI21_X1  g020(.A(G190gat), .B1(new_n208), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT28), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n206), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n211), .ZN(new_n225));
  NAND3_X1  g024(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n229));
  OR3_X1    g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G169gat), .ZN(new_n231));
  INV_X1    g030(.A(G176gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT23), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n233), .B(new_n235), .C1(new_n231), .C2(new_n232), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(KEYINPUT25), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n228), .B1(new_n227), .B2(new_n229), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n230), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n229), .A2(KEYINPUT65), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n229), .A2(KEYINPUT65), .ZN(new_n241));
  NOR3_X1   g040(.A1(new_n240), .A2(new_n241), .A3(new_n227), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT25), .B1(new_n242), .B2(new_n236), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n224), .A2(new_n239), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT70), .ZN(new_n245));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G134gat), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT69), .B1(new_n249), .B2(G127gat), .ZN(new_n250));
  INV_X1    g049(.A(G120gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G113gat), .ZN(new_n252));
  INV_X1    g051(.A(G113gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G120gat), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI22_X1  g054(.A1(new_n248), .A2(new_n250), .B1(KEYINPUT1), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT1), .B1(new_n252), .B2(new_n254), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n246), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n224), .A2(new_n239), .A3(new_n261), .A4(new_n243), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n224), .A2(new_n243), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n264), .A2(new_n261), .A3(new_n259), .A4(new_n239), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G227gat), .ZN(new_n267));
  INV_X1    g066(.A(G233gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n271), .A2(KEYINPUT34), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(KEYINPUT34), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT32), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n263), .A2(new_n269), .A3(new_n265), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n263), .A2(KEYINPUT71), .A3(new_n269), .A4(new_n265), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT33), .B1(new_n279), .B2(new_n280), .ZN(new_n282));
  XNOR2_X1  g081(.A(G15gat), .B(G43gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G71gat), .B(G99gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n281), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n285), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n287), .A2(KEYINPUT72), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(KEYINPUT72), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n288), .A2(KEYINPUT33), .A3(new_n289), .ZN(new_n290));
  AOI211_X1 g089(.A(new_n276), .B(new_n290), .C1(new_n279), .C2(new_n280), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n275), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT36), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n279), .A2(new_n280), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n285), .B1(new_n294), .B2(KEYINPUT32), .ZN(new_n295));
  INV_X1    g094(.A(new_n282), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n291), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(new_n274), .A3(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n292), .A2(new_n293), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n291), .B1(new_n295), .B2(new_n296), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT73), .B1(new_n301), .B2(new_n274), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n303), .B(new_n275), .C1(new_n286), .C2(new_n291), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n300), .B1(KEYINPUT36), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G1gat), .B(G29gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT0), .ZN(new_n308));
  XNOR2_X1  g107(.A(G57gat), .B(G85gat), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n308), .B(new_n309), .Z(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G141gat), .B(G148gat), .ZN(new_n312));
  INV_X1    g111(.A(G162gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G155gat), .ZN(new_n314));
  INV_X1    g113(.A(G155gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G162gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n312), .B1(KEYINPUT75), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT76), .B(G162gat), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT2), .B1(new_n319), .B2(new_n315), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n314), .A2(new_n316), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n317), .B1(new_n312), .B2(KEYINPUT2), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n323), .A2(new_n256), .A3(new_n324), .A4(new_n258), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n324), .A2(new_n323), .B1(new_n256), .B2(new_n258), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT77), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT5), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n323), .A2(new_n324), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n260), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(KEYINPUT3), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n330), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n326), .A2(KEYINPUT78), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n325), .B2(KEYINPUT4), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n325), .A2(KEYINPUT4), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n340), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n332), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n326), .A2(new_n339), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT5), .B1(new_n346), .B2(new_n343), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(KEYINPUT6), .B(new_n311), .C1(new_n345), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT79), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n338), .A2(new_n344), .ZN(new_n351));
  INV_X1    g150(.A(new_n332), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n347), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n310), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT6), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n355), .A2(KEYINPUT6), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n310), .A3(new_n354), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n350), .A2(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n244), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n244), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n364), .B2(new_n361), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT74), .B(G197gat), .ZN(new_n366));
  INV_X1    g165(.A(G204gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G211gat), .B(G218gat), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT22), .ZN(new_n370));
  INV_X1    g169(.A(G211gat), .ZN(new_n371));
  INV_X1    g170(.A(G218gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n368), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n369), .B1(new_n368), .B2(new_n373), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n365), .A2(new_n376), .ZN(new_n377));
  OAI221_X1 g176(.A(new_n362), .B1(new_n375), .B2(new_n374), .C1(new_n364), .C2(new_n361), .ZN(new_n378));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  AND3_X1   g180(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n378), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n383), .B2(KEYINPUT37), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT37), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n377), .A2(new_n378), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n382), .B1(new_n387), .B2(KEYINPUT38), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT38), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n384), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n360), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392));
  INV_X1    g191(.A(G50gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n368), .A2(new_n373), .ZN(new_n398));
  INV_X1    g197(.A(new_n369), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n368), .A2(new_n369), .A3(new_n373), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT29), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n333), .B1(new_n402), .B2(KEYINPUT3), .ZN(new_n403));
  INV_X1    g202(.A(G22gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n363), .B1(new_n333), .B2(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n376), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n404), .B1(new_n403), .B2(new_n406), .ZN(new_n409));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n403), .B2(KEYINPUT81), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n363), .B1(new_n374), .B2(new_n375), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n334), .B1(new_n413), .B2(new_n335), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n415));
  OAI211_X1 g214(.A(G228gat), .B(G233gat), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n406), .ZN(new_n417));
  OAI21_X1  g216(.A(G22gat), .B1(new_n417), .B2(new_n414), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(new_n407), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n397), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n411), .B1(new_n408), .B2(new_n409), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n416), .A2(new_n418), .A3(new_n407), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n396), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n381), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n383), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(KEYINPUT30), .A3(new_n427), .ZN(new_n428));
  OR3_X1    g227(.A1(new_n383), .A2(KEYINPUT30), .A3(new_n425), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT40), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n336), .A2(new_n337), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n346), .A2(new_n343), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n330), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n310), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n435), .B1(new_n328), .B2(new_n331), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n434), .B2(new_n330), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n431), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n311), .B1(new_n345), .B2(new_n348), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n434), .A2(new_n330), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n438), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n444), .A2(KEYINPUT40), .A3(new_n310), .A4(new_n436), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n441), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n424), .B1(new_n430), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n442), .A2(new_n359), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n356), .B1(new_n355), .B2(KEYINPUT6), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n349), .A2(KEYINPUT79), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n428), .A2(new_n429), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n391), .A2(new_n447), .B1(new_n454), .B2(new_n424), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n424), .B1(new_n301), .B2(new_n274), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n357), .A2(new_n350), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n457), .A2(new_n449), .B1(new_n429), .B2(new_n428), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n302), .A2(new_n456), .A3(new_n304), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT35), .ZN(new_n460));
  INV_X1    g259(.A(new_n424), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n292), .A2(new_n299), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n458), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n306), .A2(new_n455), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n466));
  XNOR2_X1  g265(.A(G15gat), .B(G22gat), .ZN(new_n467));
  INV_X1    g266(.A(G1gat), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n468), .A2(KEYINPUT16), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n467), .A2(new_n468), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT84), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT83), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(G8gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n467), .A2(new_n469), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n468), .B2(new_n467), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT83), .B1(new_n476), .B2(KEYINPUT84), .ZN(new_n477));
  INV_X1    g276(.A(G8gat), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n476), .B2(KEYINPUT83), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n474), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G29gat), .ZN(new_n481));
  INV_X1    g280(.A(G36gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT14), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(G29gat), .B2(G36gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT82), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n483), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n487), .B(new_n489), .C1(new_n481), .C2(new_n482), .ZN(new_n490));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n486), .B1(new_n492), .B2(new_n493), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n491), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT88), .B1(new_n480), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n501));
  XOR2_X1   g300(.A(G15gat), .B(G22gat), .Z(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G1gat), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n503), .B2(new_n475), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n473), .B1(new_n503), .B2(new_n475), .ZN(new_n505));
  OAI22_X1  g304(.A1(KEYINPUT83), .A2(new_n504), .B1(new_n505), .B2(new_n478), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n490), .A2(new_n494), .B1(new_n497), .B2(new_n496), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT88), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .A4(new_n474), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n480), .A2(new_n499), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n500), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G229gat), .A2(G233gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT85), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT13), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n506), .B(new_n474), .C1(new_n507), .C2(KEYINPUT17), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n499), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n510), .B(new_n513), .C1(new_n516), .C2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n480), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT17), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n499), .A2(new_n517), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n525), .A2(KEYINPUT18), .A3(new_n510), .A4(new_n513), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n515), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n515), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G197gat), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT11), .B(G169gat), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT12), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n527), .A2(new_n529), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n527), .B1(new_n529), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n466), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n515), .A2(new_n526), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n539), .B(new_n521), .C1(new_n528), .C2(new_n534), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n527), .A2(new_n529), .A3(new_n535), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT89), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n465), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT21), .ZN(new_n546));
  OR2_X1    g345(.A1(G57gat), .A2(G64gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(G57gat), .A2(G64gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT91), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT92), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n547), .A2(new_n555), .A3(new_n548), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n550), .A2(new_n553), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G71gat), .ZN(new_n558));
  INV_X1    g357(.A(G78gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n561), .A2(KEYINPUT90), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(KEYINPUT90), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n557), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n553), .A2(new_n554), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n560), .A2(new_n561), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n567), .A2(new_n549), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n522), .B1(new_n546), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n571), .B(new_n572), .Z(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n578), .B(new_n579), .Z(new_n580));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n578), .B(new_n579), .ZN(new_n583));
  INV_X1    g382(.A(new_n581), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G183gat), .B(G211gat), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n582), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n582), .B2(new_n585), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n574), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n582), .A2(new_n585), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n586), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n582), .A2(new_n587), .A3(new_n585), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n593), .A3(new_n573), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n597));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(G99gat), .A2(G106gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT97), .B(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(KEYINPUT8), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(G85gat), .A3(G92gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT7), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n604), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n611), .B(KEYINPUT7), .ZN(new_n615));
  INV_X1    g414(.A(new_n604), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n615), .A2(new_n616), .A3(new_n607), .A4(new_n608), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n524), .A2(new_n523), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G190gat), .B(G218gat), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n507), .B2(new_n618), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n623), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n625), .B1(new_n623), .B2(new_n628), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n600), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n633), .A2(new_n599), .A3(new_n629), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n595), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n557), .A2(new_n564), .B1(new_n566), .B2(new_n568), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n637), .A2(KEYINPUT10), .A3(new_n617), .A4(new_n614), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n614), .A2(new_n617), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n641), .A2(KEYINPUT100), .A3(KEYINPUT10), .A4(new_n637), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n637), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n570), .A2(new_n618), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT99), .B(KEYINPUT10), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n644), .B2(new_n645), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(G176gat), .B(G204gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n653), .B(new_n654), .Z(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n655), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n649), .B(KEYINPUT101), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n643), .B2(new_n647), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n659), .B2(new_n651), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n636), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n545), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n452), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(new_n468), .ZN(G1324gat));
  INV_X1    g464(.A(new_n663), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n478), .B1(new_n666), .B2(new_n430), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT16), .B(G8gat), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n663), .A2(new_n453), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT42), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(KEYINPUT42), .B2(new_n669), .ZN(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n663), .B2(new_n306), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n292), .A2(new_n299), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(G15gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n672), .B1(new_n663), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n663), .A2(new_n461), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NAND2_X1  g478(.A1(new_n590), .A2(new_n594), .ZN(new_n680));
  INV_X1    g479(.A(new_n635), .ZN(new_n681));
  INV_X1    g480(.A(new_n661), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n460), .A2(new_n464), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n305), .A2(KEYINPUT36), .ZN(new_n685));
  INV_X1    g484(.A(new_n300), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n455), .A3(new_n686), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n544), .B(new_n683), .C1(new_n684), .C2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n481), .A3(new_n360), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n684), .A2(new_n687), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n691), .B2(new_n681), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  AOI211_X1 g492(.A(new_n693), .B(new_n635), .C1(new_n684), .C2(new_n687), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n682), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n540), .A2(new_n541), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n695), .A2(new_n360), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n690), .B1(new_n481), .B2(new_n700), .ZN(G1328gat));
  NOR2_X1   g500(.A1(new_n453), .A2(G36gat), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n688), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n688), .A2(KEYINPUT102), .A3(new_n702), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT103), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n706), .B1(new_n705), .B2(new_n707), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n430), .A3(new_n699), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(G36gat), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n712), .ZN(G1329gat));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n693), .B1(new_n465), .B2(new_n635), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n681), .ZN(new_n716));
  INV_X1    g515(.A(new_n306), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .A4(new_n699), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G43gat), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n674), .A2(G43gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n688), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n683), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n691), .A2(new_n543), .A3(new_n723), .A4(new_n721), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT105), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n719), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(G43gat), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n718), .B2(KEYINPUT106), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n695), .A2(new_n732), .A3(new_n717), .A4(new_n699), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n720), .B1(new_n688), .B2(new_n721), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n724), .A2(KEYINPUT105), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT47), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n714), .B(new_n729), .C1(new_n734), .C2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n733), .B2(new_n731), .ZN(new_n739));
  INV_X1    g538(.A(new_n728), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n719), .B2(new_n726), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT107), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n742), .ZN(G1330gat));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n715), .A2(new_n716), .A3(new_n424), .A4(new_n699), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n744), .B1(new_n746), .B2(KEYINPUT109), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n424), .A2(new_n393), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT108), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n745), .A2(G50gat), .B1(new_n688), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n747), .B(new_n750), .ZN(G1331gat));
  NOR3_X1   g550(.A1(new_n636), .A2(new_n697), .A3(new_n682), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(new_n691), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n360), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n691), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT110), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n430), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n759));
  XOR2_X1   g558(.A(KEYINPUT49), .B(G64gat), .Z(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n758), .B2(new_n760), .ZN(G1333gat));
  NAND3_X1  g560(.A1(new_n757), .A2(G71gat), .A3(new_n717), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n558), .B1(new_n756), .B2(new_n674), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT50), .ZN(G1334gat));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n757), .A2(new_n766), .A3(new_n424), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n753), .A2(KEYINPUT110), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n756), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n424), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT112), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT111), .B(G78gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1335gat));
  NOR2_X1   g574(.A1(new_n595), .A2(new_n697), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n691), .A2(new_n681), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n691), .A2(KEYINPUT51), .A3(new_n681), .A4(new_n776), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(new_n781), .B2(new_n780), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n360), .A2(new_n605), .A3(new_n661), .ZN(new_n784));
  INV_X1    g583(.A(new_n695), .ZN(new_n785));
  INV_X1    g584(.A(new_n776), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n682), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n785), .A2(new_n452), .A3(new_n788), .ZN(new_n789));
  OAI22_X1  g588(.A1(new_n783), .A2(new_n784), .B1(new_n789), .B2(new_n605), .ZN(G1336gat));
  NAND4_X1  g589(.A1(new_n715), .A2(new_n716), .A3(new_n430), .A4(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G92gat), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n453), .A2(G92gat), .A3(new_n682), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n792), .B(new_n793), .C1(new_n783), .C2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n779), .B2(new_n780), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n792), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT52), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(G1337gat));
  INV_X1    g601(.A(G99gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n673), .A2(new_n803), .A3(new_n661), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n785), .A2(new_n306), .A3(new_n788), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n783), .A2(new_n804), .B1(new_n805), .B2(new_n803), .ZN(G1338gat));
  OR3_X1    g605(.A1(new_n461), .A2(G106gat), .A3(new_n682), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n783), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n695), .A2(new_n424), .A3(new_n787), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G106gat), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n779), .A2(new_n780), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n807), .B(KEYINPUT116), .Z(new_n814));
  AOI22_X1  g613(.A1(new_n809), .A2(G106gat), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI22_X1  g614(.A1(new_n808), .A2(new_n812), .B1(new_n811), .B2(new_n815), .ZN(G1339gat));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n655), .B1(new_n659), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n643), .A2(new_n658), .A3(new_n647), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT117), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n643), .A2(new_n647), .A3(new_n821), .A4(new_n658), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n817), .B1(new_n648), .B2(new_n649), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n823), .A2(KEYINPUT118), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT118), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n818), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(KEYINPUT55), .B(new_n818), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n829), .A2(new_n697), .A3(new_n656), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n527), .A2(new_n535), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n511), .A2(new_n514), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n513), .B1(new_n525), .B2(new_n510), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n832), .B1(new_n533), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n661), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n681), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n836), .A2(new_n632), .A3(new_n634), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n839), .A2(new_n829), .A3(new_n656), .A4(new_n830), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n680), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n595), .A2(new_n698), .A3(new_n635), .A4(new_n682), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(new_n462), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n452), .A2(new_n430), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n543), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n847), .A2(new_n848), .A3(G113gat), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n847), .B2(G113gat), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n302), .A2(new_n456), .A3(new_n304), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n844), .A2(new_n360), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT120), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n844), .A2(new_n854), .A3(new_n360), .A4(new_n851), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n453), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n697), .A2(new_n253), .ZN(new_n858));
  OAI22_X1  g657(.A1(new_n849), .A2(new_n850), .B1(new_n857), .B2(new_n858), .ZN(G1340gat));
  NAND2_X1  g658(.A1(new_n845), .A2(new_n846), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(new_n251), .A3(new_n682), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n856), .A2(new_n453), .A3(new_n661), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n251), .ZN(G1341gat));
  INV_X1    g662(.A(G127gat), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n860), .A2(new_n864), .A3(new_n680), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n430), .B(new_n680), .C1(new_n853), .C2(new_n855), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867));
  AOI21_X1  g666(.A(G127gat), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT121), .B1(new_n857), .B2(new_n680), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(G1342gat));
  OAI21_X1  g669(.A(G134gat), .B1(new_n860), .B2(new_n635), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n635), .A2(new_n430), .A3(G134gat), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n873), .B1(new_n853), .B2(new_n855), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT122), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n874), .A2(new_n875), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n874), .A2(new_n875), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .A4(new_n871), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n882), .ZN(G1343gat));
  NAND2_X1  g682(.A1(new_n306), .A2(new_n846), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n461), .B1(new_n842), .B2(new_n843), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n829), .A2(new_n543), .A3(new_n656), .A4(new_n830), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n681), .B1(new_n888), .B2(new_n837), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n840), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n680), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n461), .B1(new_n893), .B2(new_n843), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n887), .B1(new_n894), .B2(new_n886), .ZN(new_n895));
  OAI21_X1  g694(.A(G141gat), .B1(new_n895), .B2(new_n544), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n306), .A2(new_n424), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n430), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n844), .A2(new_n898), .A3(new_n360), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n899), .A2(G141gat), .A3(new_n544), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(KEYINPUT58), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n697), .B(new_n887), .C1(new_n894), .C2(new_n886), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n900), .B1(new_n904), .B2(G141gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n902), .B1(new_n903), .B2(new_n905), .ZN(G1344gat));
  INV_X1    g705(.A(G148gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(KEYINPUT59), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(new_n895), .B2(new_n682), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n886), .B1(new_n844), .B2(new_n424), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n461), .A2(KEYINPUT57), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n680), .B1(new_n889), .B2(new_n841), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n595), .A2(new_n544), .A3(new_n635), .A4(new_n682), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR4_X1   g714(.A1(new_n910), .A2(new_n682), .A3(new_n915), .A4(new_n884), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT59), .B1(new_n916), .B2(new_n907), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n909), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n899), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n907), .A3(new_n661), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1345gat));
  OAI21_X1  g720(.A(G155gat), .B1(new_n895), .B2(new_n680), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n315), .A3(new_n595), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1346gat));
  INV_X1    g723(.A(new_n319), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n895), .B2(new_n635), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n319), .A3(new_n681), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n360), .A2(new_n453), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT124), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n845), .A2(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(new_n231), .A3(new_n544), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n360), .B1(new_n842), .B2(new_n843), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n851), .A2(new_n430), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n697), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n933), .A2(new_n938), .ZN(G1348gat));
  OAI21_X1  g738(.A(G176gat), .B1(new_n932), .B2(new_n682), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n937), .A2(new_n232), .A3(new_n661), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1349gat));
  INV_X1    g741(.A(new_n932), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n209), .B1(new_n943), .B2(new_n595), .ZN(new_n944));
  NOR4_X1   g743(.A1(new_n936), .A2(new_n218), .A3(new_n219), .A4(new_n680), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n944), .A2(new_n945), .A3(KEYINPUT60), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT60), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1350gat));
  NAND3_X1  g747(.A1(new_n937), .A2(new_n211), .A3(new_n681), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n943), .A2(new_n681), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(G190gat), .ZN(new_n952));
  AOI211_X1 g751(.A(KEYINPUT61), .B(new_n211), .C1(new_n943), .C2(new_n681), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(G1351gat));
  AND4_X1   g753(.A1(new_n306), .A2(new_n934), .A3(new_n424), .A4(new_n430), .ZN(new_n955));
  XNOR2_X1  g754(.A(KEYINPUT125), .B(G197gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n697), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT126), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n913), .A2(new_n914), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(new_n911), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n717), .A2(new_n930), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n960), .B(new_n961), .C1(new_n886), .C2(new_n885), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n962), .A2(new_n544), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n958), .B1(new_n963), .B2(new_n956), .ZN(G1352gat));
  NAND3_X1  g763(.A1(new_n955), .A2(new_n367), .A3(new_n661), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT62), .Z(new_n966));
  OAI21_X1  g765(.A(G204gat), .B1(new_n962), .B2(new_n682), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n955), .A2(new_n371), .A3(new_n595), .ZN(new_n969));
  INV_X1    g768(.A(new_n961), .ZN(new_n970));
  NOR4_X1   g769(.A1(new_n910), .A2(new_n680), .A3(new_n915), .A4(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n371), .B1(new_n971), .B2(KEYINPUT127), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n973), .B1(new_n962), .B2(new_n680), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n844), .A2(new_n424), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n915), .B1(new_n976), .B2(KEYINPUT57), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n977), .A2(KEYINPUT127), .A3(new_n595), .A4(new_n961), .ZN(new_n978));
  AND4_X1   g777(.A1(KEYINPUT63), .A2(new_n974), .A3(G211gat), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n969), .B1(new_n975), .B2(new_n979), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n962), .B2(new_n635), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n955), .A2(new_n372), .A3(new_n681), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


