//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1240;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  OR2_X1    g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(new_n464), .A2(new_n471), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n470), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G138), .B(new_n471), .C1(new_n462), .C2(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .A3(G138), .A4(new_n471), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n486), .A2(G126), .A3(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n485), .A2(new_n487), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G164));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G651), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n495));
  INV_X1    g070(.A(G651), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(KEYINPUT6), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(KEYINPUT67), .A3(G651), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G50), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n498), .ZN(new_n503));
  INV_X1    g078(.A(new_n494), .ZN(new_n504));
  OR2_X1    g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G88), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n511), .A2(new_n496), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n502), .A2(new_n510), .A3(new_n512), .ZN(G166));
  NAND3_X1  g088(.A1(new_n499), .A2(G89), .A3(new_n507), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n499), .A2(G51), .A3(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(G63), .A2(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT7), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n519), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n507), .A2(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n514), .A2(new_n515), .A3(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  INV_X1    g098(.A(G64), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n524), .B1(new_n505), .B2(new_n506), .ZN(new_n525));
  AND2_X1   g100(.A1(G77), .A2(G543), .ZN(new_n526));
  OAI21_X1  g101(.A(G651), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n503), .A2(G90), .A3(new_n507), .A4(new_n504), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n503), .A2(G52), .A3(G543), .A4(new_n504), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT68), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(G171));
  INV_X1    g109(.A(G56), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(new_n505), .B2(new_n506), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n537));
  AND2_X1   g112(.A1(G68), .A2(G543), .ZN(new_n538));
  OR3_X1    g113(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(G651), .A3(new_n540), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n503), .A2(G43), .A3(G543), .A4(new_n504), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n503), .A2(G81), .A3(new_n507), .A4(new_n504), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT70), .ZN(new_n544));
  AOI21_X1  g119(.A(KEYINPUT70), .B1(new_n542), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT71), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT72), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(new_n554));
  XOR2_X1   g129(.A(new_n554), .B(KEYINPUT73), .Z(G188));
  NAND2_X1  g130(.A1(new_n508), .A2(KEYINPUT75), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n499), .A2(new_n557), .A3(new_n507), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(G91), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT74), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n562), .B1(new_n563), .B2(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n501), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n496), .ZN(new_n567));
  OAI211_X1 g142(.A(KEYINPUT74), .B(new_n560), .C1(new_n500), .C2(new_n562), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n559), .A2(new_n565), .A3(new_n567), .A4(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  NAND3_X1  g145(.A1(new_n502), .A2(new_n512), .A3(new_n510), .ZN(G303));
  OR2_X1    g146(.A1(new_n507), .A2(G74), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n501), .A2(G49), .B1(G651), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n556), .A2(G87), .A3(new_n558), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT76), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n573), .A2(new_n577), .A3(new_n574), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G288));
  AND4_X1   g155(.A1(new_n557), .A2(new_n503), .A3(new_n504), .A4(new_n507), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n557), .B1(new_n499), .B2(new_n507), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G86), .ZN(new_n584));
  AND2_X1   g159(.A1(G48), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n499), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n499), .A2(KEYINPUT77), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(new_n507), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n588), .A2(new_n589), .B1(new_n593), .B2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n584), .A2(new_n594), .ZN(G305));
  XNOR2_X1  g170(.A(KEYINPUT78), .B(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n501), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n496), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n509), .A2(G85), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(G290));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NOR2_X1   g177(.A1(G301), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n591), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G651), .ZN(new_n607));
  INV_X1    g182(.A(G54), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n500), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n556), .A2(G92), .A3(new_n558), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n556), .A2(KEYINPUT10), .A3(G92), .A4(new_n558), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT79), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(KEYINPUT80), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n614), .B(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n603), .B1(new_n621), .B2(new_n602), .ZN(G284));
  AOI21_X1  g197(.A(new_n603), .B1(new_n621), .B2(new_n602), .ZN(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  INV_X1    g199(.A(G299), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n621), .A2(new_n630), .A3(new_n628), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n630), .B1(new_n621), .B2(new_n628), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n632), .A2(new_n602), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n602), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n486), .A2(new_n472), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT82), .B(G2100), .Z(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n476), .A2(G123), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n470), .A2(G135), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n471), .A2(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G2096), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n641), .A2(new_n642), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2443), .B(G2446), .Z(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(G14), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n661), .ZN(G401));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(KEYINPUT17), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT84), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n671), .B2(KEYINPUT18), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(new_n648), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n685), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT20), .Z(new_n689));
  AOI211_X1 g264(.A(new_n687), .B(new_n689), .C1(new_n682), .C2(new_n686), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  MUX2_X1   g272(.A(G6), .B(G305), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT86), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT32), .B(G1981), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1971), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n704), .A2(G23), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n575), .B2(G16), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT33), .B(G1976), .Z(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n709), .A2(new_n711), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n707), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n702), .A2(new_n703), .A3(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n704), .A2(G24), .ZN(new_n718));
  INV_X1    g293(.A(G290), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n704), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1986), .Z(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n476), .A2(G119), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n470), .A2(G131), .ZN(new_n725));
  OR2_X1    g300(.A1(G95), .A2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n723), .B1(new_n729), .B2(new_n722), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT35), .B(G1991), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT85), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n716), .A2(new_n717), .A3(new_n721), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT36), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT87), .ZN(new_n736));
  OR3_X1    g311(.A1(new_n736), .A2(G4), .A3(G16), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(G4), .B2(G16), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n616), .A2(new_n620), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n737), .B(new_n738), .C1(new_n739), .C2(new_n704), .ZN(new_n740));
  INV_X1    g315(.A(G1348), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n476), .A2(G129), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n472), .A2(G105), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G141), .B2(new_n470), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT90), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT26), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(new_n722), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n722), .B2(G32), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n722), .A2(G35), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G162), .B2(new_n722), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT29), .B(G2090), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n755), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n722), .A2(G27), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G164), .B2(new_n722), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2078), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n722), .A2(G26), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT28), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n476), .A2(G128), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n470), .A2(G140), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n471), .A2(G116), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n767), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n766), .B1(new_n771), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2067), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT31), .B(G11), .Z(new_n774));
  INV_X1    g349(.A(G28), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT30), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(KEYINPUT30), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n773), .B(new_n778), .C1(new_n722), .C2(new_n647), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n761), .A2(new_n764), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n547), .A2(G16), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G16), .B2(G19), .ZN(new_n782));
  INV_X1    g357(.A(G1341), .ZN(new_n783));
  NOR2_X1   g358(.A1(G171), .A2(new_n704), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G5), .B2(new_n704), .ZN(new_n785));
  INV_X1    g360(.A(G1961), .ZN(new_n786));
  OAI22_X1  g361(.A1(new_n782), .A2(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n786), .B2(new_n785), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n722), .A2(G33), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT25), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n470), .A2(G139), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(G115), .A2(G2104), .ZN(new_n794));
  INV_X1    g369(.A(G127), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n464), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n791), .B(new_n793), .C1(G2105), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT88), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n789), .B1(new_n798), .B2(new_n722), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G2072), .Z(new_n800));
  INV_X1    g375(.A(G34), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n801), .A2(KEYINPUT24), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(KEYINPUT24), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n722), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G160), .B2(new_n722), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT89), .Z(new_n806));
  INV_X1    g381(.A(G2084), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n704), .A2(G21), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G168), .B2(new_n704), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G1966), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(G1966), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n808), .A2(new_n809), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n783), .B2(new_n782), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n780), .A2(new_n788), .A3(new_n800), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n704), .A2(G20), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT23), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n625), .B2(new_n704), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT91), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(G1956), .Z(new_n821));
  NOR3_X1   g396(.A1(new_n742), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n735), .A2(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  NAND2_X1  g399(.A1(new_n621), .A2(G559), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT38), .Z(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n505), .B2(new_n506), .ZN(new_n828));
  AND2_X1   g403(.A1(G80), .A2(G543), .ZN(new_n829));
  OAI21_X1  g404(.A(G651), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n503), .A2(G93), .A3(new_n507), .A4(new_n504), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n503), .A2(G55), .A3(G543), .A4(new_n504), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT92), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n546), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n542), .A2(new_n543), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT70), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT70), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n843), .A2(new_n541), .B1(new_n834), .B2(new_n836), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n826), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n826), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(G860), .B1(new_n848), .B2(KEYINPUT39), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n846), .A2(new_n850), .A3(new_n847), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT93), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n849), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n833), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(new_n798), .B(new_n750), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n638), .B(new_n728), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n771), .B(new_n491), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n476), .A2(G130), .B1(G142), .B2(new_n470), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n471), .A2(KEYINPUT94), .A3(G118), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT94), .B1(new_n471), .B2(G118), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n865), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n862), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n861), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n647), .B(new_n474), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n481), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(G37), .B1(new_n869), .B2(new_n871), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  OAI22_X1  g450(.A1(new_n632), .A2(new_n633), .B1(new_n838), .B2(new_n844), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT81), .B1(new_n739), .B2(G559), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n877), .A2(new_n631), .A3(new_n845), .ZN(new_n878));
  INV_X1    g453(.A(new_n609), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT10), .B1(new_n583), .B2(G92), .ZN(new_n880));
  INV_X1    g455(.A(new_n613), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n625), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT95), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n612), .A2(new_n613), .ZN(new_n885));
  AND4_X1   g460(.A1(new_n884), .A2(new_n885), .A3(G299), .A4(new_n879), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n614), .B2(G299), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n876), .A2(new_n878), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n885), .A2(G299), .A3(new_n879), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n614), .A2(G299), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n891), .B1(new_n882), .B2(new_n625), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n886), .B2(new_n887), .ZN(new_n897));
  AOI22_X1  g472(.A1(new_n876), .A2(new_n878), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(G166), .A2(new_n575), .ZN(new_n899));
  NAND3_X1  g474(.A1(G303), .A2(new_n574), .A3(new_n573), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(G290), .A2(new_n584), .A3(new_n594), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(G290), .B1(new_n584), .B2(new_n594), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(G305), .A2(new_n719), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n906), .A2(new_n900), .A3(new_n899), .A4(new_n902), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(KEYINPUT96), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(KEYINPUT42), .Z(new_n910));
  NOR3_X1   g485(.A1(new_n890), .A2(new_n898), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n910), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n876), .A2(new_n878), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n897), .A2(new_n895), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n912), .B1(new_n915), .B2(new_n889), .ZN(new_n916));
  OAI21_X1  g491(.A(G868), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n833), .A2(new_n602), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(G295));
  OAI21_X1  g494(.A(new_n910), .B1(new_n890), .B2(new_n898), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n915), .A2(new_n889), .A3(new_n912), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n602), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n918), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT97), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT97), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n917), .A2(new_n925), .A3(new_n918), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(G331));
  AOI21_X1  g502(.A(G168), .B1(new_n531), .B2(new_n533), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n531), .A2(G168), .A3(new_n533), .ZN(new_n929));
  OAI22_X1  g504(.A1(new_n838), .A2(new_n844), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n843), .A2(new_n541), .A3(new_n834), .A4(new_n836), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n546), .A2(new_n837), .ZN(new_n932));
  NAND2_X1  g507(.A1(G171), .A2(G286), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n531), .A2(G168), .A3(new_n533), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n891), .B1(new_n930), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n883), .A2(new_n892), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n908), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND4_X1   g513(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n934), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n931), .A2(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT41), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n892), .A2(KEYINPUT95), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n614), .A2(new_n884), .A3(G299), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n894), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n938), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n930), .A2(new_n935), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n897), .A2(new_n947), .A3(new_n895), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n942), .A2(new_n943), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n949), .A2(new_n883), .A3(new_n935), .A4(new_n930), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n908), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n946), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G37), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n905), .A2(new_n907), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n948), .A2(new_n956), .A3(new_n950), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n952), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n954), .B1(new_n958), .B2(new_n953), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n937), .B(KEYINPUT41), .C1(new_n939), .C2(new_n940), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n956), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n936), .A2(new_n888), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n955), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n956), .B1(new_n948), .B2(new_n950), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT98), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT98), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n946), .A2(new_n952), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n969), .A3(KEYINPUT43), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT99), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n967), .A2(new_n969), .A3(KEYINPUT99), .A4(KEYINPUT43), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n952), .A2(new_n953), .A3(new_n957), .A4(new_n955), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT44), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  AND4_X1   g551(.A1(KEYINPUT100), .A2(new_n972), .A3(new_n973), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n970), .B2(new_n971), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT100), .B1(new_n978), .B2(new_n973), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n961), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT101), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT101), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n982), .B(new_n961), .C1(new_n977), .C2(new_n979), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(G397));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n491), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT108), .ZN(new_n989));
  INV_X1    g564(.A(G2090), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n467), .A2(G40), .A3(new_n473), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n491), .A2(new_n987), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n986), .B1(new_n491), .B2(new_n987), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n996), .A2(KEYINPUT107), .A3(new_n991), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n989), .B(new_n990), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n991), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n491), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT102), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n491), .A2(KEYINPUT102), .A3(KEYINPUT45), .A4(new_n987), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1971), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n998), .A2(KEYINPUT109), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT109), .B1(new_n998), .B2(new_n1007), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G303), .A2(G8), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT103), .B(KEYINPUT55), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n985), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n998), .A2(new_n1007), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n998), .A2(KEYINPUT109), .A3(new_n1007), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(G8), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(KEYINPUT110), .A3(new_n1014), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1016), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT121), .ZN(new_n1024));
  INV_X1    g599(.A(G2078), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1000), .A2(new_n1003), .A3(new_n1025), .A4(new_n1004), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n1029));
  INV_X1    g604(.A(new_n991), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n1030), .A3(new_n988), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n786), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1027), .A2(G2078), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1000), .A2(new_n1003), .A3(new_n1004), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1024), .B1(new_n1028), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1037), .A2(KEYINPUT121), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(G171), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1001), .A2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n491), .A2(KEYINPUT112), .A3(KEYINPUT45), .A4(new_n987), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1000), .A2(new_n1041), .A3(new_n1042), .A4(new_n1033), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1037), .A2(G301), .A3(new_n1032), .A4(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1044), .A2(KEYINPUT54), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT122), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT122), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1039), .A2(new_n1048), .A3(new_n1045), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n992), .A2(new_n991), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n1010), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n509), .A2(G86), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n594), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(G1981), .ZN(new_n1056));
  INV_X1    g631(.A(G1981), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n584), .A2(new_n1057), .A3(new_n594), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT49), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1053), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1056), .A2(KEYINPUT49), .A3(new_n1058), .ZN(new_n1062));
  INV_X1    g637(.A(G1976), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT104), .B1(new_n575), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT104), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n573), .A2(new_n1065), .A3(new_n574), .A4(G1976), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(new_n1052), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1061), .A2(new_n1062), .B1(KEYINPUT52), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1052), .A2(new_n1066), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n576), .A2(new_n1063), .A3(new_n578), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1064), .A4(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1069), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1058), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1057), .B1(new_n594), .B2(new_n1054), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1060), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(new_n1052), .A3(new_n1062), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1067), .A2(KEYINPUT52), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1073), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT111), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n993), .A2(new_n990), .A3(new_n988), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1010), .B1(new_n1007), .B2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1074), .A2(new_n1081), .B1(new_n1015), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1032), .A2(new_n1043), .ZN(new_n1086));
  AOI21_X1  g661(.A(G301), .B1(new_n1086), .B2(new_n1037), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1028), .A2(new_n1035), .A3(G171), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT120), .B(new_n1085), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1023), .A2(new_n1050), .A3(new_n1084), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1000), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1095));
  INV_X1    g670(.A(G1966), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n993), .A2(new_n807), .A3(new_n988), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(G168), .A2(new_n1010), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT118), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1010), .B1(new_n1108), .B2(new_n1100), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1105), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1110), .B(G8), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT51), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1107), .A2(G8), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(new_n1105), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1106), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT123), .B1(new_n1094), .B2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(G299), .B(KEYINPUT57), .Z(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  OR2_X1    g696(.A1(new_n1121), .A2(KEYINPUT115), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1005), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT108), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n988), .B(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n995), .ZN(new_n1128));
  INV_X1    g703(.A(new_n997), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1125), .B1(new_n1130), .B2(G1956), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1121), .A2(KEYINPUT115), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1122), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1125), .B(new_n1120), .C1(new_n1130), .C2(G1956), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(KEYINPUT61), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1131), .A2(new_n1121), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT61), .B1(new_n1136), .B2(new_n1134), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  INV_X1    g713(.A(G2067), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1031), .A2(new_n741), .B1(new_n1139), .B2(new_n1051), .ZN(new_n1140));
  OR3_X1    g715(.A1(new_n615), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n615), .B2(new_n1138), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1141), .A2(new_n1142), .B1(new_n1138), .B2(new_n615), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT58), .B(G1341), .Z(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n992), .B2(new_n991), .ZN(new_n1147));
  INV_X1    g722(.A(G1996), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1123), .A2(KEYINPUT116), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT116), .B1(new_n1123), .B2(new_n1148), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1147), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT117), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1153), .B(new_n1147), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1145), .B1(new_n1155), .B2(new_n547), .ZN(new_n1156));
  AOI211_X1 g731(.A(KEYINPUT59), .B(new_n546), .C1(new_n1152), .C2(new_n1154), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1135), .B(new_n1144), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n615), .A2(new_n1140), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1134), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1158), .A2(new_n1133), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(G8), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1104), .B1(new_n1162), .B2(KEYINPUT119), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1116), .B1(new_n1163), .B2(new_n1112), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1117), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n1164), .A2(new_n1165), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1083), .A2(new_n1015), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1069), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1169));
  AND4_X1   g744(.A1(new_n1069), .A2(new_n1078), .A3(new_n1073), .A4(new_n1079), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1047), .A2(new_n1049), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1166), .A2(new_n1167), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1119), .A2(new_n1161), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1078), .A2(new_n1063), .A3(new_n579), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1058), .B(KEYINPUT106), .Z(new_n1177));
  AND2_X1   g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1052), .B(KEYINPUT105), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  OAI22_X1  g755(.A1(new_n1178), .A2(new_n1180), .B1(new_n1168), .B2(new_n1080), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1115), .A2(G286), .ZN(new_n1183));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n1172), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1080), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1083), .A2(new_n1015), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT63), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1083), .B2(new_n1015), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1185), .A2(new_n1186), .A3(new_n1183), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(KEYINPUT113), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1080), .A2(G286), .A3(new_n1115), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT113), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1191), .A2(new_n1192), .A3(new_n1188), .A4(new_n1186), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  OAI211_X1 g769(.A(KEYINPUT114), .B(new_n1182), .C1(new_n1184), .C2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT114), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1022), .ZN(new_n1197));
  AOI21_X1  g772(.A(KEYINPUT110), .B1(new_n1021), .B2(new_n1014), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1084), .B(new_n1183), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1194), .B1(new_n1199), .B2(new_n1187), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1196), .B1(new_n1200), .B2(new_n1181), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1166), .A2(KEYINPUT62), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1118), .A2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1202), .A2(new_n1204), .A3(new_n1087), .A4(new_n1172), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1175), .A2(new_n1195), .A3(new_n1201), .A4(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n992), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1207), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n750), .B(new_n1148), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n771), .B(new_n1139), .ZN(new_n1210));
  OR2_X1    g785(.A1(new_n729), .A2(new_n731), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n729), .A2(new_n731), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g788(.A(G290), .B(G1986), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1208), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1206), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1208), .A2(new_n1148), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT46), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  XOR2_X1   g794(.A(new_n1219), .B(KEYINPUT124), .Z(new_n1220));
  INV_X1    g795(.A(new_n1208), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1221), .B1(new_n751), .B2(new_n1210), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1222), .B1(new_n1218), .B2(new_n1217), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g799(.A(new_n1224), .B(KEYINPUT47), .ZN(new_n1225));
  NAND4_X1  g800(.A1(new_n1209), .A2(new_n729), .A3(new_n731), .A4(new_n1210), .ZN(new_n1226));
  OR2_X1    g801(.A1(new_n771), .A2(G2067), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1221), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  OR3_X1    g803(.A1(new_n1221), .A2(G1986), .A3(G290), .ZN(new_n1229));
  INV_X1    g804(.A(new_n1229), .ZN(new_n1230));
  AOI22_X1  g805(.A1(KEYINPUT48), .A2(new_n1230), .B1(new_n1213), .B2(new_n1208), .ZN(new_n1231));
  OR2_X1    g806(.A1(new_n1230), .A2(KEYINPUT48), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1228), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1225), .A2(new_n1233), .ZN(new_n1234));
  XOR2_X1   g809(.A(new_n1234), .B(KEYINPUT125), .Z(new_n1235));
  NAND2_X1  g810(.A1(new_n1216), .A2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g811(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1238));
  NAND4_X1  g812(.A1(new_n874), .A2(new_n696), .A3(new_n959), .A4(new_n1238), .ZN(G225));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1240));
  XNOR2_X1  g814(.A(G225), .B(new_n1240), .ZN(G308));
endmodule


