//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT75), .B(G125), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n189), .A3(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(G125), .A2(G140), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n192), .B1(new_n188), .B2(G140), .ZN(new_n193));
  OAI211_X1 g007(.A(G146), .B(new_n191), .C1(new_n193), .C2(new_n189), .ZN(new_n194));
  XNOR2_X1  g008(.A(G125), .B(G140), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  OR2_X1    g013(.A1(KEYINPUT69), .A2(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT69), .A2(G128), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n199), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT23), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT69), .A2(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT69), .A2(G128), .ZN(new_n206));
  OAI211_X1 g020(.A(KEYINPUT23), .B(G119), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT74), .ZN(new_n208));
  INV_X1    g022(.A(G110), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT23), .B1(new_n210), .B2(G119), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(G119), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n204), .A2(new_n208), .A3(new_n209), .A4(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n202), .A2(new_n212), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT24), .B(G110), .Z(new_n216));
  OR2_X1    g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n198), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G125), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT75), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT75), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G125), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n222), .A3(G140), .ZN(new_n223));
  INV_X1    g037(.A(new_n192), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n189), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AND4_X1   g039(.A1(new_n189), .A2(new_n220), .A3(new_n222), .A4(new_n190), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n196), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n194), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n204), .A2(new_n213), .A3(new_n208), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G110), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n215), .A2(new_n216), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT76), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n227), .A2(new_n194), .B1(new_n215), .B2(new_n216), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT76), .A3(new_n230), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n218), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  INV_X1    g052(.A(G221), .ZN(new_n239));
  INV_X1    g053(.A(G953), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT72), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G953), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n239), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT22), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(G234), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n245), .B1(new_n244), .B2(G234), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n238), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n248), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(G137), .A3(new_n246), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT77), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT77), .B1(new_n249), .B2(new_n251), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n237), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n249), .A2(new_n251), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI211_X1 g071(.A(new_n218), .B(new_n257), .C1(new_n234), .C2(new_n236), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n187), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT25), .ZN(new_n260));
  INV_X1    g074(.A(G217), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(G234), .B2(new_n187), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n234), .A2(new_n236), .ZN(new_n263));
  INV_X1    g077(.A(new_n218), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(new_n256), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n237), .B2(new_n254), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT25), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n187), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n260), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n262), .A2(G902), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(G101), .ZN(new_n274));
  AOI21_X1  g088(.A(G237), .B1(new_n241), .B2(new_n243), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G210), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n274), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT2), .B(G113), .Z(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(G116), .B(G119), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n280), .A2(new_n282), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT71), .ZN(new_n286));
  OR3_X1    g100(.A1(new_n280), .A2(KEYINPUT71), .A3(new_n282), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G131), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n291));
  INV_X1    g105(.A(G134), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT66), .A2(G134), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n238), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(G137), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n290), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT11), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT11), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT65), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n238), .A2(KEYINPUT11), .A3(G134), .ZN(new_n304));
  AND2_X1   g118(.A1(KEYINPUT66), .A2(G134), .ZN(new_n305));
  NOR2_X1   g119(.A1(KEYINPUT66), .A2(G134), .ZN(new_n306));
  OAI21_X1  g120(.A(G137), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND4_X1   g121(.A1(new_n290), .A2(new_n303), .A3(new_n304), .A4(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT64), .B1(new_n196), .B2(G143), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT64), .ZN(new_n310));
  INV_X1    g124(.A(G143), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(G146), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT1), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n196), .A2(G143), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n313), .A2(new_n314), .A3(G128), .A4(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT68), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n309), .A2(new_n312), .B1(G143), .B2(new_n196), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n319), .A2(KEYINPUT68), .A3(new_n314), .A4(G128), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n311), .A2(G146), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT70), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n200), .A2(new_n201), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n314), .B1(G143), .B2(new_n196), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT1), .B1(new_n311), .B2(G146), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n200), .A3(new_n201), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n324), .B1(new_n330), .B2(new_n323), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  AOI211_X1 g146(.A(new_n297), .B(new_n308), .C1(new_n321), .C2(new_n332), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n305), .A2(new_n306), .A3(G137), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n304), .B(new_n307), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT67), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G131), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n303), .A2(new_n338), .A3(new_n304), .A4(new_n307), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n313), .A2(G128), .A3(new_n315), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n323), .A2(new_n210), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(KEYINPUT0), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n210), .B1(new_n315), .B2(new_n322), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n345), .A2(KEYINPUT0), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n340), .A2(new_n341), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n289), .B1(new_n333), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n321), .A2(new_n332), .ZN(new_n349));
  INV_X1    g163(.A(new_n297), .ZN(new_n350));
  INV_X1    g164(.A(new_n308), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n347), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n352), .A2(new_n353), .A3(new_n288), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n279), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n279), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n278), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT31), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n297), .B1(new_n321), .B2(new_n332), .ZN(new_n360));
  AOI211_X1 g174(.A(KEYINPUT30), .B(new_n347), .C1(new_n360), .C2(new_n351), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n352), .B2(new_n353), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n289), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n354), .A3(new_n277), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n358), .A2(new_n359), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G472), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n364), .A2(KEYINPUT31), .A3(new_n354), .A4(new_n277), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n366), .A2(new_n367), .A3(new_n187), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT73), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n187), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n372), .A2(new_n366), .A3(new_n373), .A4(new_n367), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT32), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n354), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n288), .B1(new_n352), .B2(new_n353), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT28), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n277), .A3(new_n356), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n277), .B1(new_n364), .B2(new_n354), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n187), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n381), .A2(new_n382), .ZN(new_n386));
  OAI21_X1  g200(.A(G472), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n372), .A2(new_n366), .A3(KEYINPUT32), .A4(new_n367), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n272), .B1(new_n377), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G113), .B(G122), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G237), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n242), .A2(G953), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n240), .A2(KEYINPUT72), .ZN(new_n396));
  OAI211_X1 g210(.A(G214), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(KEYINPUT93), .A3(G143), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT93), .A2(G143), .ZN(new_n399));
  OR2_X1    g213(.A1(KEYINPUT93), .A2(G143), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n275), .A2(G214), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n290), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT18), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n398), .A2(KEYINPUT18), .A3(new_n401), .A4(G131), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n193), .A2(G146), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n197), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n403), .A2(new_n405), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT94), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n406), .A2(new_n408), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT94), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n403), .A4(new_n405), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n228), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n398), .A2(KEYINPUT17), .A3(new_n401), .A4(G131), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n402), .B(new_n290), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n415), .B(new_n416), .C1(new_n417), .C2(KEYINPUT17), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n393), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT96), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n418), .A3(new_n393), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT96), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n420), .B(new_n187), .C1(new_n423), .C2(new_n419), .ZN(new_n424));
  MUX2_X1   g238(.A(new_n195), .B(new_n193), .S(KEYINPUT19), .Z(new_n425));
  OAI211_X1 g239(.A(new_n417), .B(new_n194), .C1(G146), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n414), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n393), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(G475), .B1(new_n429), .B2(new_n421), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT95), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n414), .A2(new_n393), .A3(new_n418), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n393), .B1(new_n414), .B2(new_n426), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n430), .A2(new_n434), .A3(new_n435), .A4(new_n187), .ZN(new_n436));
  INV_X1    g250(.A(G475), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(new_n187), .C1(new_n432), .C2(new_n433), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT95), .B1(new_n429), .B2(new_n421), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n438), .B1(new_n439), .B2(KEYINPUT20), .ZN(new_n440));
  AOI221_X4 g254(.A(KEYINPUT97), .B1(G475), .B2(new_n424), .C1(new_n436), .C2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT97), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n436), .A2(new_n440), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n424), .A2(G475), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n325), .A2(G143), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n293), .A2(new_n294), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n311), .A2(G128), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT98), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT80), .B(G107), .ZN(new_n452));
  XNOR2_X1  g266(.A(G116), .B(G122), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT13), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n446), .B1(new_n455), .B2(new_n448), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT13), .B1(new_n311), .B2(G128), .ZN(new_n457));
  OAI21_X1  g271(.A(G134), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n451), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G107), .ZN(new_n460));
  INV_X1    g274(.A(G116), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n461), .A2(G122), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n460), .B1(new_n462), .B2(KEYINPUT14), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT14), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n453), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g279(.A1(new_n463), .A2(new_n465), .B1(new_n452), .B2(new_n453), .ZN(new_n466));
  INV_X1    g280(.A(new_n449), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n447), .B1(new_n446), .B2(new_n448), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(KEYINPUT9), .B(G234), .Z(new_n470));
  AND3_X1   g284(.A1(new_n470), .A2(G217), .A3(new_n240), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n459), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n459), .B2(new_n469), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n187), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G478), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n474), .A2(KEYINPUT99), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT99), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(new_n187), .C1(new_n472), .C2(new_n473), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n479), .B1(new_n483), .B2(new_n478), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n441), .A2(new_n445), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT3), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n392), .B2(KEYINPUT79), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT79), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT3), .ZN(new_n489));
  NOR2_X1   g303(.A1(KEYINPUT80), .A2(G107), .ZN(new_n490));
  AND2_X1   g304(.A1(KEYINPUT80), .A2(G107), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n487), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G101), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n392), .A2(G107), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n460), .A2(G104), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT3), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n495), .B1(new_n452), .B2(G104), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G101), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT81), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT81), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n349), .A2(KEYINPUT10), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n340), .A2(new_n341), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT10), .ZN(new_n507));
  INV_X1    g321(.A(new_n319), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n329), .A2(G128), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n318), .A2(new_n320), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n507), .B1(new_n510), .B2(new_n500), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n492), .A2(new_n494), .A3(new_n496), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G101), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n344), .A2(new_n346), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT4), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(new_n516), .A3(G101), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n504), .A2(new_n506), .A3(new_n511), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n241), .A2(new_n243), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G227), .ZN(new_n521));
  XNOR2_X1  g335(.A(G110), .B(G140), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT86), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n321), .A2(new_n332), .A3(new_n500), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n508), .A2(new_n509), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n500), .B1(new_n321), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n505), .B(new_n526), .C1(new_n527), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT83), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n505), .B1(new_n527), .B2(new_n529), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT12), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n321), .A2(new_n332), .A3(new_n500), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n500), .B2(new_n510), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT83), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n505), .A4(new_n526), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n531), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n519), .A2(new_n540), .A3(new_n523), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n525), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT87), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n504), .A2(new_n511), .A3(new_n518), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n545), .A2(KEYINPUT85), .A3(new_n505), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT85), .B1(new_n545), .B2(new_n505), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n519), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n523), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n525), .A2(new_n539), .A3(KEYINPUT87), .A4(new_n541), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G469), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n187), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n539), .A2(new_n519), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n549), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT84), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n524), .B(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n546), .A2(new_n547), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n556), .B(G469), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(G469), .A2(G902), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n554), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n239), .B1(new_n470), .B2(new_n187), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT78), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT88), .B(KEYINPUT5), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n283), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G113), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n461), .A2(G119), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n568), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n567), .A2(new_n570), .B1(new_n282), .B2(new_n280), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n501), .A2(new_n503), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT89), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n289), .A2(new_n514), .A3(new_n517), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT89), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n501), .A2(new_n575), .A3(new_n503), .A4(new_n571), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(G110), .B(G122), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n573), .A2(new_n574), .A3(new_n578), .A4(new_n576), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(KEYINPUT6), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT6), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n577), .A2(new_n583), .A3(new_n579), .ZN(new_n584));
  INV_X1    g398(.A(new_n188), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n349), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G224), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(G953), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n585), .B1(new_n344), .B2(new_n346), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n586), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n188), .B1(new_n321), .B2(new_n332), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n588), .B1(new_n593), .B2(new_n590), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n582), .A2(new_n584), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT7), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n589), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n592), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n497), .A2(new_n499), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n570), .B(KEYINPUT91), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n282), .A2(KEYINPUT5), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n600), .B(new_n285), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n600), .B2(new_n571), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n578), .B(KEYINPUT90), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT8), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n586), .A2(new_n597), .A3(new_n589), .A4(new_n591), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n599), .A2(new_n581), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n609), .A2(new_n187), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n596), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G210), .B1(G237), .B2(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT92), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n596), .A2(new_n610), .A3(new_n612), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n616), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT92), .ZN(new_n619));
  OAI21_X1  g433(.A(G214), .B1(G237), .B2(G902), .ZN(new_n620));
  INV_X1    g434(.A(G952), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n621), .A2(KEYINPUT100), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(KEYINPUT100), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n240), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(G234), .B2(G237), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  AOI211_X1 g440(.A(new_n187), .B(new_n520), .C1(G234), .C2(G237), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT21), .B(G898), .Z(new_n629));
  OAI21_X1  g443(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n617), .A2(new_n619), .A3(new_n620), .A4(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n390), .A2(new_n485), .A3(new_n565), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G101), .ZN(G3));
  NOR2_X1   g448(.A1(new_n472), .A2(new_n473), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT33), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n636), .A2(new_n476), .A3(G902), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n483), .A2(G478), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT20), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n187), .A2(new_n430), .B1(new_n434), .B2(new_n435), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n444), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT97), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n443), .A2(new_n442), .A3(new_n444), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n639), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n620), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n614), .B2(new_n616), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n630), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n367), .B1(new_n372), .B2(new_n366), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n370), .B2(new_n374), .ZN(new_n652));
  INV_X1    g466(.A(new_n272), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n652), .A2(new_n562), .A3(new_n653), .A4(new_n564), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT34), .B(G104), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  INV_X1    g471(.A(new_n654), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n438), .A2(new_n435), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n430), .A2(KEYINPUT20), .A3(new_n187), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n444), .A2(new_n484), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n648), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  AND3_X1   g480(.A1(new_n358), .A2(new_n359), .A3(new_n365), .ZN(new_n667));
  OAI21_X1  g481(.A(G472), .B1(new_n667), .B2(new_n371), .ZN(new_n668));
  INV_X1    g482(.A(new_n237), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT101), .B1(new_n254), .B2(KEYINPUT36), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n254), .A2(KEYINPUT101), .A3(KEYINPUT36), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n672), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n237), .A3(new_n670), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n673), .A2(new_n675), .A3(new_n270), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n269), .A2(new_n676), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n375), .A2(new_n668), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n485), .A2(new_n565), .A3(new_n678), .A4(new_n632), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT37), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n209), .ZN(G12));
  AOI21_X1  g495(.A(KEYINPUT32), .B1(new_n370), .B2(new_n374), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n387), .A2(new_n388), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n562), .A2(new_n564), .ZN(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n627), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n626), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n661), .A2(new_n647), .A3(new_n677), .A4(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n684), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT102), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  OAI21_X1  g506(.A(new_n278), .B1(new_n378), .B2(new_n379), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n365), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(KEYINPUT103), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(G902), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n694), .A2(KEYINPUT103), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n367), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n377), .A2(new_n388), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n677), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n688), .B(KEYINPUT39), .Z(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n565), .A2(KEYINPUT104), .A3(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(new_n685), .B2(new_n703), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n702), .B1(new_n708), .B2(KEYINPUT40), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n617), .A2(new_n619), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT38), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n484), .B1(new_n441), .B2(new_n445), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT40), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n705), .A2(new_n714), .A3(new_n707), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n709), .A2(new_n620), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  INV_X1    g531(.A(new_n639), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n718), .B(new_n688), .C1(new_n441), .C2(new_n445), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n377), .A2(new_n389), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n647), .A2(new_n677), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n720), .A2(new_n721), .A3(new_n565), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  NAND2_X1  g538(.A1(new_n552), .A2(new_n187), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(G469), .ZN(new_n726));
  INV_X1    g540(.A(new_n563), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n554), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n390), .A2(new_n645), .A3(new_n649), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND4_X1  g546(.A1(new_n721), .A2(new_n663), .A3(new_n729), .A4(new_n653), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  NOR2_X1   g548(.A1(new_n728), .A2(new_n648), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n485), .A3(new_n721), .A4(new_n677), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  INV_X1    g551(.A(new_n484), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n643), .B2(new_n644), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n653), .A2(new_n369), .A3(new_n668), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n735), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  AND4_X1   g556(.A1(new_n554), .A2(new_n726), .A3(new_n727), .A4(new_n647), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n668), .A2(new_n677), .A3(new_n369), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT105), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n668), .A2(new_n677), .A3(KEYINPUT105), .A4(new_n369), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n645), .A2(new_n743), .A3(new_n748), .A4(new_n688), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n646), .B1(new_n617), .B2(new_n619), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT106), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n560), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n524), .B(KEYINPUT84), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n546), .A2(new_n547), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n755), .A2(new_n756), .B1(new_n555), .B2(new_n549), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT106), .A3(G469), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n554), .A2(new_n754), .A3(new_n758), .A4(new_n561), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n759), .A2(new_n727), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n390), .A2(new_n752), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n751), .B1(new_n761), .B2(new_n719), .ZN(new_n762));
  INV_X1    g576(.A(new_n752), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n719), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n369), .A2(new_n376), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT107), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n272), .B1(new_n766), .B2(new_n389), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n764), .A2(new_n767), .A3(KEYINPUT42), .A4(new_n760), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G131), .ZN(G33));
  INV_X1    g584(.A(new_n688), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n662), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n390), .A2(new_n772), .A3(new_n752), .A4(new_n760), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n752), .B(new_n653), .C1(new_n682), .C2(new_n683), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(KEYINPUT108), .A3(new_n772), .A4(new_n760), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n643), .A2(new_n644), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n782), .B2(new_n639), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n441), .A2(new_n445), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(KEYINPUT43), .A3(new_n718), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n652), .B(new_n701), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n763), .B1(new_n786), .B2(KEYINPUT44), .ZN(new_n787));
  INV_X1    g601(.A(new_n554), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n789), .B(G469), .C1(new_n757), .C2(KEYINPUT45), .ZN(new_n790));
  NAND2_X1  g604(.A1(KEYINPUT45), .A2(G469), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n560), .A2(KEYINPUT109), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n757), .A2(KEYINPUT45), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n561), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT46), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n788), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n561), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n563), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT110), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n800), .A3(new_n704), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n797), .A2(new_n798), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n727), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT110), .B1(new_n803), .B2(new_n703), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n783), .A2(new_n785), .ZN(new_n805));
  INV_X1    g619(.A(new_n652), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n806), .A3(new_n677), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n787), .A2(new_n801), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G137), .ZN(G39));
  XNOR2_X1  g625(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n803), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n721), .A2(new_n653), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n799), .A2(new_n812), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n764), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  INV_X1    g632(.A(new_n624), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n805), .A2(new_n625), .A3(new_n740), .ZN(new_n820));
  INV_X1    g634(.A(new_n743), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n820), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n814), .A2(new_n816), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n726), .A2(new_n554), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n564), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n752), .B(new_n823), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT50), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n711), .A2(new_n646), .A3(new_n729), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT115), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n711), .A2(new_n831), .A3(new_n646), .A4(new_n729), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n828), .B1(new_n833), .B2(new_n820), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n823), .A2(KEYINPUT50), .A3(new_n832), .A4(new_n830), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n827), .A2(KEYINPUT51), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n763), .A2(new_n728), .ZN(new_n838));
  INV_X1    g652(.A(new_n388), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n682), .A2(new_n698), .A3(new_n839), .ZN(new_n840));
  AND4_X1   g654(.A1(new_n653), .A2(new_n838), .A3(new_n625), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n784), .A3(new_n639), .ZN(new_n842));
  INV_X1    g656(.A(new_n748), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n805), .A2(new_n625), .A3(new_n838), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT117), .Z(new_n846));
  AOI21_X1  g660(.A(new_n822), .B1(new_n837), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n841), .A2(new_n645), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n730), .A2(new_n736), .A3(new_n741), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n643), .A2(new_n644), .A3(new_n484), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n718), .B1(new_n441), .B2(new_n445), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n658), .A3(new_n632), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n633), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n679), .A2(new_n733), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n849), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n762), .A2(new_n768), .B1(new_n775), .B2(new_n778), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n721), .A2(new_n738), .A3(new_n677), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n444), .A2(new_n659), .A3(new_n660), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n858), .A2(new_n685), .A3(new_n859), .A4(new_n771), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n759), .A2(new_n727), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n843), .A2(new_n719), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n752), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n856), .A2(new_n857), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n721), .A2(new_n565), .A3(new_n772), .A4(new_n722), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n721), .A2(new_n565), .A3(new_n722), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n749), .B(new_n865), .C1(new_n719), .C2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n760), .A2(new_n739), .A3(new_n647), .A4(new_n688), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT52), .B1(new_n868), .B2(new_n702), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT112), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n749), .A2(new_n865), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n484), .B(new_n647), .C1(new_n441), .C2(new_n445), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n873), .A2(new_n771), .A3(new_n861), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n840), .A2(new_n677), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT112), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n871), .A2(new_n876), .A3(new_n877), .A4(new_n723), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n868), .A2(new_n702), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n872), .B1(new_n867), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n870), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT53), .B1(new_n864), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n856), .A2(new_n857), .A3(new_n863), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n874), .A2(new_n875), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n871), .A2(new_n723), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n867), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n885), .A2(new_n872), .B1(new_n886), .B2(new_n876), .ZN(new_n887));
  XNOR2_X1  g701(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n883), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT54), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n769), .A2(new_n779), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n654), .B1(new_n851), .B2(new_n850), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n643), .A2(new_n644), .A3(new_n738), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n685), .A3(new_n631), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n893), .A2(new_n632), .B1(new_n895), .B2(new_n390), .ZN(new_n896));
  INV_X1    g710(.A(new_n650), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n684), .A2(new_n272), .A3(new_n728), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n712), .A2(new_n648), .A3(new_n728), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n897), .A2(new_n898), .B1(new_n899), .B2(new_n740), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n679), .A2(new_n733), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n896), .A2(new_n900), .A3(new_n901), .A4(new_n736), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n892), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(new_n881), .A3(KEYINPUT53), .A4(new_n863), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n889), .B1(new_n883), .B2(new_n887), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n847), .A2(new_n848), .A3(new_n891), .A4(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n845), .B1(new_n834), .B2(new_n835), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n827), .B(KEYINPUT114), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT51), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n805), .A2(new_n625), .A3(new_n767), .A4(new_n838), .ZN(new_n914));
  NOR2_X1   g728(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n914), .B(new_n915), .Z(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(KEYINPUT118), .B2(KEYINPUT48), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n908), .A2(new_n913), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(G952), .A2(G953), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n782), .A2(new_n639), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n711), .A2(new_n920), .A3(new_n653), .A4(new_n620), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n825), .B(KEYINPUT49), .Z(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n564), .A3(new_n840), .ZN(new_n923));
  OAI22_X1  g737(.A1(new_n918), .A2(new_n919), .B1(new_n921), .B2(new_n923), .ZN(G75));
  NAND2_X1  g738(.A1(new_n582), .A2(new_n584), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n595), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT55), .Z(new_n927));
  INV_X1    g741(.A(G210), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n928), .B(new_n187), .C1(new_n904), .C2(new_n905), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n929), .B2(KEYINPUT56), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n187), .B1(new_n904), .B2(new_n905), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(G210), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT56), .ZN(new_n933));
  INV_X1    g747(.A(new_n927), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n520), .A2(G952), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n930), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n930), .A2(new_n935), .A3(KEYINPUT119), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G51));
  NAND2_X1  g756(.A1(new_n561), .A2(KEYINPUT57), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n906), .B1(new_n904), .B2(new_n905), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n561), .A2(KEYINPUT57), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n552), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n794), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n931), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n936), .B1(new_n948), .B2(new_n950), .ZN(G54));
  NAND3_X1  g765(.A1(new_n931), .A2(KEYINPUT58), .A3(G475), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n429), .A2(new_n421), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n952), .A2(new_n954), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n936), .ZN(G60));
  INV_X1    g771(.A(new_n636), .ZN(new_n958));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n958), .B(new_n961), .C1(new_n944), .C2(new_n945), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT120), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n960), .B1(new_n891), .B2(new_n907), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(new_n958), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT53), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n870), .A2(new_n878), .A3(new_n880), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n883), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n880), .B1(new_n867), .B2(new_n869), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n903), .A2(new_n970), .A3(new_n863), .A4(new_n888), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n906), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n961), .B1(new_n944), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(KEYINPUT120), .A3(new_n636), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n936), .B(new_n963), .C1(new_n966), .C2(new_n974), .ZN(G63));
  NAND2_X1  g789(.A1(new_n904), .A2(new_n905), .ZN(new_n976));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT60), .Z(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n266), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n673), .A2(new_n675), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n981), .B(new_n937), .C1(new_n982), .C2(new_n979), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(G66));
  INV_X1    g799(.A(new_n629), .ZN(new_n986));
  OAI21_X1  g800(.A(G953), .B1(new_n986), .B2(new_n587), .ZN(new_n987));
  INV_X1    g801(.A(new_n520), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n987), .B1(new_n856), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT121), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n925), .B1(G898), .B2(new_n520), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(G69));
  INV_X1    g806(.A(KEYINPUT124), .ZN(new_n993));
  INV_X1    g807(.A(G227), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n988), .B1(new_n994), .B2(new_n686), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n361), .A2(new_n363), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(new_n425), .Z(new_n997));
  INV_X1    g811(.A(KEYINPUT122), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n769), .A2(new_n998), .A3(new_n779), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n998), .B1(new_n769), .B2(new_n779), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n810), .B(new_n817), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n873), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n804), .A2(new_n767), .A3(new_n801), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n886), .ZN(new_n1004));
  OAI21_X1  g818(.A(KEYINPUT123), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n810), .A2(new_n817), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT123), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n1003), .A2(new_n886), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1000), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n857), .A2(new_n998), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1011), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n988), .B(new_n997), .C1(new_n1005), .C2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n777), .A2(new_n705), .A3(new_n707), .A4(new_n852), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n805), .A2(KEYINPUT44), .A3(new_n806), .A4(new_n677), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n809), .A2(new_n752), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n804), .A2(new_n801), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n817), .B(new_n1014), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT62), .ZN(new_n1019));
  AND3_X1   g833(.A1(new_n716), .A2(new_n1019), .A3(new_n886), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1019), .B1(new_n716), .B2(new_n886), .ZN(new_n1021));
  NOR3_X1   g835(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n997), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n988), .B1(new_n997), .B2(new_n686), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n993), .B(new_n995), .C1(new_n1013), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1025), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1005), .A2(new_n1012), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n997), .A2(new_n988), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n995), .A2(new_n993), .ZN(new_n1031));
  OR2_X1    g845(.A1(new_n995), .A2(new_n993), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1027), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n1026), .A2(new_n1033), .ZN(G72));
  NAND2_X1  g848(.A1(new_n364), .A2(new_n354), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1035), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n1036), .A2(new_n278), .ZN(new_n1037));
  NOR4_X1   g851(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .A4(new_n902), .ZN(new_n1038));
  XNOR2_X1  g852(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1039));
  NAND2_X1  g853(.A1(G472), .A2(G902), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT126), .Z(new_n1042));
  INV_X1    g856(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1037), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(KEYINPUT127), .ZN(new_n1045));
  INV_X1    g859(.A(KEYINPUT127), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n1046), .B(new_n1037), .C1(new_n1038), .C2(new_n1043), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1005), .A2(new_n1012), .A3(new_n856), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1049), .A2(new_n1042), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1050), .A2(new_n1036), .A3(new_n278), .ZN(new_n1051));
  INV_X1    g865(.A(new_n365), .ZN(new_n1052));
  OAI221_X1 g866(.A(new_n1041), .B1(new_n1052), .B2(new_n384), .C1(new_n882), .C2(new_n890), .ZN(new_n1053));
  AND4_X1   g867(.A1(new_n937), .A2(new_n1048), .A3(new_n1051), .A4(new_n1053), .ZN(G57));
endmodule


