//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT70), .B(G116), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n192), .B1(new_n194), .B2(G119), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT2), .B(G113), .Z(new_n196));
  AND2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n195), .A2(new_n196), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT66), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n203), .A3(G143), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT68), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n204), .A2(new_n210), .A3(new_n205), .A4(new_n207), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G134), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G137), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n215), .A2(new_n222), .A3(new_n216), .A4(new_n219), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n201), .A2(new_n203), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n206), .B2(G146), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n200), .A2(KEYINPUT65), .A3(G143), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n225), .A2(new_n206), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n205), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n229), .A2(KEYINPUT67), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT66), .B(G146), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n200), .A2(KEYINPUT65), .A3(G143), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT65), .B1(new_n200), .B2(G143), .ZN(new_n237));
  OAI22_X1  g051(.A1(new_n235), .A2(G143), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n234), .B1(new_n238), .B2(new_n231), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n212), .B(new_n224), .C1(new_n233), .C2(new_n239), .ZN(new_n240));
  OR2_X1    g054(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n243), .A2(new_n204), .A3(G128), .A4(new_n207), .ZN(new_n244));
  INV_X1    g058(.A(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n242), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n245), .B1(new_n204), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n244), .B1(new_n247), .B2(new_n229), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n218), .A2(G137), .ZN(new_n249));
  OAI21_X1  g063(.A(G131), .B1(new_n249), .B2(new_n214), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n223), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n240), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n199), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n223), .A2(new_n250), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n235), .A2(G143), .B1(new_n241), .B2(new_n242), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n238), .B1(new_n256), .B2(new_n245), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n255), .B1(new_n257), .B2(new_n244), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT67), .B1(new_n229), .B2(new_n232), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n238), .A2(new_n234), .A3(new_n231), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n259), .A2(new_n260), .B1(new_n209), .B2(new_n211), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n258), .B1(new_n261), .B2(new_n224), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT71), .B1(new_n262), .B2(KEYINPUT30), .ZN(new_n263));
  AND4_X1   g077(.A1(KEYINPUT71), .A2(new_n240), .A3(KEYINPUT30), .A4(new_n251), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n254), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT72), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT26), .B(G101), .Z(new_n267));
  INV_X1    g081(.A(G237), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(G210), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n267), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n275), .B(new_n254), .C1(new_n263), .C2(new_n264), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n262), .A2(new_n199), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n266), .A2(new_n274), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n199), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n252), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n199), .B1(new_n240), .B2(new_n251), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT28), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT28), .B1(new_n262), .B2(new_n199), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n278), .A2(KEYINPUT31), .B1(new_n273), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n276), .A2(new_n277), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n274), .A4(new_n266), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n187), .B(new_n189), .C1(new_n286), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n278), .A2(KEYINPUT31), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n285), .A2(new_n273), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT32), .B1(new_n294), .B2(new_n188), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n297));
  INV_X1    g111(.A(G472), .ZN(new_n298));
  INV_X1    g112(.A(new_n281), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n277), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n283), .B1(new_n300), .B2(KEYINPUT28), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT29), .A3(new_n274), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT30), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n305), .B1(new_n252), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n262), .A2(KEYINPUT71), .A3(KEYINPUT30), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n275), .B1(new_n309), .B2(new_n254), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n273), .B1(new_n287), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT29), .B1(new_n301), .B2(new_n274), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n304), .B1(new_n313), .B2(KEYINPUT74), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  AOI211_X1 g130(.A(new_n297), .B(new_n298), .C1(new_n314), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(KEYINPUT74), .ZN(new_n318));
  INV_X1    g132(.A(new_n304), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT75), .B1(new_n320), .B2(G472), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n296), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G475), .ZN(new_n323));
  XNOR2_X1  g137(.A(G125), .B(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT16), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n326), .A2(G140), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(KEYINPUT16), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n200), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n325), .B(G146), .C1(KEYINPUT16), .C2(new_n327), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT80), .B(G143), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n268), .A2(new_n269), .A3(G214), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n268), .A2(new_n269), .A3(G214), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(KEYINPUT80), .B2(new_n206), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT17), .A3(G131), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(G131), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n335), .A2(new_n337), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n222), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n332), .B(new_n339), .C1(new_n343), .C2(KEYINPUT17), .ZN(new_n344));
  XNOR2_X1  g158(.A(G113), .B(G122), .ZN(new_n345));
  INV_X1    g159(.A(G104), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT18), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n341), .B1(new_n348), .B2(new_n222), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n235), .A2(new_n324), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n200), .B2(new_n324), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n349), .B(new_n351), .C1(new_n340), .C2(new_n348), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n344), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n347), .B1(new_n344), .B2(new_n352), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n303), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n323), .B1(new_n356), .B2(KEYINPUT82), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT82), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n358), .B(new_n303), .C1(new_n354), .C2(new_n355), .ZN(new_n359));
  NOR2_X1   g173(.A1(G475), .A2(G902), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n324), .B(KEYINPUT19), .Z(new_n361));
  OAI21_X1  g175(.A(new_n330), .B1(new_n361), .B2(new_n225), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT81), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n330), .B(new_n364), .C1(new_n361), .C2(new_n225), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n343), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n347), .B1(new_n366), .B2(new_n352), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n360), .B1(new_n354), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT20), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT20), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n370), .B(new_n360), .C1(new_n354), .C2(new_n367), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n357), .A2(new_n359), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G952), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G953), .ZN(new_n374));
  NAND2_X1  g188(.A1(G234), .A2(G237), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(G902), .A3(G953), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT21), .B(G898), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT9), .B(G234), .ZN(new_n383));
  INV_X1    g197(.A(G217), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n383), .A2(new_n384), .A3(G953), .ZN(new_n385));
  INV_X1    g199(.A(G122), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G116), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(KEYINPUT83), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n193), .A2(new_n386), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n390), .B2(KEYINPUT14), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G107), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G107), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n390), .A2(new_n395), .A3(new_n388), .ZN(new_n396));
  XNOR2_X1  g210(.A(G128), .B(G143), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(new_n218), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(KEYINPUT13), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n245), .A2(KEYINPUT13), .A3(G143), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(new_n218), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n400), .A2(new_n402), .B1(new_n218), .B2(new_n397), .ZN(new_n403));
  INV_X1    g217(.A(new_n396), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n395), .B1(new_n390), .B2(new_n388), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n385), .B1(new_n399), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n399), .A2(new_n406), .A3(new_n385), .ZN(new_n409));
  AOI21_X1  g223(.A(G902), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G478), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT15), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n410), .B(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n372), .A2(new_n382), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n224), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n346), .A2(G107), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n346), .A2(G107), .ZN(new_n418));
  OAI21_X1  g232(.A(G101), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT3), .B1(new_n346), .B2(G107), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n395), .A3(G104), .ZN(new_n422));
  INV_X1    g236(.A(G101), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n420), .A2(new_n422), .A3(new_n423), .A4(new_n416), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n257), .A2(new_n244), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n204), .A2(new_n207), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT1), .B1(new_n206), .B2(G146), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G128), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n244), .ZN(new_n431));
  INV_X1    g245(.A(new_n425), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n415), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n434), .B(KEYINPUT12), .Z(new_n435));
  INV_X1    g249(.A(KEYINPUT10), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n425), .A2(new_n436), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n433), .A2(new_n436), .B1(new_n248), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n212), .B1(new_n233), .B2(new_n239), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n420), .A2(new_n422), .A3(new_n416), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G101), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT4), .A3(new_n424), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(KEYINPUT4), .B2(new_n441), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n438), .B(new_n415), .C1(new_n439), .C2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G140), .ZN(new_n445));
  INV_X1    g259(.A(G227), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(G953), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n445), .B(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n435), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n433), .A2(new_n436), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n248), .A2(new_n437), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n439), .A2(new_n443), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n224), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n449), .B1(new_n456), .B2(new_n444), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G469), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n303), .ZN(new_n460));
  INV_X1    g274(.A(new_n444), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n448), .B1(new_n435), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n456), .A2(new_n449), .A3(new_n444), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G469), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n459), .A2(new_n303), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n460), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G210), .B1(G237), .B2(G902), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT79), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n261), .A2(G125), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n248), .A2(new_n326), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G224), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(G953), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n475), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n471), .A2(new_n477), .A3(new_n472), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(new_n191), .ZN(new_n481));
  INV_X1    g295(.A(G113), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n191), .B(new_n480), .C1(new_n193), .C2(new_n190), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n195), .A2(new_n196), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n432), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n199), .B2(new_n443), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n489));
  XNOR2_X1  g303(.A(G110), .B(G122), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n488), .A2(new_n491), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n490), .B(new_n487), .C1(new_n199), .C2(new_n443), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(KEYINPUT6), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n479), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n303), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n477), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n476), .A2(new_n478), .A3(new_n499), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n471), .A2(new_n498), .A3(new_n477), .A4(new_n472), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n485), .A2(new_n486), .A3(new_n425), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n490), .B(KEYINPUT8), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n195), .A2(KEYINPUT5), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n197), .B1(new_n504), .B2(new_n483), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n502), .B(new_n503), .C1(new_n505), .C2(new_n425), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n500), .A2(new_n501), .A3(new_n494), .A4(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n470), .B1(new_n497), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n496), .A2(new_n507), .A3(new_n303), .A4(new_n469), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G221), .B1(new_n383), .B2(G902), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n512), .B(KEYINPUT77), .Z(new_n513));
  OAI21_X1  g327(.A(G214), .B1(G237), .B2(G902), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n414), .A2(new_n468), .A3(new_n511), .A4(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n245), .A2(KEYINPUT23), .A3(G119), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n190), .A2(G128), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n190), .A2(G128), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n519), .B(new_n520), .C1(new_n521), .C2(KEYINPUT23), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n245), .A2(G119), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n520), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT24), .B(G110), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n522), .A2(G110), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n331), .A2(new_n528), .ZN(new_n529));
  OAI22_X1  g343(.A1(new_n525), .A2(new_n527), .B1(new_n522), .B2(G110), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n330), .A3(new_n350), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(KEYINPUT76), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT22), .B(G137), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n529), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n529), .B2(new_n531), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(G902), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT25), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n384), .B1(G234), .B2(new_n303), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n542), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n322), .A2(new_n518), .A3(new_n546), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT84), .B(G101), .Z(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(G3));
  NAND2_X1  g363(.A1(new_n294), .A2(new_n303), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G472), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n189), .B1(new_n286), .B2(new_n290), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n513), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n546), .A2(new_n468), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n495), .A2(new_n492), .ZN(new_n558));
  AOI21_X1  g372(.A(G902), .B1(new_n558), .B2(new_n479), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT85), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n469), .A4(new_n507), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n510), .A2(KEYINPUT85), .ZN(new_n562));
  INV_X1    g376(.A(new_n469), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n497), .B2(new_n508), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n514), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT86), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n410), .B2(G478), .ZN(new_n568));
  INV_X1    g382(.A(new_n409), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n303), .B1(new_n569), .B2(new_n407), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(KEYINPUT86), .A3(new_n411), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT33), .B1(new_n569), .B2(new_n407), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT33), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n408), .A2(new_n573), .A3(new_n409), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n411), .A2(G902), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n568), .A2(new_n571), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n357), .A2(new_n359), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n369), .A2(new_n371), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n566), .A2(new_n381), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n557), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G104), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(G6));
  INV_X1    g401(.A(new_n566), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT88), .ZN(new_n589));
  INV_X1    g403(.A(new_n413), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n372), .A2(new_n589), .A3(new_n382), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n372), .A2(new_n590), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT88), .B1(new_n592), .B2(new_n381), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n557), .A2(new_n588), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G107), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G9));
  NAND2_X1  g410(.A1(new_n529), .A2(new_n531), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n597), .A2(KEYINPUT89), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(KEYINPUT89), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OR3_X1    g414(.A1(new_n600), .A2(KEYINPUT36), .A3(new_n535), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n600), .B1(KEYINPUT36), .B2(new_n535), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n544), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n540), .B2(new_n541), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n517), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n552), .B1(new_n550), .B2(G472), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT37), .B(G110), .Z(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G12));
  NAND2_X1  g423(.A1(new_n468), .A2(new_n555), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT90), .B(G900), .Z(new_n612));
  AOI21_X1  g426(.A(new_n377), .B1(new_n379), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n372), .A2(new_n590), .A3(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n566), .A2(new_n604), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n322), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT91), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n322), .A2(KEYINPUT91), .A3(new_n611), .A4(new_n616), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT92), .B(G128), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G30));
  XNOR2_X1  g437(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n511), .B(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n372), .A2(new_n413), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(new_n604), .A3(new_n514), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n613), .B(KEYINPUT39), .Z(new_n628));
  NAND2_X1  g442(.A1(new_n611), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT95), .Z(new_n630));
  AOI211_X1 g444(.A(new_n625), .B(new_n627), .C1(new_n630), .C2(KEYINPUT40), .ZN(new_n631));
  INV_X1    g445(.A(new_n278), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n300), .A2(new_n273), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT94), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n303), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(G472), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n296), .A2(new_n636), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n630), .A2(KEYINPUT40), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n631), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G143), .ZN(G45));
  NOR3_X1   g454(.A1(new_n372), .A2(new_n577), .A3(new_n613), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT96), .B1(new_n642), .B2(new_n566), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT96), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n641), .A2(new_n565), .A3(new_n644), .A4(new_n514), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n604), .ZN(new_n647));
  AND4_X1   g461(.A1(new_n322), .A2(new_n646), .A3(new_n611), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n200), .ZN(G48));
  INV_X1    g463(.A(new_n460), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n459), .B1(new_n458), .B2(new_n303), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n650), .A2(new_n651), .A3(new_n513), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n566), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n582), .A2(new_n545), .A3(new_n381), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n322), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT41), .B(G113), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G15));
  AND2_X1   g472(.A1(new_n322), .A2(new_n654), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n593), .A2(new_n546), .A3(new_n591), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G116), .ZN(G18));
  NAND2_X1  g476(.A1(new_n372), .A2(new_n413), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n604), .A2(new_n663), .A3(new_n381), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G119), .ZN(G21));
  INV_X1    g480(.A(KEYINPUT97), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n274), .B1(new_n285), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n301), .A2(KEYINPUT97), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n278), .A2(KEYINPUT31), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT98), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n290), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n292), .A2(new_n673), .A3(new_n671), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n188), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n675), .A2(new_n551), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n626), .A2(new_n565), .A3(new_n514), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT99), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n626), .A2(new_n565), .A3(new_n679), .A4(new_n514), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n653), .A2(new_n381), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n676), .A2(new_n681), .A3(new_n682), .A4(new_n546), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G122), .ZN(G24));
  NAND3_X1  g498(.A1(new_n588), .A2(new_n652), .A3(new_n641), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n675), .A2(new_n551), .A3(new_n647), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n675), .A2(new_n551), .A3(KEYINPUT100), .A4(new_n647), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(new_n326), .ZN(G27));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n295), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n552), .A2(KEYINPUT102), .A3(KEYINPUT32), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n693), .A2(new_n694), .A3(new_n291), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT29), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n285), .B2(new_n273), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n266), .A2(new_n276), .A3(new_n277), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n697), .B1(new_n698), .B2(new_n273), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n319), .B1(new_n699), .B2(new_n315), .ZN(new_n700));
  INV_X1    g514(.A(new_n316), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n297), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n320), .A2(KEYINPUT75), .A3(G472), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n545), .B1(new_n695), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT101), .B1(new_n468), .B2(new_n555), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n511), .A2(new_n515), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n468), .A2(KEYINPUT101), .A3(new_n555), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n641), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n710), .ZN(new_n714));
  INV_X1    g528(.A(new_n709), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n714), .A2(new_n707), .A3(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n322), .A2(new_n716), .A3(new_n546), .A4(new_n641), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n706), .A2(new_n713), .B1(new_n717), .B2(new_n712), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n222), .ZN(G33));
  AOI21_X1  g533(.A(new_n545), .B1(new_n705), .B2(new_n296), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n615), .B(KEYINPUT103), .Z(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(KEYINPUT104), .A3(new_n716), .A4(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n322), .A2(new_n716), .A3(new_n546), .A4(new_n721), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G134), .ZN(G36));
  NAND2_X1  g541(.A1(new_n464), .A2(KEYINPUT45), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n462), .A2(new_n463), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n459), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n466), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n460), .B1(new_n732), .B2(KEYINPUT46), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n555), .A3(new_n628), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT105), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n735), .A2(new_n738), .A3(new_n555), .A4(new_n628), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n715), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  NAND2_X1  g555(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n581), .A2(new_n577), .ZN(new_n744));
  MUX2_X1   g558(.A(new_n742), .B(new_n743), .S(new_n744), .Z(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n554), .A3(new_n647), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT107), .B1(new_n746), .B2(new_n741), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n746), .A2(KEYINPUT107), .A3(new_n741), .ZN(new_n748));
  OAI221_X1 g562(.A(new_n740), .B1(new_n741), .B2(new_n746), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n735), .B(new_n555), .C1(KEYINPUT108), .C2(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n735), .A2(new_n555), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n709), .A2(new_n545), .A3(new_n641), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n322), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  NOR2_X1   g575(.A1(new_n648), .A2(new_n690), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n610), .A2(new_n647), .A3(new_n613), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n637), .A2(new_n681), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n621), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n762), .A2(new_n621), .A3(KEYINPUT52), .A4(new_n764), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n322), .B(new_n654), .C1(new_n660), .C2(new_n664), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n683), .A3(new_n656), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n718), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n582), .A2(new_n592), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n511), .A2(new_n774), .A3(new_n382), .A4(new_n514), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n557), .A2(new_n775), .B1(new_n605), .B2(new_n606), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n715), .A2(new_n663), .A3(new_n613), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n322), .A2(new_n611), .A3(new_n647), .A4(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n778), .A3(new_n547), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n711), .B1(new_n688), .B2(new_n689), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n772), .A2(new_n773), .A3(new_n726), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n780), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n776), .A2(new_n778), .A3(new_n547), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n726), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n706), .A2(new_n713), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n717), .A2(new_n712), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n770), .A2(new_n656), .A3(new_n683), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT109), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n769), .A2(new_n782), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT53), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n767), .A2(new_n794), .A3(new_n768), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n765), .A2(KEYINPUT110), .A3(new_n766), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n791), .A2(new_n782), .A3(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n793), .B(KEYINPUT54), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT111), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n795), .A2(new_n796), .ZN(new_n802));
  INV_X1    g616(.A(new_n799), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n805), .A3(KEYINPUT54), .A4(new_n793), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n772), .A2(KEYINPUT112), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n772), .A2(KEYINPUT112), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n781), .A2(KEYINPUT53), .A3(new_n726), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n802), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n792), .A2(new_n798), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n625), .B1(new_n815), .B2(KEYINPUT50), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n653), .A2(KEYINPUT113), .A3(new_n514), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT113), .B1(new_n653), .B2(new_n514), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT50), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n650), .A2(new_n651), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n513), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n755), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n823), .B1(new_n826), .B2(new_n715), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n745), .A2(new_n377), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n828), .A2(new_n546), .A3(new_n676), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n688), .A2(new_n689), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n652), .A2(new_n709), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n827), .A2(new_n829), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n835));
  INV_X1    g649(.A(new_n637), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n546), .A3(new_n377), .A4(new_n832), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n372), .A2(new_n577), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n837), .A2(new_n838), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n829), .A2(new_n819), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n840), .B2(new_n821), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n834), .A2(new_n835), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n835), .B1(new_n834), .B2(new_n841), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n833), .A2(new_n706), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT48), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n374), .B1(new_n837), .B2(new_n582), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n654), .B2(new_n829), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n842), .A2(new_n843), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n801), .A2(new_n806), .A3(new_n814), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n373), .A2(new_n269), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n824), .B(KEYINPUT49), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n546), .A2(new_n516), .A3(new_n744), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n836), .A2(new_n625), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n852), .A2(KEYINPUT116), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(G75));
  XNOR2_X1  g674(.A(new_n558), .B(new_n479), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT55), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT56), .B1(new_n863), .B2(KEYINPUT118), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n303), .B1(new_n811), .B2(new_n813), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n470), .ZN(new_n866));
  OAI221_X1 g680(.A(new_n864), .B1(KEYINPUT118), .B2(new_n863), .C1(new_n866), .C2(KEYINPUT117), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n269), .A2(G952), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT56), .B1(new_n865), .B2(G210), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n871), .B1(new_n872), .B2(new_n863), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n869), .A2(new_n873), .ZN(G51));
  AND3_X1   g688(.A1(new_n865), .A2(new_n728), .A3(new_n731), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n466), .B(KEYINPUT119), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT57), .Z(new_n877));
  INV_X1    g691(.A(new_n814), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n812), .B1(new_n811), .B2(new_n813), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n875), .B1(new_n880), .B2(new_n458), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT120), .B1(new_n881), .B2(new_n870), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n883));
  INV_X1    g697(.A(new_n458), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n811), .A2(new_n813), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n814), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n884), .B1(new_n887), .B2(new_n877), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n883), .B(new_n871), .C1(new_n888), .C2(new_n875), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n882), .A2(new_n889), .ZN(G54));
  OR2_X1    g704(.A1(new_n354), .A2(new_n367), .ZN(new_n891));
  AND2_X1   g705(.A1(KEYINPUT58), .A2(G475), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n865), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n891), .B1(new_n865), .B2(new_n892), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n893), .A2(new_n894), .A3(new_n870), .ZN(G60));
  XNOR2_X1  g709(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n411), .A2(new_n303), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n896), .B(new_n897), .Z(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n806), .A2(new_n814), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n802), .A2(new_n803), .B1(KEYINPUT53), .B2(new_n792), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n805), .B1(new_n901), .B2(KEYINPUT54), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n575), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n898), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n878), .B2(new_n879), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n905), .A2(KEYINPUT122), .A3(new_n871), .A4(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n801), .A2(new_n806), .A3(new_n814), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n575), .B1(new_n910), .B2(new_n899), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n871), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n908), .A2(new_n913), .ZN(G63));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT60), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n811), .B2(new_n813), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n601), .A2(new_n602), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n870), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n538), .B(KEYINPUT123), .Z(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n917), .B2(new_n918), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(KEYINPUT61), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n921), .B(new_n924), .ZN(G66));
  OAI21_X1  g739(.A(G953), .B1(new_n380), .B2(new_n474), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n776), .A2(new_n547), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n771), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n928), .B2(G953), .ZN(new_n929));
  INV_X1    g743(.A(new_n558), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(G898), .B2(new_n269), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n929), .B(new_n931), .ZN(G69));
  NAND2_X1  g746(.A1(new_n252), .A2(new_n253), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n309), .A2(new_n933), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(new_n361), .Z(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI211_X1 g750(.A(G900), .B(G953), .C1(new_n936), .C2(G227), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(G227), .B2(new_n936), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n737), .A2(new_n739), .B1(new_n680), .B2(new_n678), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n706), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n760), .A2(new_n788), .A3(new_n726), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n762), .A2(new_n621), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n749), .A2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n943), .A2(new_n749), .A3(KEYINPUT126), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n941), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(G953), .B1(new_n948), .B2(new_n936), .ZN(new_n949));
  AOI211_X1 g763(.A(new_n715), .B(new_n630), .C1(new_n582), .C2(new_n592), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n720), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n951), .A2(KEYINPUT125), .A3(new_n749), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT125), .B1(new_n951), .B2(new_n749), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n760), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n639), .A2(new_n943), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT62), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n935), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n938), .B1(new_n949), .B2(new_n957), .ZN(G72));
  NOR2_X1   g772(.A1(new_n698), .A2(new_n274), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n948), .A2(new_n928), .ZN(new_n960));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT63), .Z(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n959), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n964), .A2(new_n871), .ZN(new_n965));
  INV_X1    g779(.A(new_n901), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n273), .B1(new_n288), .B2(new_n266), .ZN(new_n967));
  NOR4_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n959), .A4(new_n963), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n928), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n954), .A2(new_n956), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n967), .B1(new_n971), .B2(new_n963), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n965), .A2(new_n969), .A3(KEYINPUT127), .A4(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n964), .A3(new_n871), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n968), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n973), .A2(new_n976), .ZN(G57));
endmodule


