

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U323 ( .A(n436), .B(n435), .Z(n546) );
  NAND2_X1 U324 ( .A1(n569), .A2(n294), .ZN(n291) );
  XOR2_X1 U325 ( .A(n320), .B(n422), .Z(n292) );
  XOR2_X1 U326 ( .A(n509), .B(KEYINPUT110), .Z(n293) );
  XOR2_X1 U327 ( .A(n411), .B(n410), .Z(n294) );
  INV_X1 U328 ( .A(KEYINPUT122), .ZN(n409) );
  NOR2_X1 U329 ( .A1(n545), .A2(n470), .ZN(n471) );
  XNOR2_X1 U330 ( .A(n409), .B(KEYINPUT54), .ZN(n410) );
  XOR2_X1 U331 ( .A(G120GAT), .B(G71GAT), .Z(n375) );
  NOR2_X1 U332 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U333 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U334 ( .A(n359), .B(n358), .ZN(n364) );
  NOR2_X1 U335 ( .A1(n475), .A2(n458), .ZN(n563) );
  INV_X1 U336 ( .A(n505), .ZN(n571) );
  NOR2_X1 U337 ( .A1(n519), .A2(n507), .ZN(n514) );
  INV_X1 U338 ( .A(n475), .ZN(n533) );
  XNOR2_X1 U339 ( .A(G183GAT), .B(KEYINPUT124), .ZN(n459) );
  XNOR2_X1 U340 ( .A(n460), .B(n459), .ZN(G1350GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n296) );
  XNOR2_X1 U342 ( .A(KEYINPUT78), .B(KEYINPUT14), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n316) );
  XOR2_X1 U344 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n298) );
  XNOR2_X1 U345 ( .A(KEYINPUT80), .B(KEYINPUT77), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U347 ( .A(KEYINPUT75), .B(G64GAT), .Z(n300) );
  XNOR2_X1 U348 ( .A(G1GAT), .B(G8GAT), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n314) );
  XOR2_X1 U351 ( .A(G22GAT), .B(G155GAT), .Z(n444) );
  XOR2_X1 U352 ( .A(n444), .B(G78GAT), .Z(n304) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G127GAT), .Z(n317) );
  XNOR2_X1 U354 ( .A(n317), .B(G211GAT), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n310) );
  XNOR2_X1 U356 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n305) );
  XNOR2_X1 U357 ( .A(n305), .B(KEYINPUT69), .ZN(n367) );
  INV_X1 U358 ( .A(KEYINPUT81), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n367), .B(n306), .ZN(n308) );
  NAND2_X1 U360 ( .A1(G231GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U362 ( .A(n310), .B(n309), .Z(n312) );
  XNOR2_X1 U363 ( .A(G183GAT), .B(G71GAT), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n579) );
  XOR2_X1 U367 ( .A(n317), .B(n375), .Z(n319) );
  NAND2_X1 U368 ( .A1(G227GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U370 ( .A(G134GAT), .B(KEYINPUT0), .Z(n422) );
  XOR2_X1 U371 ( .A(KEYINPUT83), .B(G190GAT), .Z(n322) );
  XNOR2_X1 U372 ( .A(G43GAT), .B(G99GAT), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U374 ( .A(G176GAT), .B(KEYINPUT82), .Z(n324) );
  XNOR2_X1 U375 ( .A(G169GAT), .B(G113GAT), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n292), .B(n327), .ZN(n328) );
  XOR2_X1 U379 ( .A(n328), .B(KEYINPUT84), .Z(n332) );
  XOR2_X1 U380 ( .A(G183GAT), .B(KEYINPUT19), .Z(n330) );
  XNOR2_X1 U381 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n338) );
  XNOR2_X1 U383 ( .A(n338), .B(KEYINPUT20), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n475) );
  XOR2_X1 U385 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n334) );
  NAND2_X1 U386 ( .A1(G226GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U388 ( .A(n335), .B(G92GAT), .Z(n340) );
  XOR2_X1 U389 ( .A(G64GAT), .B(KEYINPUT72), .Z(n337) );
  XNOR2_X1 U390 ( .A(G176GAT), .B(G204GAT), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n337), .B(n336), .ZN(n369) );
  XNOR2_X1 U392 ( .A(n338), .B(n369), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U394 ( .A(G36GAT), .B(G190GAT), .Z(n386) );
  XOR2_X1 U395 ( .A(n341), .B(n386), .Z(n346) );
  XOR2_X1 U396 ( .A(G169GAT), .B(G8GAT), .Z(n348) );
  XOR2_X1 U397 ( .A(KEYINPUT87), .B(G218GAT), .Z(n343) );
  XNOR2_X1 U398 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U400 ( .A(G197GAT), .B(n344), .ZN(n453) );
  XOR2_X1 U401 ( .A(n348), .B(n453), .Z(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n467) );
  XOR2_X1 U403 ( .A(G113GAT), .B(G1GAT), .Z(n428) );
  XOR2_X1 U404 ( .A(G22GAT), .B(G141GAT), .Z(n347) );
  XNOR2_X1 U405 ( .A(n428), .B(n347), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U407 ( .A(n350), .B(G50GAT), .Z(n359) );
  XOR2_X1 U408 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n352) );
  XNOR2_X1 U409 ( .A(G197GAT), .B(G15GAT), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n353), .B(G36GAT), .ZN(n357) );
  XOR2_X1 U412 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n355) );
  NAND2_X1 U413 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U415 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n361) );
  XNOR2_X1 U416 ( .A(G43GAT), .B(G29GAT), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U418 ( .A(KEYINPUT68), .B(n362), .Z(n399) );
  XNOR2_X1 U419 ( .A(n399), .B(KEYINPUT30), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n505) );
  XOR2_X1 U421 ( .A(KEYINPUT71), .B(G92GAT), .Z(n366) );
  XNOR2_X1 U422 ( .A(G99GAT), .B(G85GAT), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n395) );
  XOR2_X1 U424 ( .A(n367), .B(n395), .Z(n371) );
  XNOR2_X1 U425 ( .A(G106GAT), .B(G78GAT), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n368), .B(G148GAT), .ZN(n437) );
  XNOR2_X1 U427 ( .A(n437), .B(n369), .ZN(n370) );
  XOR2_X1 U428 ( .A(n371), .B(n370), .Z(n379) );
  XOR2_X1 U429 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n373) );
  XNOR2_X1 U430 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U432 ( .A(n375), .B(n374), .Z(n377) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n574) );
  XNOR2_X1 U436 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n574), .B(n380), .ZN(n559) );
  NAND2_X1 U438 ( .A1(n571), .A2(n559), .ZN(n381) );
  XOR2_X1 U439 ( .A(KEYINPUT46), .B(n381), .Z(n382) );
  NOR2_X1 U440 ( .A1(n579), .A2(n382), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n383), .B(KEYINPUT118), .ZN(n400) );
  XOR2_X1 U442 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n385) );
  XNOR2_X1 U443 ( .A(G134GAT), .B(G106GAT), .ZN(n384) );
  XOR2_X1 U444 ( .A(n385), .B(n384), .Z(n390) );
  XOR2_X1 U445 ( .A(KEYINPUT11), .B(n386), .Z(n388) );
  XOR2_X1 U446 ( .A(G50GAT), .B(G162GAT), .Z(n438) );
  XNOR2_X1 U447 ( .A(G218GAT), .B(n438), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n392) );
  NAND2_X1 U450 ( .A1(G232GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n394) );
  INV_X1 U452 ( .A(KEYINPUT10), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n395), .B(KEYINPUT73), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n399), .B(n398), .ZN(n461) );
  NAND2_X1 U457 ( .A1(n400), .A2(n461), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n401), .B(KEYINPUT47), .ZN(n407) );
  INV_X1 U459 ( .A(n579), .ZN(n492) );
  XNOR2_X1 U460 ( .A(KEYINPUT36), .B(KEYINPUT106), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n402), .B(n461), .ZN(n582) );
  NOR2_X1 U462 ( .A1(n492), .A2(n582), .ZN(n403) );
  XNOR2_X1 U463 ( .A(KEYINPUT45), .B(n403), .ZN(n404) );
  NAND2_X1 U464 ( .A1(n404), .A2(n574), .ZN(n405) );
  NOR2_X1 U465 ( .A1(n405), .A2(n571), .ZN(n406) );
  NOR2_X1 U466 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n408), .B(KEYINPUT48), .ZN(n548) );
  NOR2_X1 U468 ( .A1(n467), .A2(n548), .ZN(n411) );
  XOR2_X1 U469 ( .A(KEYINPUT1), .B(KEYINPUT95), .Z(n413) );
  XNOR2_X1 U470 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n436) );
  XOR2_X1 U472 ( .A(KEYINPUT91), .B(KEYINPUT96), .Z(n415) );
  XNOR2_X1 U473 ( .A(G120GAT), .B(KEYINPUT6), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U475 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n417) );
  XNOR2_X1 U476 ( .A(G57GAT), .B(KEYINPUT94), .ZN(n416) );
  XNOR2_X1 U477 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U478 ( .A(n419), .B(n418), .Z(n434) );
  XOR2_X1 U479 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n421) );
  XNOR2_X1 U480 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n448) );
  XOR2_X1 U482 ( .A(n448), .B(n422), .Z(n424) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n432) );
  XOR2_X1 U485 ( .A(G85GAT), .B(G148GAT), .Z(n426) );
  XNOR2_X1 U486 ( .A(G127GAT), .B(G162GAT), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U488 ( .A(n427), .B(G155GAT), .Z(n430) );
  XNOR2_X1 U489 ( .A(G29GAT), .B(n428), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n435) );
  INV_X1 U493 ( .A(n546), .ZN(n569) );
  XOR2_X1 U494 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U495 ( .A1(G228GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n452) );
  XOR2_X1 U497 ( .A(G204GAT), .B(KEYINPUT22), .Z(n442) );
  XNOR2_X1 U498 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U500 ( .A(n443), .B(KEYINPUT89), .Z(n446) );
  XNOR2_X1 U501 ( .A(n444), .B(KEYINPUT24), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U503 ( .A(n447), .B(KEYINPUT23), .Z(n450) );
  XNOR2_X1 U504 ( .A(n448), .B(KEYINPUT90), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n472) );
  AND2_X1 U508 ( .A1(n569), .A2(n472), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n294), .A2(n455), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n456), .B(KEYINPUT123), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n457), .B(KEYINPUT55), .ZN(n458) );
  NAND2_X1 U512 ( .A1(n579), .A2(n563), .ZN(n460) );
  XNOR2_X1 U513 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n482) );
  NAND2_X1 U514 ( .A1(n571), .A2(n574), .ZN(n495) );
  INV_X1 U515 ( .A(n461), .ZN(n564) );
  NOR2_X1 U516 ( .A1(n564), .A2(n492), .ZN(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT16), .B(n462), .ZN(n479) );
  NOR2_X1 U518 ( .A1(n533), .A2(n472), .ZN(n464) );
  XNOR2_X1 U519 ( .A(KEYINPUT101), .B(KEYINPUT26), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U521 ( .A(KEYINPUT100), .B(n465), .ZN(n570) );
  XOR2_X1 U522 ( .A(n467), .B(KEYINPUT99), .Z(n466) );
  XNOR2_X1 U523 ( .A(KEYINPUT27), .B(n466), .ZN(n474) );
  NOR2_X1 U524 ( .A1(n570), .A2(n474), .ZN(n545) );
  INV_X1 U525 ( .A(n467), .ZN(n523) );
  NAND2_X1 U526 ( .A1(n533), .A2(n523), .ZN(n468) );
  NAND2_X1 U527 ( .A1(n472), .A2(n468), .ZN(n469) );
  XNOR2_X1 U528 ( .A(KEYINPUT25), .B(n469), .ZN(n470) );
  NOR2_X1 U529 ( .A1(n546), .A2(n471), .ZN(n477) );
  XNOR2_X1 U530 ( .A(KEYINPUT28), .B(n472), .ZN(n488) );
  NAND2_X1 U531 ( .A1(n546), .A2(n488), .ZN(n473) );
  NOR2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n534) );
  AND2_X1 U533 ( .A1(n534), .A2(n475), .ZN(n476) );
  XOR2_X1 U534 ( .A(KEYINPUT102), .B(n478), .Z(n491) );
  NAND2_X1 U535 ( .A1(n479), .A2(n491), .ZN(n480) );
  XOR2_X1 U536 ( .A(KEYINPUT103), .B(n480), .Z(n507) );
  NOR2_X1 U537 ( .A1(n495), .A2(n507), .ZN(n489) );
  NAND2_X1 U538 ( .A1(n546), .A2(n489), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(G1324GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n484) );
  NAND2_X1 U541 ( .A1(n489), .A2(n523), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n485), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U545 ( .A1(n489), .A2(n533), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  INV_X1 U547 ( .A(n488), .ZN(n528) );
  NAND2_X1 U548 ( .A1(n528), .A2(n489), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U550 ( .A1(n492), .A2(n491), .ZN(n493) );
  NOR2_X1 U551 ( .A1(n493), .A2(n582), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n494), .B(KEYINPUT37), .ZN(n518) );
  NOR2_X1 U553 ( .A1(n495), .A2(n518), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n496), .B(KEYINPUT38), .ZN(n503) );
  NAND2_X1 U555 ( .A1(n546), .A2(n503), .ZN(n498) );
  XOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .Z(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n503), .A2(n523), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n501) );
  NAND2_X1 U561 ( .A1(n503), .A2(n533), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n503), .A2(n528), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n504), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U566 ( .A1(n505), .A2(n559), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n506), .B(KEYINPUT108), .ZN(n519) );
  NAND2_X1 U568 ( .A1(n514), .A2(n546), .ZN(n508) );
  XNOR2_X1 U569 ( .A(n508), .B(KEYINPUT109), .ZN(n509) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n293), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n523), .A2(n514), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT111), .Z(n513) );
  NAND2_X1 U575 ( .A1(n514), .A2(n533), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U578 ( .A1(n514), .A2(n528), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(n517), .ZN(G1335GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n521) );
  NOR2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n529), .A2(n546), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  XOR2_X1 U586 ( .A(G92GAT), .B(KEYINPUT115), .Z(n525) );
  NAND2_X1 U587 ( .A1(n529), .A2(n523), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n533), .A2(n529), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(KEYINPUT116), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(n527), .ZN(G1338GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT117), .B(KEYINPUT44), .Z(n531) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  XOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT119), .Z(n537) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U598 ( .A1(n548), .A2(n535), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n542), .A2(n571), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U602 ( .A1(n542), .A2(n559), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NAND2_X1 U604 ( .A1(n579), .A2(n542), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n540), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U608 ( .A1(n542), .A2(n564), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n571), .A2(n555), .ZN(n549) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n553) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n551) );
  NAND2_X1 U616 ( .A1(n555), .A2(n559), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n579), .A2(n555), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U621 ( .A(G162GAT), .B(KEYINPUT121), .Z(n557) );
  NAND2_X1 U622 ( .A1(n555), .A2(n564), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n563), .A2(n571), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n563), .A2(n559), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(n562), .ZN(G1349GAT) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1351GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n573) );
  NOR2_X1 U636 ( .A1(n291), .A2(n570), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n578), .A2(n571), .ZN(n572) );
  XOR2_X1 U638 ( .A(n573), .B(n572), .Z(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n576) );
  INV_X1 U640 ( .A(n578), .ZN(n581) );
  OR2_X1 U641 ( .A1(n581), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

