//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT31), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n191), .A3(G116), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n196), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n192), .A3(new_n194), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT0), .B(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(G137), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n209), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n211), .A2(G137), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n213), .A2(G134), .ZN(new_n222));
  OAI21_X1  g036(.A(G131), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT68), .B1(new_n217), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n225));
  AOI21_X1  g039(.A(G128), .B1(new_n202), .B2(new_n204), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n227), .A2(new_n201), .A3(G143), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n225), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n201), .A2(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n231), .B(KEYINPUT66), .C1(new_n207), .C2(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n207), .A2(new_n227), .A3(G128), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n224), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n217), .A2(new_n223), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT68), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n220), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT69), .B1(new_n239), .B2(KEYINPUT30), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n209), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n219), .A2(new_n217), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n206), .B(KEYINPUT64), .C1(new_n207), .C2(new_n208), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT65), .ZN(new_n246));
  INV_X1    g060(.A(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n203), .A2(G146), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(new_n230), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT66), .B1(new_n249), .B2(new_n231), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n226), .A2(new_n225), .A3(new_n228), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n234), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n237), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n242), .A2(new_n243), .A3(new_n254), .A4(new_n244), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n246), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT30), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n240), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n239), .A2(KEYINPUT69), .A3(KEYINPUT30), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n200), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n224), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n252), .A2(new_n238), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n220), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n200), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G237), .ZN(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G210), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT27), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n187), .B1(new_n261), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n272), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n263), .A2(KEYINPUT30), .A3(new_n264), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n258), .B2(new_n240), .ZN(new_n278));
  OAI211_X1 g092(.A(KEYINPUT31), .B(new_n274), .C1(new_n278), .C2(new_n200), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n265), .A2(KEYINPUT28), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT28), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n239), .A2(new_n281), .A3(new_n200), .ZN(new_n282));
  INV_X1    g096(.A(new_n200), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n280), .A2(new_n282), .B1(new_n283), .B2(new_n256), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT70), .B1(new_n284), .B2(new_n271), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n282), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n256), .A2(new_n283), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  INV_X1    g103(.A(new_n271), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n273), .A2(new_n279), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(G472), .A2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT71), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n285), .ZN(new_n296));
  AOI22_X1  g110(.A1(KEYINPUT65), .A2(new_n245), .B1(new_n252), .B2(new_n237), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT30), .B1(new_n297), .B2(new_n255), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n275), .A2(new_n276), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n260), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n283), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT31), .B1(new_n301), .B2(new_n274), .ZN(new_n302));
  AOI211_X1 g116(.A(new_n187), .B(new_n272), .C1(new_n300), .C2(new_n283), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n296), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n293), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT32), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n295), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n273), .A2(new_n279), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n294), .B1(new_n309), .B2(new_n296), .ZN(new_n310));
  OR2_X1    g124(.A1(new_n239), .A2(new_n200), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n286), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n271), .A2(KEYINPUT29), .ZN(new_n314));
  AOI21_X1  g128(.A(G902), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n284), .A2(new_n290), .ZN(new_n316));
  INV_X1    g130(.A(new_n265), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n300), .B2(new_n283), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n318), .B2(new_n290), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n315), .B1(new_n319), .B2(KEYINPUT29), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n310), .A2(KEYINPUT32), .B1(new_n320), .B2(G472), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n308), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT75), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT22), .B(G137), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G125), .B(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT16), .ZN(new_n329));
  INV_X1    g143(.A(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G125), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(KEYINPUT16), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n201), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n329), .B(G146), .C1(KEYINPUT16), .C2(new_n331), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT67), .B(G119), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(G128), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n188), .A2(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT23), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n337), .A2(G128), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G110), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT24), .B(G110), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n337), .A2(KEYINPUT73), .A3(G128), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n339), .A2(KEYINPUT73), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n335), .B(new_n343), .C1(new_n344), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n328), .A2(new_n201), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n334), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT73), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n341), .B(new_n352), .C1(new_n188), .C2(G128), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n344), .A3(new_n345), .ZN(new_n354));
  INV_X1    g168(.A(G110), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n338), .A2(new_n355), .A3(new_n340), .A4(new_n341), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n351), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n349), .B1(new_n357), .B2(KEYINPUT74), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(KEYINPUT74), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n327), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n357), .A2(KEYINPUT74), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(new_n359), .A3(new_n349), .A4(new_n326), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  AOI21_X1  g179(.A(G902), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n364), .A2(new_n365), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT72), .B(G217), .Z(new_n370));
  INV_X1    g184(.A(G902), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n370), .B1(G234), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n368), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n361), .A2(new_n363), .A3(new_n373), .A4(new_n366), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n369), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n361), .A2(new_n363), .ZN(new_n376));
  INV_X1    g190(.A(new_n372), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n371), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(KEYINPUT77), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT9), .B(G234), .ZN(new_n383));
  OAI21_X1  g197(.A(G221), .B1(new_n383), .B2(G902), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT78), .ZN(new_n385));
  XNOR2_X1  g199(.A(G110), .B(G140), .ZN(new_n386));
  INV_X1    g200(.A(G227), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(G953), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n386), .B(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT12), .B1(new_n243), .B2(KEYINPUT81), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n394));
  INV_X1    g208(.A(G107), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(G104), .ZN(new_n396));
  INV_X1    g210(.A(G101), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(G107), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n396), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n392), .A2(G107), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n395), .A2(G104), .ZN(new_n401));
  OAI21_X1  g215(.A(G101), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n226), .A2(new_n228), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n403), .B1(new_n234), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT80), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n399), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n406), .B1(new_n399), .B2(new_n402), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n207), .A2(new_n227), .A3(G128), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n229), .B2(new_n232), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n405), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n243), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n391), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n404), .A2(new_n234), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n399), .A3(new_n402), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n403), .A2(KEYINPUT80), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n399), .A2(new_n402), .A3(new_n406), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n416), .B1(new_n419), .B2(new_n252), .ZN(new_n420));
  INV_X1    g234(.A(new_n391), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n243), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n393), .A2(new_n396), .A3(new_n398), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n424), .A2(new_n425), .A3(G101), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(new_n209), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT79), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n399), .A2(KEYINPUT4), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n424), .A2(G101), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AND4_X1   g245(.A1(new_n428), .A2(new_n430), .A3(KEYINPUT4), .A4(new_n399), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n427), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT10), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n419), .B2(new_n252), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n416), .A2(KEYINPUT10), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n433), .B(new_n413), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n390), .B1(new_n423), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT10), .B1(new_n409), .B2(new_n411), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(KEYINPUT10), .B2(new_n416), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n413), .B1(new_n440), .B2(new_n433), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT82), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n390), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n437), .A2(KEYINPUT82), .A3(new_n390), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n438), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G469), .B1(new_n446), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(G469), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n443), .A2(KEYINPUT84), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n437), .A2(new_n450), .A3(new_n390), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n423), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n243), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n390), .B1(new_n454), .B2(new_n437), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(G902), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n447), .A2(KEYINPUT83), .B1(new_n448), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT83), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n459), .B(G469), .C1(new_n446), .C2(G902), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n385), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G475), .ZN(new_n462));
  INV_X1    g276(.A(new_n335), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n266), .A2(new_n267), .A3(G214), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n203), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n266), .A2(new_n267), .A3(G143), .A4(G214), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(new_n215), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT17), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI211_X1 g284(.A(new_n469), .B(new_n215), .C1(new_n465), .C2(new_n466), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n471), .A2(KEYINPUT96), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(KEYINPUT96), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n463), .A2(new_n470), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT90), .ZN(new_n475));
  INV_X1    g289(.A(G125), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(G140), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n330), .A2(G125), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(G140), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n331), .A2(new_n480), .A3(KEYINPUT90), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n350), .B1(new_n482), .B2(new_n201), .ZN(new_n483));
  INV_X1    g297(.A(new_n467), .ZN(new_n484));
  AND4_X1   g298(.A1(KEYINPUT91), .A2(new_n484), .A3(KEYINPUT18), .A4(G131), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n484), .A2(KEYINPUT91), .B1(KEYINPUT18), .B2(G131), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(G113), .B(G122), .Z(new_n488));
  XOR2_X1   g302(.A(KEYINPUT94), .B(G104), .Z(new_n489));
  XOR2_X1   g303(.A(new_n488), .B(new_n489), .Z(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT95), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n474), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n474), .A2(new_n487), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n492), .B1(new_n493), .B2(new_n490), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n462), .B1(new_n494), .B2(new_n371), .ZN(new_n495));
  INV_X1    g309(.A(new_n492), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT19), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n479), .B2(new_n481), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n328), .A2(KEYINPUT19), .ZN(new_n500));
  OAI211_X1 g314(.A(KEYINPUT92), .B(new_n201), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n334), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n331), .A2(new_n480), .A3(KEYINPUT90), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT90), .B1(new_n331), .B2(new_n480), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT19), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n500), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT92), .B1(new_n507), .B2(new_n201), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n497), .B1(new_n502), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n468), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n500), .B1(new_n482), .B2(KEYINPUT19), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(G146), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n513), .A2(KEYINPUT93), .A3(new_n334), .A4(new_n501), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n509), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n487), .ZN(new_n516));
  INV_X1    g330(.A(new_n490), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n496), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(G475), .A2(G902), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT20), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT20), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n490), .B1(new_n515), .B2(new_n487), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(new_n519), .C1(new_n523), .C2(new_n496), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n495), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G478), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(KEYINPUT15), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n370), .A2(G953), .A3(new_n383), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n193), .A2(KEYINPUT14), .A3(G122), .ZN(new_n531));
  INV_X1    g345(.A(G122), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G116), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n193), .A2(G122), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(G107), .B(new_n531), .C1(new_n535), .C2(KEYINPUT14), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n203), .A2(G128), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n247), .A2(G143), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(G134), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n211), .B1(new_n537), .B2(new_n538), .ZN(new_n541));
  OAI221_X1 g355(.A(new_n536), .B1(G107), .B2(new_n535), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT13), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n544), .A2(new_n203), .A3(G128), .ZN(new_n545));
  OAI211_X1 g359(.A(G134), .B(new_n545), .C1(new_n539), .C2(new_n544), .ZN(new_n546));
  INV_X1    g360(.A(new_n540), .ZN(new_n547));
  INV_X1    g361(.A(new_n535), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(new_n395), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n535), .A2(G107), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n546), .B(new_n547), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n542), .A2(new_n543), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n543), .B1(new_n542), .B2(new_n551), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n530), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n542), .A2(new_n551), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT97), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(new_n529), .A3(new_n552), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n528), .B1(new_n559), .B2(new_n371), .ZN(new_n560));
  AOI211_X1 g374(.A(G902), .B(new_n527), .C1(new_n555), .C2(new_n558), .ZN(new_n561));
  NAND2_X1  g375(.A1(G234), .A2(G237), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n562), .A2(G952), .A3(new_n267), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT21), .B(G898), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT98), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n562), .A2(G902), .A3(G953), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n560), .A2(new_n561), .A3(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n525), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G214), .B1(G237), .B2(G902), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(G110), .B(G122), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT86), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n426), .B1(new_n197), .B2(new_n199), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT85), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n576), .B(new_n577), .C1(new_n431), .C2(new_n432), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n192), .A2(KEYINPUT5), .A3(new_n194), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n579), .B(G113), .C1(KEYINPUT5), .C2(new_n192), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n580), .B(new_n199), .C1(new_n408), .C2(new_n407), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n430), .A2(KEYINPUT4), .A3(new_n399), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT79), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n429), .A2(new_n428), .A3(new_n430), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n577), .B1(new_n586), .B2(new_n576), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n575), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n576), .B1(new_n431), .B2(new_n432), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT85), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n573), .B(KEYINPUT86), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n578), .A4(new_n581), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n588), .A2(KEYINPUT6), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n209), .A2(G125), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT87), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT87), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n209), .A2(new_n596), .A3(G125), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n411), .A2(new_n476), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n267), .A2(G224), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g416(.A(KEYINPUT6), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n603), .B(new_n575), .C1(new_n582), .C2(new_n587), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n593), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n601), .A2(KEYINPUT7), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n599), .B2(new_n594), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT8), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n591), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n575), .A2(KEYINPUT8), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n192), .A2(KEYINPUT5), .A3(new_n194), .ZN(new_n612));
  OAI21_X1  g426(.A(G113), .B1(new_n192), .B2(KEYINPUT5), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n199), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n403), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n611), .B1(new_n581), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n599), .A2(new_n595), .A3(new_n597), .A4(new_n606), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT88), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT88), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n598), .A2(new_n619), .A3(new_n599), .A4(new_n606), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n607), .B(new_n616), .C1(new_n618), .C2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(G902), .B1(new_n621), .B2(new_n592), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n605), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(G210), .B1(G237), .B2(G902), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT89), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n625), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n605), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n572), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n570), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n322), .A2(new_n382), .A3(new_n461), .A4(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G101), .ZN(G3));
  OAI21_X1  g446(.A(G472), .B1(new_n292), .B2(G902), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n295), .A2(new_n633), .A3(new_n306), .A4(new_n382), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n443), .A2(new_n442), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n445), .A3(new_n454), .ZN(new_n636));
  INV_X1    g450(.A(new_n438), .ZN(new_n637));
  AOI21_X1  g451(.A(G902), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT83), .B1(new_n638), .B2(new_n448), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n457), .A2(new_n448), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n460), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n385), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n521), .A2(new_n524), .ZN(new_n645));
  INV_X1    g459(.A(new_n495), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n559), .B(KEYINPUT33), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n526), .A2(G902), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n559), .A2(new_n371), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n648), .A2(new_n649), .B1(new_n526), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n568), .ZN(new_n654));
  INV_X1    g468(.A(new_n628), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n627), .B1(new_n605), .B2(new_n622), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n571), .B(new_n654), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n644), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  NOR2_X1   g475(.A1(new_n560), .A2(new_n561), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n657), .A2(new_n647), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n644), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NAND4_X1  g480(.A1(new_n570), .A2(new_n641), .A3(new_n642), .A4(new_n629), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n362), .A2(new_n359), .A3(new_n349), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT36), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n326), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT99), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n668), .A2(new_n671), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n380), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n375), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n295), .A2(new_n633), .A3(new_n306), .A4(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n667), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT37), .B(G110), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  AND2_X1   g493(.A1(new_n375), .A2(new_n674), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n681));
  INV_X1    g495(.A(new_n567), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n681), .B1(new_n682), .B2(G900), .ZN(new_n683));
  INV_X1    g497(.A(new_n563), .ZN(new_n684));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n567), .A2(KEYINPUT100), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n680), .A2(new_n647), .A3(new_n662), .A4(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n322), .A2(new_n461), .A3(new_n629), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT101), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n643), .B1(new_n308), .B2(new_n321), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n629), .A4(new_n689), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  XNOR2_X1  g510(.A(new_n687), .B(KEYINPUT39), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n461), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT103), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT40), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n662), .A2(new_n572), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n647), .A2(new_n680), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT102), .ZN(new_n704));
  INV_X1    g518(.A(new_n318), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n271), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n317), .A2(new_n271), .ZN(new_n707));
  AOI21_X1  g521(.A(G902), .B1(new_n707), .B2(new_n311), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n310), .A2(KEYINPUT32), .B1(new_n709), .B2(G472), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n308), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n626), .A2(new_n628), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(KEYINPUT38), .Z(new_n714));
  NOR3_X1   g528(.A1(new_n704), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n701), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n699), .A2(new_n700), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n203), .ZN(G45));
  NOR3_X1   g533(.A1(new_n653), .A2(new_n680), .A3(new_n688), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n322), .A2(new_n461), .A3(new_n629), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G146), .ZN(G48));
  NOR2_X1   g536(.A1(new_n448), .A2(KEYINPUT104), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n457), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n443), .A2(KEYINPUT84), .B1(new_n422), .B2(new_n414), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n455), .B1(new_n726), .B2(new_n451), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n723), .B1(new_n727), .B2(G902), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(new_n728), .A3(new_n642), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n322), .A2(new_n382), .A3(new_n658), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(KEYINPUT41), .B(G113), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G15));
  INV_X1    g547(.A(new_n382), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n308), .B2(new_n321), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n663), .A3(new_n730), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  NAND2_X1  g551(.A1(new_n713), .A2(new_n571), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n675), .A2(new_n525), .A3(new_n569), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n738), .A2(new_n739), .A3(new_n729), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n322), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  NAND3_X1  g556(.A1(new_n713), .A2(new_n647), .A3(new_n702), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n725), .A2(new_n728), .A3(new_n642), .A4(new_n654), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n312), .A2(KEYINPUT105), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n290), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n312), .A2(KEYINPUT105), .ZN(new_n748));
  OAI22_X1  g562(.A1(new_n302), .A2(new_n303), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n293), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n633), .A2(new_n382), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  NOR2_X1   g567(.A1(new_n738), .A2(new_n729), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n633), .A2(new_n750), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n653), .A2(new_n688), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .A4(new_n675), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  NAND3_X1  g572(.A1(new_n626), .A2(new_n571), .A3(new_n628), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n385), .B1(new_n640), .B2(new_n447), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n756), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n310), .A2(KEYINPUT32), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n320), .A2(G472), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n307), .B1(new_n292), .B2(new_n294), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n382), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT42), .B1(new_n762), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n760), .A2(new_n761), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n735), .A2(new_n769), .A3(new_n756), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n215), .ZN(G33));
  NOR3_X1   g587(.A1(new_n647), .A2(new_n662), .A3(new_n688), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n735), .A2(new_n774), .A3(new_n770), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  OAI21_X1  g590(.A(G469), .B1(new_n446), .B2(KEYINPUT45), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(KEYINPUT45), .B2(new_n446), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT106), .ZN(new_n779));
  NAND2_X1  g593(.A1(G469), .A2(G902), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT46), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT107), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n779), .A2(new_n784), .A3(KEYINPUT46), .A4(new_n780), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n781), .A2(new_n782), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n783), .A2(new_n640), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(new_n642), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n295), .A2(new_n633), .A3(new_n306), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n680), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n652), .A2(new_n525), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n791), .B(KEYINPUT43), .Z(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT44), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n759), .B(KEYINPUT108), .Z(new_n795));
  NAND4_X1  g609(.A1(new_n788), .A2(new_n697), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  NAND3_X1  g611(.A1(new_n756), .A2(new_n734), .A3(new_n760), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n322), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n787), .A2(new_n642), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT47), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n800), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n330), .ZN(G42));
  NAND2_X1  g620(.A1(new_n725), .A2(new_n728), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(KEYINPUT49), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(KEYINPUT49), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n382), .A2(new_n642), .A3(new_n571), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n791), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n712), .A3(new_n714), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n721), .A2(new_n757), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n743), .A2(new_n675), .A3(new_n688), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n711), .A2(new_n815), .A3(new_n761), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n695), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT52), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n813), .B1(new_n694), .B2(new_n691), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n816), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n650), .A2(new_n527), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n559), .A2(new_n371), .A3(new_n528), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(KEYINPUT110), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n560), .B2(new_n561), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n629), .A2(new_n525), .A3(new_n654), .A4(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n634), .A2(new_n828), .A3(new_n643), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT111), .B1(new_n829), .B2(new_n677), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n789), .A2(new_n630), .A3(new_n461), .A4(new_n675), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n525), .A2(new_n827), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n657), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n789), .A2(new_n382), .A3(new_n461), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n322), .A2(new_n740), .B1(new_n745), .B2(new_n751), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n838), .A2(new_n631), .A3(new_n731), .ZN(new_n839));
  INV_X1    g653(.A(new_n657), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(KEYINPUT109), .A3(new_n647), .A4(new_n652), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT109), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n653), .B2(new_n657), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n644), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n844), .A2(new_n736), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n837), .A2(new_n839), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n768), .A2(new_n771), .A3(new_n775), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n760), .A2(new_n675), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n525), .A2(new_n687), .A3(new_n824), .A4(new_n826), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT112), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n692), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n755), .A2(new_n756), .A3(new_n761), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n818), .A2(new_n821), .A3(new_n846), .A4(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n838), .A2(new_n731), .A3(new_n631), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n844), .A2(new_n736), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n854), .A2(new_n860), .A3(new_n837), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(KEYINPUT53), .A3(new_n821), .A4(new_n818), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  XNOR2_X1  g678(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n730), .A2(new_n572), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(KEYINPUT114), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(KEYINPUT114), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n714), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT115), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n792), .A2(new_n563), .A3(new_n751), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n870), .A2(new_n875), .A3(new_n714), .A4(new_n871), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT50), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT116), .B1(new_n730), .B2(new_n760), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n729), .A2(new_n759), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n881), .A3(new_n684), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n792), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n755), .A2(new_n675), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT117), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n882), .A2(new_n382), .A3(new_n712), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n887), .A2(new_n647), .A3(new_n652), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n878), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n725), .A2(new_n728), .A3(new_n385), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n801), .A2(new_n804), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n874), .A2(new_n795), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n889), .B(KEYINPUT51), .C1(new_n891), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n267), .A2(G952), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n874), .B2(new_n754), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n883), .A2(new_n767), .ZN(new_n899));
  XOR2_X1   g713(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n900));
  OAI221_X1 g714(.A(new_n898), .B1(new_n653), .B2(new_n887), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n868), .A2(new_n895), .A3(new_n896), .A4(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(G952), .A2(G953), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n812), .B1(new_n903), .B2(new_n904), .ZN(G75));
  NAND2_X1  g719(.A1(new_n593), .A2(new_n604), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n602), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT55), .Z(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n863), .B2(G902), .ZN(new_n913));
  AOI211_X1 g727(.A(KEYINPUT119), .B(new_n371), .C1(new_n857), .C2(new_n862), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n915), .B2(new_n625), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n267), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n371), .B1(new_n857), .B2(new_n862), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(new_n625), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n920), .B2(new_n909), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT120), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n625), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n910), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n917), .B1(new_n924), .B2(new_n908), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n913), .A2(new_n914), .A3(new_n627), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(new_n911), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n922), .A2(new_n928), .ZN(G51));
  XOR2_X1   g743(.A(new_n780), .B(KEYINPUT57), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n863), .A2(new_n866), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n932), .B2(new_n867), .ZN(new_n933));
  INV_X1    g747(.A(new_n727), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n779), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n915), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n917), .B1(new_n935), .B2(new_n937), .ZN(G54));
  AND2_X1   g752(.A1(KEYINPUT58), .A2(G475), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n915), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n518), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n915), .B(new_n939), .C1(new_n496), .C2(new_n523), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n941), .A2(new_n918), .A3(new_n942), .ZN(G60));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n944));
  INV_X1    g758(.A(new_n648), .ZN(new_n945));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT59), .Z(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n857), .A2(new_n862), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n865), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n949), .B1(new_n951), .B2(new_n931), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n944), .B1(new_n952), .B2(new_n917), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n948), .B1(new_n932), .B2(new_n867), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(KEYINPUT121), .A3(new_n918), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n945), .B1(new_n868), .B2(new_n947), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(G63));
  XNOR2_X1  g771(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n958));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n950), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n672), .A2(new_n673), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n917), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n376), .B(KEYINPUT123), .Z(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n963), .B(KEYINPUT61), .C1(new_n961), .C2(new_n964), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(G66));
  AOI21_X1  g783(.A(new_n267), .B1(new_n565), .B2(G224), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT124), .Z(new_n971));
  INV_X1    g785(.A(new_n846), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n267), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT125), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n906), .B1(G898), .B2(new_n267), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G69));
  XNOR2_X1  g790(.A(new_n300), .B(new_n507), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT126), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n759), .B1(new_n653), .B2(new_n832), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n699), .A2(new_n735), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n796), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n805), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n819), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n718), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT62), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n978), .B1(new_n986), .B2(new_n267), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n977), .B1(new_n685), .B2(new_n267), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n767), .A2(new_n743), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n788), .A2(new_n697), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n983), .A2(new_n847), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n796), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n993), .A2(new_n805), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n989), .B1(new_n994), .B2(new_n267), .ZN(new_n995));
  OR3_X1    g809(.A1(new_n987), .A2(new_n988), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n988), .B1(new_n987), .B2(new_n995), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(G72));
  NOR3_X1   g812(.A1(new_n993), .A2(new_n805), .A3(new_n972), .ZN(new_n999));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n290), .B(new_n318), .C1(new_n999), .C2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n318), .B2(new_n290), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n863), .A2(new_n706), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1003), .A2(new_n1005), .A3(new_n918), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1001), .B1(new_n986), .B2(new_n972), .ZN(new_n1007));
  INV_X1    g821(.A(new_n706), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(KEYINPUT127), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT127), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1007), .A2(new_n1011), .A3(new_n1008), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1006), .B1(new_n1010), .B2(new_n1012), .ZN(G57));
endmodule


