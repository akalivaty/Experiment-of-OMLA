//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  XOR2_X1   g0012(.A(KEYINPUT65), .B(G244), .Z(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G107), .A2(G264), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n212), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  NAND3_X1  g0024(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n212), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n226), .B1(new_n229), .B2(KEYINPUT0), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n230), .B1(KEYINPUT0), .B2(new_n229), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n223), .B(new_n232), .C1(KEYINPUT1), .C2(new_n221), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n245), .B(new_n251), .ZN(G351));
  OAI21_X1  g0052(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  OAI211_X1 g0056(.A(G1), .B(G13), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n257), .A3(G274), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n253), .ZN(new_n259));
  INV_X1    g0059(.A(G226), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G222), .A2(G1698), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G223), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n257), .B1(new_n270), .B2(new_n214), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n261), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT70), .B(G200), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(G190), .B2(new_n272), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G1), .A2(G13), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n209), .A2(G20), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G50), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G150), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n210), .A2(G33), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(G20), .B2(new_n203), .ZN(new_n289));
  INV_X1    g0089(.A(new_n280), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n283), .B1(G50), .B2(new_n276), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT9), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n292), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n275), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(G179), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n272), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n291), .B(new_n298), .C1(G169), .C2(new_n272), .ZN(new_n299));
  XOR2_X1   g0099(.A(new_n299), .B(KEYINPUT67), .Z(new_n300));
  NAND2_X1  g0100(.A1(new_n235), .A2(G1698), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n262), .B(new_n301), .C1(G226), .C2(G1698), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G97), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n257), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G238), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n258), .B1(new_n259), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT13), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(G200), .B2(new_n309), .ZN(new_n312));
  OR3_X1    g0112(.A1(new_n276), .A2(KEYINPUT71), .A3(G68), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT71), .B1(new_n276), .B2(G68), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(KEYINPUT12), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n281), .A2(G68), .A3(new_n282), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n315), .B(new_n316), .C1(KEYINPUT12), .C2(new_n314), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n317), .A2(KEYINPUT72), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(KEYINPUT72), .ZN(new_n319));
  INV_X1    g0119(.A(new_n284), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n320), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n287), .A2(new_n214), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n280), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT11), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n318), .A2(new_n319), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n312), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n286), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n284), .B1(G20), .B2(G77), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT15), .B(G87), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT68), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n329), .B1(new_n331), .B2(new_n287), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(new_n280), .B1(new_n214), .B2(new_n277), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n281), .A2(G77), .A3(new_n282), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT69), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n279), .B1(G33), .B2(G41), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n262), .A2(G232), .A3(new_n264), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n206), .B2(new_n262), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n270), .A2(new_n305), .A3(new_n264), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n258), .C1(new_n213), .C2(new_n259), .ZN(new_n342));
  INV_X1    g0142(.A(new_n273), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n336), .B(new_n344), .C1(new_n310), .C2(new_n342), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n342), .A2(G179), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n333), .A2(new_n335), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  AND4_X1   g0151(.A1(new_n296), .A2(new_n300), .A3(new_n327), .A4(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT14), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n309), .A2(new_n353), .A3(G169), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n309), .B2(new_n297), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n353), .B1(new_n309), .B2(G169), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n325), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT16), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT74), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n255), .B2(KEYINPUT3), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT73), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n268), .B2(G33), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n268), .A2(KEYINPUT74), .A3(G33), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n255), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n361), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT7), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(G20), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n367), .B1(new_n262), .B2(G20), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n247), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G58), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n247), .ZN(new_n373));
  OAI21_X1  g0173(.A(G20), .B1(new_n373), .B2(new_n201), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n284), .A2(G159), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n359), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT7), .B1(new_n270), .B2(new_n210), .ZN(new_n378));
  AOI211_X1 g0178(.A(new_n367), .B(G20), .C1(new_n267), .C2(new_n269), .ZN(new_n379));
  OAI21_X1  g0179(.A(G68), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n376), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(KEYINPUT16), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n377), .A2(new_n280), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n281), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n328), .A2(new_n282), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n384), .A2(new_n385), .B1(new_n276), .B2(new_n328), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n264), .A2(G226), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n262), .B(new_n390), .C1(G223), .C2(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n337), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n258), .B1(new_n259), .B2(new_n235), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n348), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n257), .B1(new_n391), .B2(new_n392), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n398), .A2(new_n395), .A3(new_n297), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n388), .A2(new_n389), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n270), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n370), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n376), .B1(new_n404), .B2(G68), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n290), .B1(new_n405), .B2(KEYINPUT16), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n386), .B1(new_n406), .B2(new_n377), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT18), .B1(new_n407), .B2(new_n400), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n394), .A2(new_n396), .A3(new_n310), .ZN(new_n414));
  INV_X1    g0214(.A(G200), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n398), .B2(new_n395), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n413), .B1(new_n407), .B2(new_n417), .ZN(new_n418));
  AND4_X1   g0218(.A1(new_n383), .A2(new_n387), .A3(new_n417), .A4(new_n410), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n358), .A2(new_n409), .A3(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n267), .A2(new_n269), .A3(new_n210), .A4(G68), .ZN(new_n422));
  OR2_X1    g0222(.A1(KEYINPUT76), .A2(G97), .ZN(new_n423));
  NAND2_X1  g0223(.A1(KEYINPUT76), .A2(G97), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n287), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n422), .B1(new_n425), .B2(KEYINPUT19), .ZN(new_n426));
  XOR2_X1   g0226(.A(KEYINPUT76), .B(G97), .Z(new_n427));
  NOR2_X1   g0227(.A1(G87), .A2(G107), .ZN(new_n428));
  NAND3_X1  g0228(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n427), .A2(new_n428), .B1(new_n210), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n280), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n209), .A2(G33), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n281), .A2(KEYINPUT84), .A3(G87), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT84), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n276), .A2(new_n432), .A3(new_n279), .A4(new_n278), .ZN(new_n435));
  INV_X1    g0235(.A(G87), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n331), .A2(new_n277), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n431), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n209), .A2(G45), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n442), .A2(G250), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n257), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n257), .A2(G274), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n305), .A2(new_n264), .ZN(new_n447));
  INV_X1    g0247(.A(G244), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G1698), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n267), .A2(new_n447), .A3(new_n269), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G116), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT83), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n257), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(KEYINPUT83), .A3(new_n451), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n446), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G190), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n441), .B(new_n457), .C1(new_n456), .C2(new_n273), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n297), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n431), .B(new_n439), .C1(new_n435), .C2(new_n331), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n459), .B(new_n460), .C1(G169), .C2(new_n456), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n264), .A2(KEYINPUT4), .A3(G244), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT80), .B1(new_n270), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n267), .A2(new_n269), .A3(G250), .A4(G1698), .ZN(new_n466));
  NAND2_X1  g0266(.A1(KEYINPUT4), .A2(G244), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1698), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n267), .A4(new_n269), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n267), .A2(new_n269), .A3(G244), .A4(new_n264), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT4), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n337), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  INV_X1    g0277(.A(new_n442), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(G257), .A3(new_n257), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n477), .A2(new_n257), .A3(G274), .A4(new_n478), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n476), .A2(new_n483), .A3(new_n297), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT82), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n466), .A2(new_n465), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n486), .A2(new_n474), .A3(new_n464), .A4(new_n470), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n482), .B1(new_n487), .B2(new_n337), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT82), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(new_n297), .ZN(new_n490));
  INV_X1    g0290(.A(new_n488), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n485), .A2(new_n490), .B1(new_n348), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n206), .B1(new_n369), .B2(new_n370), .ZN(new_n493));
  AND2_X1   g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  NOR2_X1   g0294(.A1(G97), .A2(G107), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT77), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT77), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G97), .A2(G107), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n207), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n423), .A2(new_n424), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(KEYINPUT6), .A3(new_n206), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n210), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n284), .A2(G77), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n493), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT78), .B1(new_n507), .B2(new_n290), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT78), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n378), .B1(new_n366), .B2(new_n368), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n505), .B1(new_n510), .B2(new_n206), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n280), .C1(new_n511), .C2(new_n504), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n435), .A2(G97), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(G97), .B2(new_n277), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n514), .B(KEYINPUT79), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n508), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n492), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n488), .A2(new_n310), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(G200), .B2(new_n488), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(new_n508), .A3(new_n515), .A4(new_n512), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(KEYINPUT81), .A3(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n508), .A2(new_n515), .A3(new_n512), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT81), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(new_n519), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n462), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n337), .B1(new_n478), .B2(new_n477), .ZN(new_n526));
  INV_X1    g0326(.A(new_n479), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n257), .A2(G274), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n526), .A2(G270), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n262), .A2(G264), .A3(G1698), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n262), .A2(G257), .A3(new_n264), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n270), .A2(G303), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n337), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n529), .A2(new_n534), .A3(G179), .ZN(new_n535));
  MUX2_X1   g0335(.A(new_n276), .B(new_n435), .S(G116), .Z(new_n536));
  NAND2_X1  g0336(.A1(new_n465), .A2(new_n210), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n427), .B2(G33), .ZN(new_n539));
  INV_X1    g0339(.A(G116), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n278), .A2(new_n279), .B1(G20), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT20), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(G33), .B1(new_n423), .B2(new_n424), .ZN(new_n543));
  OAI211_X1 g0343(.A(KEYINPUT20), .B(new_n541), .C1(new_n543), .C2(new_n537), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n536), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n535), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n348), .B1(new_n529), .B2(new_n534), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n548), .A2(KEYINPUT21), .A3(new_n546), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT21), .B1(new_n548), .B2(new_n546), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n262), .A2(new_n210), .A3(G87), .ZN(new_n553));
  XNOR2_X1  g0353(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n287), .A2(new_n540), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT86), .B1(new_n210), .B2(G107), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT23), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT23), .ZN(new_n560));
  OAI211_X1 g0360(.A(KEYINPUT86), .B(new_n560), .C1(new_n210), .C2(G107), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n557), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n262), .A2(new_n554), .A3(new_n210), .A4(G87), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n556), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT24), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT24), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n556), .A2(new_n562), .A3(new_n566), .A4(new_n563), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n290), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n277), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT25), .B1(new_n277), .B2(new_n206), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n569), .A2(new_n570), .B1(new_n206), .B2(new_n435), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n267), .A2(new_n269), .A3(G257), .A4(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n267), .A2(new_n269), .A3(G250), .A4(new_n264), .ZN(new_n574));
  INV_X1    g0374(.A(G294), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n574), .C1(new_n255), .C2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(new_n337), .B1(new_n526), .B2(G264), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n577), .A2(G190), .A3(new_n481), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n415), .B1(new_n577), .B2(new_n481), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n529), .A2(new_n534), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n546), .B1(G200), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n479), .A2(G270), .A3(new_n257), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n481), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n337), .B2(new_n533), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G190), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n572), .A2(new_n580), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n577), .A2(new_n481), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n348), .ZN(new_n589));
  OAI221_X1 g0389(.A(new_n589), .B1(G179), .B2(new_n588), .C1(new_n568), .C2(new_n571), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n552), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n421), .A2(new_n525), .A3(new_n591), .ZN(G372));
  INV_X1    g0392(.A(KEYINPUT89), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n440), .A2(KEYINPUT88), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT88), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n431), .A2(new_n438), .A3(new_n439), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n456), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(KEYINPUT87), .A3(new_n343), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT87), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n456), .B2(new_n273), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n597), .A2(new_n457), .A3(new_n599), .A4(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n602), .A2(new_n492), .A3(new_n516), .A4(new_n461), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n461), .B1(new_n603), .B2(KEYINPUT26), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT26), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n491), .A2(new_n348), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n489), .A2(new_n476), .A3(new_n483), .A4(new_n297), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n489), .B1(new_n488), .B2(new_n297), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n522), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n462), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n605), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n593), .B1(new_n604), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n602), .A2(new_n461), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(new_n610), .A3(new_n605), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT26), .B1(new_n517), .B2(new_n462), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(KEYINPUT89), .A4(new_n461), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n488), .A2(G200), .ZN(new_n618));
  AOI211_X1 g0418(.A(G190), .B(new_n482), .C1(new_n487), .C2(new_n337), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT81), .B1(new_n516), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n524), .B1(new_n610), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n552), .A2(new_n590), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n572), .A2(new_n580), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .A4(new_n614), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n613), .A2(new_n617), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n421), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n350), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n327), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n420), .B1(new_n629), .B2(new_n357), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT90), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n389), .B1(new_n388), .B2(new_n401), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n407), .A2(KEYINPUT18), .A3(new_n400), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n402), .A2(new_n408), .A3(KEYINPUT90), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n296), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n637), .A2(new_n300), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n627), .A2(new_n638), .ZN(G369));
  NAND3_X1  g0439(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT27), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(G213), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n546), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n552), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n582), .A2(new_n586), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n649), .B(KEYINPUT91), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G330), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n590), .A2(new_n645), .ZN(new_n653));
  INV_X1    g0453(.A(new_n645), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n624), .B1(new_n572), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n653), .B1(new_n590), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n552), .A2(new_n645), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT92), .Z(new_n659));
  AOI21_X1  g0459(.A(new_n653), .B1(new_n659), .B2(new_n656), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n227), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G1), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n427), .A2(new_n540), .A3(new_n428), .ZN(new_n666));
  OAI22_X1  g0466(.A1(new_n665), .A2(new_n666), .B1(new_n224), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  AND4_X1   g0468(.A1(new_n552), .A2(new_n587), .A3(new_n590), .A4(new_n654), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n622), .A2(new_n611), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT95), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n525), .A2(KEYINPUT95), .A3(new_n669), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT31), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n456), .A2(new_n476), .A3(new_n483), .A4(new_n577), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n585), .A2(G179), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT30), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n454), .A2(new_n455), .ZN(new_n679));
  INV_X1    g0479(.A(new_n446), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n679), .A2(new_n680), .A3(new_n577), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT30), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(new_n488), .A4(new_n535), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n585), .A2(new_n456), .A3(G179), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n488), .B1(new_n481), .B2(new_n577), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n678), .A2(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT94), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n645), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n678), .A2(new_n683), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n685), .A2(new_n684), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n689), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n675), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n690), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n645), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT93), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n674), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n614), .A2(new_n623), .A3(new_n624), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n521), .B2(new_n524), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n603), .A2(KEYINPUT26), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n610), .A2(new_n605), .A3(new_n611), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n701), .A3(new_n461), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n654), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n626), .A2(new_n654), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(KEYINPUT29), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n697), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT96), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT96), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n668), .B1(new_n710), .B2(G1), .ZN(G364));
  AND2_X1   g0511(.A1(new_n210), .A2(G13), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n209), .B1(new_n712), .B2(G45), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n663), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n652), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(G330), .B2(new_n650), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G13), .A2(G33), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G20), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n649), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n715), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n662), .A2(new_n270), .ZN(new_n723));
  OR2_X1    g0523(.A1(G355), .A2(KEYINPUT97), .ZN(new_n724));
  NAND2_X1  g0524(.A1(G355), .A2(KEYINPUT97), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n662), .A2(new_n262), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(G45), .B2(new_n224), .ZN(new_n728));
  INV_X1    g0528(.A(G45), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n251), .A2(new_n729), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n726), .B1(G116), .B2(new_n227), .C1(new_n728), .C2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n279), .B1(G20), .B2(new_n348), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n720), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n722), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G179), .A2(G200), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n210), .B1(new_n735), .B2(G190), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n736), .A2(KEYINPUT102), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(KEYINPUT102), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(G20), .A2(G179), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT98), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G190), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n415), .ZN(new_n744));
  AOI22_X1  g0544(.A1(new_n740), .A2(G294), .B1(new_n744), .B2(G326), .ZN(new_n745));
  INV_X1    g0545(.A(G322), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n743), .A2(G200), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n742), .A2(new_n310), .A3(new_n415), .ZN(new_n750));
  INV_X1    g0550(.A(G311), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n210), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n735), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n262), .B(new_n752), .C1(G329), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n273), .A2(G179), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT99), .ZN(new_n758));
  INV_X1    g0558(.A(new_n753), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G283), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n758), .A2(new_n210), .A3(new_n310), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G303), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n756), .B1(new_n761), .B2(new_n762), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n742), .A2(new_n310), .A3(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(KEYINPUT101), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n767), .A2(KEYINPUT101), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n749), .B(new_n766), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n763), .A2(G87), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n760), .A2(G107), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n775), .A2(new_n262), .A3(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT100), .Z(new_n778));
  INV_X1    g0578(.A(G159), .ZN(new_n779));
  OR3_X1    g0579(.A1(new_n754), .A2(KEYINPUT32), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(KEYINPUT32), .B1(new_n754), .B2(new_n779), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n780), .B(new_n781), .C1(new_n739), .C2(new_n205), .ZN(new_n782));
  INV_X1    g0582(.A(new_n750), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G50), .A2(new_n744), .B1(new_n783), .B2(G77), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n372), .B2(new_n748), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n782), .B(new_n785), .C1(G68), .C2(new_n772), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n774), .B1(new_n778), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n732), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n721), .B(new_n734), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n717), .A2(new_n789), .ZN(G396));
  OAI21_X1  g0590(.A(new_n345), .B1(new_n336), .B2(new_n654), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n350), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n628), .A2(new_n654), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n705), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n794), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n626), .A2(new_n654), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n697), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n715), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n697), .A2(new_n795), .A3(new_n797), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n788), .A2(new_n719), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n715), .B1(new_n802), .B2(G77), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT103), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G294), .A2(new_n747), .B1(new_n744), .B2(G303), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n540), .B2(new_n750), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n760), .A2(G87), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n270), .B1(new_n754), .B2(new_n751), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n740), .B2(G97), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(new_n764), .C2(new_n206), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n806), .B(new_n810), .C1(G283), .C2(new_n772), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G137), .A2(new_n744), .B1(new_n783), .B2(G159), .ZN(new_n812));
  INV_X1    g0612(.A(G143), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n813), .B2(new_n748), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G150), .B2(new_n772), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT34), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n760), .A2(G68), .ZN(new_n817));
  INV_X1    g0617(.A(G132), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n262), .B1(new_n754), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n740), .B2(G58), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n817), .B(new_n820), .C1(new_n764), .C2(new_n202), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n815), .B2(KEYINPUT34), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n811), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n804), .B1(new_n823), .B2(new_n788), .C1(new_n796), .C2(new_n719), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n801), .A2(new_n824), .ZN(G384));
  NAND2_X1  g0625(.A1(new_n501), .A2(new_n503), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT35), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n225), .A2(new_n540), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n826), .B2(KEYINPUT35), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT104), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n827), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT36), .ZN(new_n833));
  OR3_X1    g0633(.A1(new_n373), .A2(new_n224), .A3(new_n214), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n209), .B(G13), .C1(new_n834), .C2(new_n246), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n693), .A2(KEYINPUT94), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n686), .A2(new_n687), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n837), .A2(KEYINPUT31), .A3(new_n645), .A4(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n692), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT95), .B1(new_n525), .B2(new_n669), .ZN(new_n841));
  AND4_X1   g0641(.A1(KEYINPUT95), .A2(new_n622), .A3(new_n611), .A4(new_n669), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n643), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT16), .B1(new_n380), .B2(new_n381), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT106), .B1(new_n845), .B2(new_n290), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT106), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n847), .B(new_n280), .C1(new_n405), .C2(KEYINPUT16), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n846), .A2(new_n382), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n387), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n844), .B(new_n850), .C1(new_n420), .C2(new_n409), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n383), .A2(new_n387), .A3(new_n417), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n850), .B2(new_n401), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n850), .A2(new_n844), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n388), .A2(new_n401), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n388), .A2(new_n844), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n383), .A2(new_n387), .A3(new_n417), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n851), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n851), .B(KEYINPUT38), .C1(new_n856), .C2(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n357), .A2(KEYINPUT105), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT105), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n868), .B(new_n325), .C1(new_n355), .C2(new_n356), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n326), .A2(new_n654), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n312), .B2(new_n326), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n867), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n870), .B1(new_n355), .B2(new_n356), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n794), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n843), .A2(new_n866), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT40), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT110), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(KEYINPUT110), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n865), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT108), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n418), .B2(new_n419), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n407), .A2(new_n417), .A3(new_n410), .ZN(new_n885));
  OAI211_X1 g0685(.A(KEYINPUT108), .B(new_n885), .C1(new_n853), .C2(new_n413), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n634), .A2(new_n884), .A3(new_n635), .A4(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n858), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n882), .B1(new_n893), .B2(KEYINPUT109), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT109), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n887), .A2(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(KEYINPUT38), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n876), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n843), .A2(new_n874), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n881), .A2(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n421), .A2(new_n843), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(G330), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT107), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n872), .A2(new_n873), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  AOI221_X4 g0708(.A(new_n908), .B1(new_n865), .B2(new_n864), .C1(new_n797), .C2(new_n793), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n844), .B1(new_n634), .B2(new_n635), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n908), .B1(new_n797), .B2(new_n793), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n912), .B2(new_n866), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT107), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n893), .A2(KEYINPUT109), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(new_n897), .A3(new_n865), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n645), .B1(new_n867), .B2(new_n869), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n866), .A2(new_n917), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n911), .A2(new_n914), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n706), .A2(new_n421), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n638), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n923), .B(new_n926), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n905), .A2(new_n927), .B1(new_n209), .B2(new_n712), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n905), .A2(new_n927), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n836), .B1(new_n928), .B2(new_n929), .ZN(G367));
  NOR2_X1   g0730(.A1(new_n597), .A2(new_n654), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n614), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n461), .B2(new_n932), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT43), .Z(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n521), .A2(new_n524), .B1(new_n516), .B2(new_n645), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n517), .A2(new_n654), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT111), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n517), .B1(new_n941), .B2(new_n590), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n654), .ZN(new_n943));
  INV_X1    g0743(.A(new_n939), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n656), .A3(new_n659), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT42), .Z(new_n946));
  AOI21_X1  g0746(.A(new_n936), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT112), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n943), .A2(new_n946), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n948), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n947), .A2(KEYINPUT112), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT113), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n953), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT113), .ZN(new_n956));
  INV_X1    g0756(.A(new_n949), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n950), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n955), .A2(new_n956), .A3(new_n958), .A4(new_n948), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n657), .A2(new_n941), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n954), .A2(new_n961), .A3(new_n959), .ZN(new_n964));
  INV_X1    g0764(.A(new_n657), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(KEYINPUT114), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n660), .A2(new_n944), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT45), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n660), .A2(new_n944), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n966), .B(new_n971), .Z(new_n972));
  XNOR2_X1  g0772(.A(new_n659), .B(new_n656), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n651), .B(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n972), .A2(new_n975), .B1(new_n708), .B2(new_n709), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n663), .B(KEYINPUT41), .Z(new_n977));
  OAI21_X1  g0777(.A(new_n713), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n963), .A2(new_n964), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n727), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n733), .B1(new_n227), .B2(new_n331), .C1(new_n980), .C2(new_n241), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n981), .A2(new_n715), .ZN(new_n982));
  INV_X1    g0782(.A(new_n720), .ZN(new_n983));
  INV_X1    g0783(.A(new_n744), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n984), .A2(new_n751), .B1(new_n206), .B2(new_n739), .ZN(new_n985));
  XNOR2_X1  g0785(.A(KEYINPUT115), .B(G317), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n262), .B1(new_n755), .B2(new_n986), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n765), .B2(new_n748), .C1(new_n761), .C2(new_n427), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n985), .B(new_n988), .C1(G283), .C2(new_n783), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n763), .A2(G116), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT46), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n989), .B(new_n991), .C1(new_n575), .C2(new_n771), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n739), .A2(new_n247), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n984), .A2(new_n813), .B1(new_n202), .B2(new_n750), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(new_n772), .C2(G159), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n763), .A2(G58), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n760), .A2(G77), .ZN(new_n997));
  INV_X1    g0797(.A(G137), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n262), .B1(new_n754), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n747), .B2(G150), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n992), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(KEYINPUT116), .B(KEYINPUT47), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n982), .B1(new_n983), .B2(new_n934), .C1(new_n1004), .C2(new_n788), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n979), .A2(new_n1005), .ZN(G387));
  AOI21_X1  g0806(.A(new_n974), .B1(new_n708), .B2(new_n709), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n708), .A2(new_n709), .A3(new_n974), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n663), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n975), .A2(new_n714), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n984), .A2(new_n746), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n747), .B2(new_n986), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n765), .B2(new_n750), .C1(new_n751), .C2(new_n771), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT48), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n764), .A2(new_n575), .B1(new_n739), .B2(new_n762), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(KEYINPUT49), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n262), .B1(new_n755), .B2(G326), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n540), .C2(new_n761), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT49), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n764), .A2(new_n214), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n739), .A2(new_n331), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n270), .B1(new_n755), .B2(G150), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n761), .C2(new_n205), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G50), .A2(new_n747), .B1(new_n783), .B2(G68), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n779), .B2(new_n984), .C1(new_n771), .C2(new_n286), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1024), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n732), .B1(new_n1023), .B2(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n238), .A2(new_n729), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1032), .A2(new_n727), .B1(new_n666), .B2(new_n723), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n328), .A2(new_n202), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT50), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n729), .B1(new_n247), .B2(new_n214), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1035), .A2(new_n666), .A3(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1033), .A2(new_n1037), .B1(G107), .B2(new_n227), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n722), .B1(new_n1038), .B2(new_n733), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1031), .B(new_n1039), .C1(new_n656), .C2(new_n983), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1011), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1010), .A2(new_n1041), .ZN(G393));
  XNOR2_X1  g0842(.A(new_n971), .B(new_n657), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n714), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n733), .B1(new_n227), .B2(new_n427), .C1(new_n980), .C2(new_n245), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n715), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G150), .A2(new_n744), .B1(new_n747), .B2(G159), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT51), .Z(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n202), .B2(new_n771), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n262), .B1(new_n813), .B2(new_n754), .C1(new_n750), .C2(new_n286), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n739), .A2(new_n214), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n807), .B(new_n1052), .C1(new_n764), .C2(new_n247), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n772), .A2(G303), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n270), .B1(new_n746), .B2(new_n754), .C1(new_n750), .C2(new_n575), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G116), .B2(new_n740), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n763), .A2(G283), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1054), .A2(new_n776), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G311), .A2(new_n747), .B1(new_n744), .B2(G317), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1049), .A2(new_n1053), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1046), .B1(new_n1061), .B2(new_n732), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n940), .B2(new_n983), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n966), .B(new_n971), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n663), .B1(new_n1008), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1043), .A2(new_n1007), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1044), .B(new_n1063), .C1(new_n1065), .C2(new_n1066), .ZN(G390));
  AOI21_X1  g0867(.A(new_n919), .B1(new_n894), .B2(new_n897), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n703), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1069), .A2(new_n792), .B1(new_n628), .B2(new_n654), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1068), .B1(new_n1070), .B2(new_n908), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n912), .A2(new_n919), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n920), .B1(new_n916), .B2(new_n917), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n843), .ZN(new_n1075));
  INV_X1    g0875(.A(G330), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n794), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1075), .A2(new_n908), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n696), .A2(new_n907), .A3(new_n1077), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1071), .B(new_n1081), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n714), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT118), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n421), .A2(G330), .A3(new_n843), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT117), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n902), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n925), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n797), .A2(new_n793), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n907), .B1(new_n696), .B2(new_n1077), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1079), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n908), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n1081), .A3(new_n1070), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1091), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1086), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1080), .A2(new_n1091), .A3(new_n1097), .A4(new_n1082), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n663), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n715), .B1(new_n802), .B2(new_n328), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n817), .B1(new_n575), .B2(new_n754), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1103), .B(KEYINPUT120), .Z(new_n1104));
  AOI21_X1  g0904(.A(new_n262), .B1(new_n763), .B2(G87), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1105), .A2(KEYINPUT119), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n984), .A2(new_n762), .B1(new_n427), .B2(new_n750), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1051), .B(new_n1107), .C1(G116), .C2(new_n747), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1105), .A2(KEYINPUT119), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n772), .A2(G107), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n763), .A2(G150), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT53), .ZN(new_n1113));
  INV_X1    g0913(.A(G128), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1114), .A2(new_n984), .B1(new_n748), .B2(new_n818), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT54), .B(G143), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1115), .B1(new_n783), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n760), .A2(G50), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n772), .A2(G137), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n739), .A2(new_n779), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n270), .B(new_n1121), .C1(G125), .C2(new_n755), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .A4(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1104), .A2(new_n1111), .B1(new_n1113), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1102), .B1(new_n1124), .B2(new_n732), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n1073), .B2(new_n719), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1085), .A2(new_n1101), .A3(new_n1126), .ZN(G378));
  OAI21_X1  g0927(.A(new_n922), .B1(new_n913), .B2(KEYINPUT107), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n909), .A2(new_n906), .A3(new_n910), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1076), .B1(new_n898), .B2(new_n899), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n296), .A2(new_n299), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n291), .A2(new_n844), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1134), .B(new_n1135), .Z(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT110), .B1(new_n875), .B2(new_n876), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n875), .A2(KEYINPUT110), .A3(new_n876), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1131), .B(new_n1136), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1136), .B1(new_n881), .B2(new_n1131), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1130), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1136), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1138), .A2(new_n1137), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n900), .A2(G330), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1146), .A2(new_n923), .A3(new_n1139), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1142), .A2(KEYINPUT122), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT122), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(new_n923), .A3(new_n1149), .A4(new_n1139), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n714), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n715), .B1(new_n802), .B2(G50), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n270), .B2(new_n256), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n256), .B(new_n270), .C1(new_n754), .C2(new_n762), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1024), .A2(new_n993), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n747), .A2(G107), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n331), .B2(new_n750), .C1(new_n984), .C2(new_n540), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G97), .B2(new_n772), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1156), .B(new_n1159), .C1(new_n372), .C2(new_n761), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT58), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1154), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n740), .A2(G150), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n748), .A2(new_n1114), .B1(new_n998), .B2(new_n750), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(G125), .C2(new_n744), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n818), .B2(new_n771), .C1(new_n764), .C2(new_n1116), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G33), .B(G41), .C1(new_n755), .C2(G124), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1167), .B(new_n1168), .C1(new_n779), .C2(new_n761), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1162), .B1(new_n1161), .B2(new_n1160), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1152), .B1(new_n1171), .B2(new_n732), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1143), .B2(new_n719), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT121), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1151), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT123), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT123), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1151), .A2(new_n1177), .A3(new_n1174), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT124), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1142), .A2(new_n1179), .A3(new_n1147), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1100), .B2(new_n1091), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1146), .A2(new_n923), .A3(KEYINPUT124), .A4(new_n1139), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1180), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1184), .A2(new_n663), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1100), .A2(new_n1091), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1148), .A2(new_n1150), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1181), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1176), .A2(new_n1178), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(G375));
  NAND2_X1  g0990(.A1(new_n908), .A2(new_n718), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n715), .B1(new_n802), .B2(G68), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n262), .B1(new_n754), .B2(new_n1114), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n744), .B2(G132), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1194), .B1(new_n761), .B2(new_n372), .C1(new_n764), .C2(new_n779), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n740), .A2(G50), .B1(G150), .B2(new_n783), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n998), .B2(new_n748), .C1(new_n771), .C2(new_n1116), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(G294), .A2(new_n744), .B1(new_n783), .B2(G107), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n762), .B2(new_n748), .C1(new_n771), .C2(new_n540), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n763), .A2(G97), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n262), .B1(new_n755), .B2(G303), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1200), .A2(new_n997), .A3(new_n1025), .A4(new_n1201), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n1195), .A2(new_n1197), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1192), .B1(new_n1203), .B2(new_n732), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1097), .A2(new_n714), .B1(new_n1191), .B2(new_n1204), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n977), .B(KEYINPUT125), .Z(new_n1206));
  NAND2_X1  g1006(.A1(new_n1098), .A2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1091), .A2(new_n1097), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1205), .B1(new_n1207), .B2(new_n1208), .ZN(G381));
  INV_X1    g1009(.A(G378), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1189), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(G396), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1010), .A2(new_n1212), .A3(new_n1041), .ZN(new_n1213));
  OR4_X1    g1013(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1213), .ZN(new_n1214));
  OR3_X1    g1014(.A1(new_n1211), .A2(G387), .A3(new_n1214), .ZN(G407));
  OAI211_X1 g1015(.A(G407), .B(G213), .C1(G343), .C2(new_n1211), .ZN(G409));
  AOI21_X1  g1016(.A(new_n1212), .B1(new_n1010), .B2(new_n1041), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(G390), .A3(new_n1213), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1044), .A2(new_n1063), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n664), .B1(new_n972), .B2(new_n1007), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1066), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1220), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1010), .A2(new_n1212), .A3(new_n1041), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1223), .B1(new_n1224), .B2(new_n1217), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1219), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(G387), .A2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n979), .A2(new_n1219), .A3(new_n1225), .A4(new_n1005), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1188), .A2(new_n663), .A3(new_n1184), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1177), .B1(new_n1151), .B2(new_n1174), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1151), .A2(new_n1177), .A3(new_n1174), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1230), .B(G378), .C1(new_n1231), .C2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1180), .A2(new_n714), .A3(new_n1183), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1206), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1174), .B(new_n1234), .C1(new_n1187), .C2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1210), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1233), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n644), .A2(G213), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1208), .A2(KEYINPUT60), .A3(new_n1098), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n663), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1208), .B1(KEYINPUT60), .B2(new_n1098), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1205), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n801), .A3(new_n824), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G384), .B(new_n1205), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1238), .A2(new_n1239), .A3(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT126), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1238), .A2(KEYINPUT126), .A3(new_n1239), .A4(new_n1247), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT62), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1239), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(G2897), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1246), .B(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1237), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1189), .B2(G378), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n1257), .B2(new_n1253), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1253), .B(new_n1246), .C1(new_n1233), .C2(new_n1237), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1258), .B(new_n1259), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1229), .B1(new_n1252), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1250), .A2(new_n1264), .A3(new_n1251), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1229), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1261), .A2(KEYINPUT63), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1263), .A2(new_n1269), .ZN(G405));
  AND3_X1   g1070(.A1(new_n1227), .A2(new_n1247), .A3(new_n1228), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1247), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT127), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1229), .A2(new_n1246), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT127), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1227), .A2(new_n1247), .A3(new_n1228), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G375), .A2(new_n1210), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1233), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1273), .A2(new_n1277), .A3(new_n1233), .A4(new_n1279), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G402));
endmodule


