//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT67), .A2(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(G143), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n189), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n192), .A2(new_n193), .A3(G128), .A4(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n197), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n190), .A2(new_n191), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(new_n199), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n196), .B1(new_n198), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G137), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n204), .A2(G137), .ZN(new_n207));
  OAI21_X1  g021(.A(G131), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n204), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n205), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n208), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n210), .A2(new_n205), .A3(new_n212), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n214), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n192), .A2(KEYINPUT0), .A3(G128), .A4(new_n195), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT0), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(new_n197), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(KEYINPUT66), .A2(KEYINPUT0), .A3(G128), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT66), .B1(KEYINPUT0), .B2(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(G143), .B1(new_n190), .B2(new_n191), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n225), .B(new_n228), .C1(new_n229), .C2(new_n200), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n219), .A2(new_n220), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n216), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g046(.A(G116), .B(G119), .Z(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n234), .A2(new_n235), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT69), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n234), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT68), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n234), .A2(new_n235), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .A4(new_n233), .ZN(new_n243));
  XNOR2_X1  g057(.A(G116), .B(G119), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n238), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n232), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT28), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n230), .A2(new_n220), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n249), .A2(new_n219), .B1(new_n203), .B2(new_n215), .ZN(new_n250));
  INV_X1    g064(.A(new_n246), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n232), .A2(new_n246), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n248), .B1(new_n254), .B2(KEYINPUT28), .ZN(new_n255));
  NOR2_X1   g069(.A1(G237), .A2(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G210), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n257), .B(KEYINPUT27), .Z(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n261), .A2(KEYINPUT29), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT75), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n255), .A2(new_n266), .A3(new_n262), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n248), .ZN(new_n269));
  XOR2_X1   g083(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n270));
  NAND2_X1  g084(.A1(new_n254), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n271), .A3(new_n261), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n273));
  OR2_X1    g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n275), .B(new_n276), .C1(new_n250), .C2(KEYINPUT64), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT30), .B1(new_n250), .B2(new_n275), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT70), .B1(new_n232), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n246), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n252), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n260), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT29), .B1(new_n272), .B2(new_n273), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n274), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n268), .B1(new_n286), .B2(KEYINPUT74), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n274), .A2(new_n284), .A3(new_n288), .A4(new_n285), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n187), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n282), .A2(new_n261), .A3(new_n252), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT31), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n269), .A2(new_n271), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n260), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n247), .B1(new_n281), .B2(new_n246), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT31), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n261), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n292), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G472), .A2(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(KEYINPUT32), .A3(new_n299), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT32), .B1(new_n298), .B2(new_n299), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n290), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT22), .B(G137), .ZN(new_n309));
  INV_X1    g123(.A(G221), .ZN(new_n310));
  INV_X1    g124(.A(G234), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n310), .A2(new_n311), .A3(G953), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n309), .B(new_n312), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(KEYINPUT77), .Z(new_n316));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(G128), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT23), .B1(new_n197), .B2(G119), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n197), .A2(KEYINPUT78), .A3(G119), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(G119), .B(G128), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT24), .B(G110), .Z(new_n325));
  OAI22_X1  g139(.A1(new_n323), .A2(G110), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT79), .B(G125), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  INV_X1    g142(.A(G140), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(G125), .A2(G140), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n327), .B2(G140), .ZN(new_n332));
  OAI211_X1 g146(.A(G146), .B(new_n330), .C1(new_n332), .C2(new_n328), .ZN(new_n333));
  AND2_X1   g147(.A1(KEYINPUT67), .A2(G146), .ZN(new_n334));
  NOR2_X1   g148(.A1(KEYINPUT67), .A2(G146), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(G125), .A2(G140), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n338), .A2(new_n331), .A3(new_n339), .ZN(new_n340));
  OR2_X1    g154(.A1(G125), .A2(G140), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT80), .B1(new_n341), .B2(new_n337), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n336), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n326), .A2(new_n333), .A3(new_n343), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n323), .A2(G110), .B1(new_n324), .B2(new_n325), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n330), .B1(new_n332), .B2(new_n328), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n189), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n333), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(KEYINPUT81), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n344), .B2(new_n349), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n314), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n313), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT25), .B1(new_n356), .B2(G902), .ZN(new_n357));
  OAI21_X1  g171(.A(G217), .B1(new_n311), .B2(G902), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT76), .ZN(new_n359));
  AOI21_X1  g173(.A(G902), .B1(new_n354), .B2(new_n355), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n359), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n356), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT82), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n357), .A2(new_n362), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n370));
  INV_X1    g184(.A(new_n367), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n308), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G210), .B1(G237), .B2(G902), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT91), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n377));
  INV_X1    g191(.A(G104), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n378), .B2(G107), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT3), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G104), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n378), .A2(G107), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n379), .A2(new_n382), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n378), .A2(G107), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n381), .A2(G104), .ZN(new_n387));
  OAI21_X1  g201(.A(G101), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n318), .A3(G116), .ZN(new_n391));
  OAI211_X1 g205(.A(G113), .B(new_n391), .C1(new_n233), .C2(new_n390), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n389), .A2(new_n245), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n379), .A2(new_n382), .A3(new_n384), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(G101), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n394), .A2(KEYINPUT83), .A3(new_n395), .A4(G101), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n395), .B1(new_n394), .B2(G101), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n398), .A2(new_n399), .B1(new_n385), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n393), .B1(new_n401), .B2(new_n246), .ZN(new_n402));
  XNOR2_X1  g216(.A(G110), .B(G122), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n377), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n246), .ZN(new_n405));
  INV_X1    g219(.A(new_n393), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n403), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  XOR2_X1   g224(.A(KEYINPUT79), .B(G125), .Z(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n230), .B2(new_n220), .ZN(new_n412));
  OAI22_X1  g226(.A1(new_n412), .A2(KEYINPUT90), .B1(new_n203), .B2(new_n327), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G953), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G224), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(KEYINPUT90), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n417), .ZN(new_n419));
  OAI211_X1 g233(.A(G224), .B(new_n415), .C1(new_n419), .C2(new_n413), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n407), .A2(new_n377), .A3(new_n408), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n410), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n402), .A2(new_n403), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT7), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n419), .B2(new_n413), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n403), .B(KEYINPUT8), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n389), .B1(new_n245), .B2(new_n392), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n393), .B2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n420), .A2(new_n424), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n414), .A2(KEYINPUT7), .A3(new_n416), .A4(new_n417), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n265), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n376), .B1(new_n423), .B2(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n424), .A2(new_n426), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n435), .A2(new_n420), .A3(new_n431), .A4(new_n429), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n410), .A2(new_n421), .A3(new_n422), .ZN(new_n437));
  INV_X1    g251(.A(new_n376), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n265), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  XNOR2_X1  g255(.A(G113), .B(G122), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(new_n378), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G237), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n415), .A3(G214), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n199), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n256), .A2(G143), .A3(G214), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G131), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n213), .A3(new_n448), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n333), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT19), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n340), .B2(new_n342), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT19), .B(new_n341), .C1(new_n411), .C2(new_n329), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n336), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT93), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT93), .A4(new_n336), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n453), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(KEYINPUT18), .A2(G131), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n449), .B(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n339), .B1(new_n338), .B2(new_n331), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n341), .A2(KEYINPUT80), .A3(new_n337), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n201), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n332), .A2(G146), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(new_n468), .B2(KEYINPUT92), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT92), .B1(new_n332), .B2(G146), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n464), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n444), .B1(new_n461), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n449), .B(new_n462), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n332), .A2(G146), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n343), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n474), .B1(new_n477), .B2(new_n470), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n449), .A2(KEYINPUT17), .A3(G131), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT17), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n450), .A2(new_n480), .A3(new_n451), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n347), .A2(new_n333), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n482), .A3(new_n443), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(G475), .A2(G902), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n441), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n485), .ZN(new_n487));
  AOI211_X1 g301(.A(KEYINPUT20), .B(new_n487), .C1(new_n473), .C2(new_n483), .ZN(new_n488));
  INV_X1    g302(.A(G475), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n478), .A2(new_n482), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n444), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n491), .B2(new_n483), .ZN(new_n492));
  OAI22_X1  g306(.A1(new_n486), .A2(new_n488), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT94), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n199), .A2(G128), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n197), .A2(G143), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n495), .A2(new_n496), .A3(new_n204), .ZN(new_n497));
  INV_X1    g311(.A(G122), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G116), .ZN(new_n499));
  INV_X1    g313(.A(G116), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G122), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G107), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n501), .A3(new_n381), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n497), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT13), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n495), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n496), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n495), .A2(new_n506), .ZN(new_n509));
  OAI21_X1  g323(.A(G134), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n500), .A2(KEYINPUT14), .A3(G122), .ZN(new_n512));
  OAI211_X1 g326(.A(G107), .B(new_n512), .C1(new_n502), .C2(KEYINPUT14), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n204), .B1(new_n495), .B2(new_n496), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n513), .B(new_n504), .C1(new_n497), .C2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n494), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT9), .B(G234), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(G217), .A3(new_n415), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n511), .A2(new_n515), .A3(new_n494), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n522), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n520), .B1(new_n524), .B2(new_n516), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n525), .A3(new_n265), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n528), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n523), .A2(new_n525), .A3(new_n265), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n493), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n415), .A2(G952), .ZN(new_n534));
  NAND2_X1  g348(.A1(G234), .A2(G237), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(G902), .A3(G953), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT21), .B(G898), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(G214), .B1(G237), .B2(G902), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n440), .A2(new_n533), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n310), .B1(new_n519), .B2(new_n265), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G469), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G140), .ZN(new_n549));
  INV_X1    g363(.A(G227), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(G953), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n549), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n385), .A2(new_n388), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n553), .B(new_n196), .C1(new_n198), .C2(new_n202), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n192), .A2(new_n195), .ZN(new_n555));
  OAI21_X1  g369(.A(G128), .B1(new_n200), .B2(new_n193), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT84), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n557), .A2(new_n558), .A3(new_n196), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n389), .B1(new_n558), .B2(new_n196), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT12), .A3(new_n219), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT86), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n219), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT12), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n561), .A2(KEYINPUT86), .A3(KEYINPUT12), .A4(new_n219), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT87), .ZN(new_n570));
  INV_X1    g384(.A(new_n219), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT10), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n553), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n401), .A2(new_n249), .B1(new_n203), .B2(new_n573), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n196), .A2(new_n558), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n194), .B1(new_n336), .B2(G143), .ZN(new_n576));
  INV_X1    g390(.A(new_n556), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n196), .B(new_n558), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(new_n578), .A3(new_n389), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT85), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n579), .A2(new_n580), .A3(new_n572), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n579), .B2(new_n572), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n571), .B(new_n574), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n569), .A2(new_n570), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n570), .B1(new_n569), .B2(new_n583), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n552), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n574), .B1(new_n581), .B2(new_n582), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n219), .ZN(new_n588));
  INV_X1    g402(.A(new_n552), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(new_n583), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n548), .B1(new_n591), .B2(new_n265), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT88), .B(G469), .Z(new_n593));
  NAND2_X1  g407(.A1(new_n583), .A2(new_n589), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT89), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n583), .A2(KEYINPUT89), .A3(new_n589), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n569), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n589), .B1(new_n588), .B2(new_n583), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AOI211_X1 g414(.A(G902), .B(new_n593), .C1(new_n598), .C2(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n545), .B(new_n547), .C1(new_n592), .C2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n374), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  OAI21_X1  g419(.A(new_n547), .B1(new_n592), .B2(new_n601), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI211_X1 g421(.A(KEYINPUT82), .B(new_n367), .C1(new_n362), .C2(new_n357), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n370), .B1(new_n369), .B2(new_n371), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n298), .A2(new_n265), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G472), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n300), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n607), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n375), .B1(new_n423), .B2(new_n433), .ZN(new_n616));
  INV_X1    g430(.A(new_n375), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n436), .A2(new_n437), .A3(new_n265), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n543), .A3(new_n618), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n523), .A2(new_n525), .A3(KEYINPUT33), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT33), .B1(new_n523), .B2(new_n525), .ZN(new_n621));
  OAI211_X1 g435(.A(G478), .B(new_n265), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n526), .A2(new_n527), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n493), .A2(new_n624), .ZN(new_n625));
  NOR4_X1   g439(.A1(new_n615), .A2(new_n541), .A3(new_n619), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT34), .B(G104), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  AND3_X1   g442(.A1(new_n616), .A2(new_n543), .A3(new_n618), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n478), .A2(new_n482), .A3(new_n443), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n459), .A2(new_n460), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n478), .B1(new_n631), .B2(new_n453), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n630), .B1(new_n632), .B2(new_n444), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT20), .B1(new_n633), .B2(new_n487), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT95), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n484), .A2(new_n441), .A3(new_n485), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n491), .A2(new_n483), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n489), .B1(new_n638), .B2(new_n265), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(KEYINPUT95), .B2(new_n488), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n637), .A2(new_n640), .A3(new_n532), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n629), .A2(new_n542), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n615), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n381), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT96), .B(KEYINPUT35), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  XNOR2_X1  g460(.A(new_n350), .B(KEYINPUT81), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n314), .A2(KEYINPUT36), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n647), .A2(KEYINPUT36), .A3(new_n314), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n365), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n369), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n612), .A2(new_n653), .A3(new_n300), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT97), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n612), .A2(new_n653), .A3(KEYINPUT97), .A4(new_n300), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n603), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  NAND2_X1  g474(.A1(new_n287), .A2(new_n289), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G472), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n298), .A2(KEYINPUT32), .A3(new_n299), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n663), .A2(new_n306), .A3(KEYINPUT72), .ZN(new_n664));
  INV_X1    g478(.A(new_n307), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n537), .B1(new_n539), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n641), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n606), .A2(new_n619), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n666), .A2(new_n653), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  XOR2_X1   g487(.A(new_n668), .B(KEYINPUT39), .Z(new_n674));
  OAI211_X1 g488(.A(new_n547), .B(new_n674), .C1(new_n592), .C2(new_n601), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n305), .A2(new_n307), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n283), .A2(new_n261), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n678), .B1(new_n261), .B2(new_n254), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n679), .B2(KEYINPUT100), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(KEYINPUT100), .B2(new_n679), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G472), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n684));
  INV_X1    g498(.A(new_n653), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT99), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n440), .B(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n639), .B1(new_n634), .B2(new_n636), .ZN(new_n689));
  INV_X1    g503(.A(new_n532), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n543), .A2(new_n685), .A3(new_n688), .A4(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n676), .A2(new_n683), .A3(new_n684), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  NAND3_X1  g508(.A1(new_n493), .A2(new_n624), .A3(new_n669), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT101), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n666), .A2(new_n653), .A3(new_n671), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NAND2_X1  g513(.A1(new_n598), .A2(new_n600), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n548), .B1(new_n700), .B2(new_n265), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n601), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n625), .A2(new_n541), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n702), .A2(new_n547), .A3(new_n629), .A4(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n374), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND2_X1  g522(.A1(new_n702), .A2(new_n547), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n642), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n666), .A2(new_n610), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  AND2_X1   g526(.A1(new_n567), .A2(new_n568), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n595), .A2(new_n594), .B1(new_n713), .B2(new_n564), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n599), .B1(new_n714), .B2(new_n597), .ZN(new_n715));
  OAI21_X1  g529(.A(G469), .B1(new_n715), .B2(G902), .ZN(new_n716));
  INV_X1    g530(.A(new_n593), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n700), .A2(new_n265), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n716), .A2(new_n629), .A3(new_n718), .A4(new_n547), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n689), .A2(new_n690), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n719), .A2(new_n720), .A3(new_n541), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n666), .A2(new_n653), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  AOI21_X1  g537(.A(KEYINPUT102), .B1(new_n611), .B2(G472), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n726));
  AOI211_X1 g540(.A(new_n726), .B(new_n187), .C1(new_n298), .C2(new_n265), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n691), .A2(new_n542), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n719), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n363), .A2(new_n367), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n292), .B(new_n297), .C1(new_n261), .C2(new_n255), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n299), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n729), .A2(new_n731), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  OAI211_X1 g550(.A(new_n734), .B(new_n653), .C1(new_n724), .C2(new_n727), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n719), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n697), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  AND3_X1   g555(.A1(new_n434), .A2(new_n439), .A3(new_n543), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n547), .B(new_n742), .C1(new_n592), .C2(new_n601), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n696), .A3(new_n744), .ZN(new_n745));
  OR3_X1    g559(.A1(new_n663), .A2(new_n306), .A3(KEYINPUT104), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT104), .B1(new_n663), .B2(new_n306), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n662), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n745), .A2(new_n748), .A3(new_n732), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n308), .A2(new_n373), .A3(new_n696), .A4(new_n743), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  INV_X1    g567(.A(new_n743), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n666), .A2(new_n610), .A3(new_n670), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  AOI21_X1  g570(.A(new_n493), .B1(new_n623), .B2(new_n622), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT43), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n613), .A2(KEYINPUT106), .A3(new_n653), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT106), .B1(new_n613), .B2(new_n653), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT44), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n548), .B1(new_n591), .B2(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n765), .A2(KEYINPUT105), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n586), .A2(KEYINPUT45), .A3(new_n590), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n765), .A2(KEYINPUT105), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(G469), .A2(G902), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n601), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n770), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n546), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n434), .A2(new_n439), .A3(new_n543), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT107), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n763), .A2(new_n775), .A3(new_n674), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  XNOR2_X1  g593(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n770), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT46), .B1(new_n769), .B2(new_n770), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n782), .A2(new_n783), .A3(new_n601), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(new_n784), .B2(new_n546), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n773), .A2(new_n774), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n547), .A3(new_n780), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n666), .A2(new_n610), .A3(new_n696), .A4(new_n776), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n785), .A2(new_n787), .A3(KEYINPUT109), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NAND2_X1  g608(.A1(new_n729), .A2(new_n734), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n758), .A2(new_n537), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n795), .A2(new_n363), .A3(new_n367), .A4(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n709), .A2(new_n543), .A3(new_n688), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n702), .A2(new_n547), .A3(new_n742), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n373), .A2(new_n802), .A3(new_n536), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n305), .A2(new_n307), .B1(G472), .B2(new_n681), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n805), .A2(new_n493), .A3(new_n624), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n796), .A2(new_n802), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n806), .B1(new_n738), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT116), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n785), .A2(new_n787), .ZN(new_n811));
  INV_X1    g625(.A(new_n702), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(new_n547), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n777), .A3(new_n797), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT51), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n748), .A2(new_n732), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n807), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n817), .B(KEYINPUT48), .Z(new_n818));
  NAND2_X1  g632(.A1(new_n797), .A2(new_n739), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n819), .B(new_n534), .C1(new_n625), .C2(new_n805), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n814), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n801), .A2(KEYINPUT51), .A3(new_n808), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n815), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n629), .A2(new_n691), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n653), .A2(new_n827), .A3(new_n668), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n607), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n826), .B1(new_n829), .B2(new_n804), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n619), .A2(new_n689), .A3(new_n690), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n685), .A2(new_n669), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n606), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n683), .A2(new_n833), .A3(KEYINPUT115), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n672), .A2(new_n698), .A3(new_n740), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT52), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n672), .A2(new_n740), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n830), .A2(new_n834), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n698), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n738), .A2(new_n697), .A3(new_n754), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n532), .A2(new_n668), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n637), .A2(new_n640), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT113), .B1(new_n742), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n637), .A2(new_n640), .A3(new_n845), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT113), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n776), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n606), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n666), .A2(new_n852), .A3(new_n653), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n755), .A2(new_n844), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n752), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n440), .A2(new_n544), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n720), .B(KEYINPUT112), .C1(new_n624), .C2(new_n689), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n625), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n856), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n607), .A2(new_n610), .A3(new_n614), .A4(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n658), .A2(new_n735), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n374), .B1(new_n603), .B2(new_n705), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n862), .A2(new_n711), .A3(new_n863), .A4(new_n722), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n843), .B1(new_n855), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n722), .A2(new_n711), .ZN(new_n866));
  AOI221_X4 g680(.A(new_n373), .B1(new_n704), .B2(new_n602), .C1(new_n677), .C2(new_n662), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n658), .A2(new_n735), .A3(new_n861), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT114), .A3(new_n752), .A4(new_n854), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n842), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n838), .A2(new_n839), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n865), .A2(new_n870), .ZN(new_n876));
  INV_X1    g690(.A(new_n842), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT53), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT54), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n872), .A2(KEYINPUT53), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n869), .A2(new_n752), .A3(new_n854), .ZN(new_n881));
  OR3_X1    g695(.A1(new_n880), .A2(new_n842), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n882), .B(new_n883), .C1(KEYINPUT53), .C2(new_n871), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n825), .A2(new_n885), .B1(G952), .B2(G953), .ZN(new_n886));
  AND4_X1   g700(.A1(new_n732), .A2(new_n547), .A3(new_n543), .A4(new_n757), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT110), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n688), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n888), .B2(new_n887), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n812), .A2(KEYINPUT49), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n812), .A2(KEYINPUT49), .ZN(new_n892));
  NOR4_X1   g706(.A1(new_n890), .A2(new_n683), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT111), .Z(new_n894));
  NAND2_X1  g708(.A1(new_n886), .A2(new_n894), .ZN(G75));
  NOR3_X1   g709(.A1(new_n880), .A2(new_n842), .A3(new_n881), .ZN(new_n896));
  OAI211_X1 g710(.A(G210), .B(G902), .C1(new_n878), .C2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n410), .A2(new_n422), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n421), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n423), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT55), .Z(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n903), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n897), .A2(new_n898), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n415), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n904), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT117), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n904), .A2(new_n911), .A3(new_n906), .A4(new_n908), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(G51));
  XOR2_X1   g727(.A(new_n770), .B(KEYINPUT57), .Z(new_n914));
  NOR2_X1   g728(.A1(new_n878), .A2(new_n896), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n883), .ZN(new_n916));
  INV_X1    g730(.A(new_n884), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n700), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n915), .A2(new_n265), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n769), .B(KEYINPUT118), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n907), .B1(new_n919), .B2(new_n922), .ZN(G54));
  NAND2_X1  g737(.A1(KEYINPUT58), .A2(G475), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n484), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  NOR4_X1   g740(.A1(new_n915), .A2(new_n265), .A3(new_n633), .A4(new_n924), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n907), .ZN(G60));
  OR2_X1    g742(.A1(new_n620), .A2(new_n621), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT119), .ZN(new_n930));
  XNOR2_X1  g744(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n931));
  NAND2_X1  g745(.A1(G478), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n930), .B(new_n933), .C1(new_n916), .C2(new_n917), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n908), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n930), .B1(new_n885), .B2(new_n933), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(G63));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT60), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n356), .B1(new_n915), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n882), .B1(KEYINPUT53), .B2(new_n871), .ZN(new_n941));
  INV_X1    g755(.A(new_n939), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n650), .A2(new_n651), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT121), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n941), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n940), .A2(new_n908), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT61), .B1(new_n946), .B2(KEYINPUT122), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n947), .B(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n540), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n415), .B1(new_n950), .B2(G224), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n864), .B2(new_n415), .ZN(new_n952));
  INV_X1    g766(.A(G898), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n900), .B1(new_n953), .B2(G953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n952), .B(new_n954), .ZN(G69));
  AND2_X1   g769(.A1(new_n455), .A2(new_n456), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n281), .B(new_n956), .Z(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n693), .ZN(new_n959));
  OAI21_X1  g773(.A(KEYINPUT62), .B1(new_n836), .B2(new_n959), .ZN(new_n960));
  OR3_X1    g774(.A1(new_n836), .A2(new_n959), .A3(KEYINPUT62), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n776), .B1(new_n857), .B2(new_n859), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n374), .A2(new_n607), .A3(new_n674), .A4(new_n962), .ZN(new_n963));
  AND4_X1   g777(.A1(new_n778), .A2(new_n960), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n793), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n958), .B1(new_n965), .B2(new_n415), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n775), .A2(new_n674), .A3(new_n816), .A4(new_n831), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n752), .A2(new_n755), .ZN(new_n968));
  INV_X1    g782(.A(new_n836), .ZN(new_n969));
  AND4_X1   g783(.A1(new_n778), .A2(new_n967), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n793), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n415), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n957), .B1(G900), .B2(G953), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n966), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(G953), .B1(new_n550), .B2(new_n667), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(new_n958), .B2(KEYINPUT123), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n974), .B(new_n977), .ZN(G72));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n793), .A2(new_n869), .A3(new_n970), .ZN(new_n980));
  XNOR2_X1  g794(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n981));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(KEYINPUT125), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n295), .A2(new_n260), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT126), .Z(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(KEYINPUT125), .B1(new_n980), .B2(new_n983), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n793), .A2(new_n964), .A3(new_n869), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n983), .ZN(new_n991));
  INV_X1    g805(.A(new_n678), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n678), .A2(new_n983), .A3(new_n985), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n875), .B2(new_n878), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n993), .A2(new_n908), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n979), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n980), .A2(new_n983), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT125), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n1000), .A2(new_n984), .A3(new_n986), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n995), .A2(new_n908), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1001), .A2(new_n1002), .A3(KEYINPUT127), .A4(new_n993), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n997), .A2(new_n1003), .ZN(G57));
endmodule


