//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n193), .B2(new_n187), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(G146), .B(new_n189), .C1(new_n193), .C2(new_n187), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G119), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT24), .B(G110), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n201), .A2(G128), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n202), .B(new_n206), .C1(new_n207), .C2(KEYINPUT23), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n205), .B1(G110), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n198), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT72), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n190), .A2(new_n192), .A3(new_n195), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n197), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n203), .A2(new_n204), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n208), .B2(G110), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  AND4_X1   g030(.A1(new_n211), .A2(new_n215), .A3(new_n197), .A4(new_n212), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n210), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G137), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT73), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT73), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n219), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n222), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n224), .A2(new_n227), .A3(KEYINPUT74), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT74), .B1(new_n224), .B2(new_n227), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n218), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n224), .A2(new_n227), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n231), .B(new_n210), .C1(new_n216), .C2(new_n217), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G217), .ZN(new_n234));
  INV_X1    g048(.A(G902), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(G234), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(G902), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n228), .A2(new_n229), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n215), .A2(new_n197), .A3(new_n212), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT72), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n213), .A2(new_n211), .A3(new_n215), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n241), .A2(new_n242), .B1(new_n198), .B2(new_n209), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n232), .B(new_n235), .C1(new_n239), .C2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n230), .A2(KEYINPUT25), .A3(new_n235), .A4(new_n232), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n246), .A2(KEYINPUT75), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT75), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n244), .A2(new_n249), .A3(new_n245), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n236), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n238), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT0), .A3(G128), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT64), .B1(new_n195), .B2(G143), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n255), .A3(G146), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT0), .B(G128), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n254), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n254), .B(new_n264), .C1(new_n260), .C2(new_n261), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT11), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(G137), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(G137), .ZN(new_n269));
  INV_X1    g083(.A(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT11), .A3(G134), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n268), .A2(new_n271), .A3(new_n274), .A4(new_n269), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n263), .A2(new_n265), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT67), .B1(new_n201), .B2(G116), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n279));
  INV_X1    g093(.A(G116), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(G119), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(KEYINPUT2), .A2(G113), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT2), .A2(G113), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n280), .A2(G119), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n282), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n285), .B1(new_n282), .B2(new_n287), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n195), .A2(G143), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n255), .A2(G146), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n199), .B1(new_n292), .B2(KEYINPUT1), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n260), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n269), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n267), .A2(G137), .ZN(new_n298));
  OAI21_X1  g112(.A(G131), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n275), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n277), .A2(new_n290), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G237), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n221), .A3(G210), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT27), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT26), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT27), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n303), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n305), .A2(new_n309), .A3(G101), .ZN(new_n310));
  AOI21_X1  g124(.A(G101), .B1(new_n305), .B2(new_n309), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n301), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n296), .A2(new_n275), .A3(new_n299), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n257), .A2(new_n259), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n261), .B1(new_n315), .B2(new_n292), .ZN(new_n316));
  AND4_X1   g130(.A1(KEYINPUT0), .A2(new_n292), .A3(new_n293), .A4(G128), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT65), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n254), .B(new_n319), .C1(new_n260), .C2(new_n261), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n276), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n314), .B1(new_n321), .B2(KEYINPUT66), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT66), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n318), .A2(new_n323), .A3(new_n276), .A4(new_n320), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT30), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n277), .A2(KEYINPUT30), .A3(new_n300), .ZN(new_n326));
  INV_X1    g140(.A(new_n290), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n313), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT31), .ZN(new_n330));
  INV_X1    g144(.A(G101), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n307), .A2(new_n308), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n304), .A2(KEYINPUT26), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n305), .A2(new_n309), .A3(G101), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n334), .A2(KEYINPUT69), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT69), .B1(new_n334), .B2(new_n335), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT28), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n301), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n277), .A2(KEYINPUT28), .A3(new_n290), .A4(new_n300), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n290), .B1(new_n322), .B2(new_n324), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n339), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT31), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n346), .B(new_n313), .C1(new_n325), .C2(new_n328), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n330), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT70), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT32), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT32), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n277), .A2(new_n300), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n327), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n341), .A2(new_n342), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n312), .A2(KEYINPUT29), .ZN(new_n360));
  OAI211_X1 g174(.A(KEYINPUT71), .B(new_n235), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n235), .B1(new_n359), .B2(new_n360), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT71), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n321), .A2(KEYINPUT66), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n300), .A3(new_n324), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n327), .A3(new_n326), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n312), .B1(new_n369), .B2(new_n301), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n366), .A2(new_n327), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n371), .A2(new_n338), .A3(new_n341), .A4(new_n342), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n361), .B(new_n364), .C1(new_n370), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G472), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n252), .B1(new_n356), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT9), .B(G234), .ZN(new_n378));
  OAI21_X1  g192(.A(G221), .B1(new_n378), .B2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT79), .B(G469), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(KEYINPUT76), .A2(G104), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(KEYINPUT76), .A2(G104), .ZN(new_n385));
  NOR2_X1   g199(.A1(KEYINPUT3), .A2(G107), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(KEYINPUT3), .A2(G107), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G101), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(KEYINPUT3), .A2(G107), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(G104), .B2(new_n386), .ZN(new_n396));
  OR2_X1    g210(.A1(KEYINPUT76), .A2(G104), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n391), .A3(new_n383), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n398), .A3(new_n331), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n401), .B(G101), .C1(new_n387), .C2(new_n393), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n263), .A2(new_n400), .A3(new_n265), .A4(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n397), .A2(new_n390), .A3(new_n383), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n331), .B1(G104), .B2(G107), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT10), .A3(new_n296), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n294), .B1(new_n295), .B2(new_n253), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n399), .A3(new_n406), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT10), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n411), .A2(KEYINPUT77), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT77), .B1(new_n411), .B2(new_n412), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n403), .B(new_n409), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n276), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n412), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT77), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n411), .A2(KEYINPUT77), .A3(new_n412), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n276), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n409), .A4(new_n403), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G140), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n221), .A2(G227), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(KEYINPUT80), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n296), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n407), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n422), .B1(new_n430), .B2(new_n411), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(KEYINPUT12), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n427), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n423), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n428), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n416), .B2(new_n423), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(KEYINPUT80), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n235), .B(new_n382), .C1(new_n438), .C2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n436), .B1(new_n435), .B2(new_n423), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n416), .A2(new_n423), .A3(new_n436), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G469), .B1(new_n444), .B2(G902), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n380), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G214), .B1(G237), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G210), .B1(G237), .B2(G902), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n450), .B(KEYINPUT88), .Z(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(KEYINPUT87), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n429), .A2(new_n191), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n262), .A2(G125), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n221), .A2(G224), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT84), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n459), .B(KEYINPUT83), .Z(new_n460));
  XNOR2_X1  g274(.A(new_n456), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT81), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT81), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n282), .A2(new_n287), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G113), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n469), .B2(new_n286), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n286), .B1(new_n278), .B2(new_n281), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n285), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n471), .A2(new_n473), .A3(new_n399), .A4(new_n406), .ZN(new_n474));
  XNOR2_X1  g288(.A(G110), .B(G122), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n399), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n402), .B1(new_n288), .B2(new_n289), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n474), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT6), .ZN(new_n479));
  INV_X1    g293(.A(new_n475), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n282), .A2(new_n287), .ZN(new_n481));
  INV_X1    g295(.A(new_n285), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n331), .B1(new_n396), .B2(new_n398), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n483), .A2(new_n473), .B1(new_n484), .B2(new_n401), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n467), .A2(new_n470), .B1(new_n285), .B2(new_n472), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n485), .A2(new_n400), .B1(new_n408), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n480), .B1(new_n487), .B2(KEYINPUT82), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n479), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n475), .B1(new_n489), .B2(new_n490), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(KEYINPUT82), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(KEYINPUT6), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n461), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n475), .B(KEYINPUT8), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n470), .B1(new_n481), .B2(new_n462), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n408), .A2(new_n473), .A3(new_n499), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n500), .A2(KEYINPUT85), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n408), .A2(new_n486), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(KEYINPUT85), .B2(new_n500), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n498), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n505), .A2(KEYINPUT86), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n454), .A2(new_n455), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n505), .B2(new_n459), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n459), .A2(new_n505), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n454), .A2(new_n455), .A3(new_n509), .A4(new_n506), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n478), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n235), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n453), .B1(new_n496), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n461), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n493), .A2(KEYINPUT6), .A3(new_n494), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n493), .A2(new_n494), .B1(KEYINPUT6), .B2(new_n478), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n501), .A2(new_n503), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n497), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n508), .A2(new_n478), .A3(new_n510), .ZN(new_n520));
  AOI21_X1  g334(.A(G902), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n453), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n449), .B1(new_n513), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n302), .A2(new_n221), .A3(G214), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n255), .ZN(new_n527));
  NOR2_X1   g341(.A1(G237), .A2(G953), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(G143), .A3(G214), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n274), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n196), .A3(new_n197), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n274), .A3(new_n529), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(new_n530), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n532), .A2(KEYINPUT92), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT92), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n531), .A2(new_n196), .A3(new_n538), .A4(new_n197), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n527), .A2(new_n529), .ZN(new_n540));
  NAND2_X1  g354(.A1(KEYINPUT18), .A2(G131), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT89), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n540), .A2(new_n545), .A3(new_n542), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n193), .A2(G146), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n212), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n540), .B2(new_n542), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n537), .A2(new_n539), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(G113), .B(G122), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n392), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n554), .B(KEYINPUT91), .Z(new_n555));
  INV_X1    g369(.A(new_n554), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT90), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n193), .B1(new_n557), .B2(KEYINPUT19), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT19), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(KEYINPUT90), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n193), .A2(KEYINPUT90), .A3(new_n559), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n195), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n534), .A2(new_n530), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n197), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n547), .A2(new_n551), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n552), .A2(new_n555), .B1(new_n556), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(G475), .A2(G902), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT20), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n532), .A2(KEYINPUT92), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n535), .A2(new_n536), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n573), .A3(new_n539), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n566), .A3(new_n555), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n567), .A2(new_n556), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT20), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n569), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n574), .A2(new_n566), .A3(new_n555), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n554), .B1(new_n574), .B2(new_n566), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n235), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n571), .A2(new_n579), .B1(G475), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n221), .A2(G952), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(G234), .B2(G237), .ZN(new_n585));
  NAND2_X1  g399(.A1(G234), .A2(G237), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(G902), .A3(G953), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT94), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT21), .B(G898), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n280), .A2(G122), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n390), .B1(new_n592), .B2(KEYINPUT14), .ZN(new_n593));
  XNOR2_X1  g407(.A(G116), .B(G122), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT14), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n593), .A2(new_n596), .B1(new_n390), .B2(new_n594), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n199), .A2(G143), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT93), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n255), .A2(G128), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n267), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n267), .B1(new_n599), .B2(new_n600), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n598), .B(KEYINPUT93), .Z(new_n605));
  INV_X1    g419(.A(KEYINPUT13), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n600), .B(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G134), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n594), .B(new_n390), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n601), .A3(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n378), .A2(new_n234), .A3(G953), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n604), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(new_n604), .B2(new_n610), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n235), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT15), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n615), .A3(G478), .ZN(new_n616));
  INV_X1    g430(.A(G478), .ZN(new_n617));
  OAI221_X1 g431(.A(new_n235), .B1(KEYINPUT15), .B2(new_n617), .C1(new_n612), .C2(new_n613), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n583), .A2(new_n591), .A3(new_n620), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n447), .A2(new_n525), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n377), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  INV_X1    g438(.A(G472), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n348), .B2(new_n235), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n348), .B2(new_n349), .ZN(new_n627));
  INV_X1    g441(.A(new_n252), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n627), .A2(new_n628), .A3(new_n446), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n517), .A2(new_n451), .A3(new_n521), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n452), .B1(new_n496), .B2(new_n512), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n631), .A3(new_n448), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n582), .A2(G475), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n578), .B1(new_n577), .B2(new_n569), .ZN(new_n634));
  AOI211_X1 g448(.A(KEYINPUT20), .B(new_n570), .C1(new_n575), .C2(new_n576), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n613), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n604), .A2(new_n610), .A3(new_n611), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n639));
  NAND3_X1  g453(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  OAI22_X1  g455(.A1(new_n612), .A2(new_n613), .B1(KEYINPUT95), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n640), .A2(new_n642), .A3(G478), .A4(new_n235), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n614), .A2(new_n617), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n636), .A2(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n632), .A2(new_n646), .A3(new_n590), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n629), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  INV_X1    g464(.A(KEYINPUT96), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n633), .B(new_n619), .C1(new_n634), .C2(new_n635), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n651), .B1(new_n653), .B2(new_n591), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n652), .A2(KEYINPUT96), .A3(new_n590), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n654), .A2(new_n632), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n629), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NOR3_X1   g473(.A1(new_n228), .A2(new_n229), .A3(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n218), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n237), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(new_n248), .B2(new_n251), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n246), .A2(KEYINPUT75), .A3(new_n247), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n236), .A3(new_n250), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(KEYINPUT97), .A3(new_n662), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n621), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n669), .A2(new_n627), .A3(new_n446), .A4(new_n524), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT37), .B(G110), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT98), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n672), .B(KEYINPUT99), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n670), .B(new_n673), .ZN(G12));
  NAND2_X1  g488(.A1(new_n665), .A2(new_n668), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n675), .A2(new_n446), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT32), .B1(new_n350), .B2(new_n351), .ZN(new_n677));
  AOI211_X1 g491(.A(KEYINPUT70), .B(new_n353), .C1(new_n348), .C2(new_n349), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n376), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n585), .B1(new_n588), .B2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n632), .A2(new_n652), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT100), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n199), .ZN(G30));
  XOR2_X1   g500(.A(new_n682), .B(KEYINPUT39), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n446), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT40), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n689), .A2(KEYINPUT101), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(KEYINPUT101), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n338), .B1(new_n301), .B2(new_n358), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n369), .B2(new_n313), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n356), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n513), .A2(new_n523), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT38), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n513), .A2(new_n523), .A3(KEYINPUT38), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n583), .A2(new_n620), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n448), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n696), .A2(new_n675), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n690), .A2(new_n691), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT102), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n255), .ZN(G45));
  NOR3_X1   g521(.A1(new_n632), .A2(new_n646), .A3(new_n682), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n680), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  INV_X1    g524(.A(new_n377), .ZN(new_n711));
  INV_X1    g525(.A(new_n415), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n427), .B1(new_n712), .B2(new_n422), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n439), .A2(KEYINPUT80), .B1(new_n713), .B2(new_n435), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n424), .A2(new_n427), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT80), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(G902), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(G469), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n441), .B(new_n379), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n711), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n647), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND2_X1  g538(.A1(new_n721), .A2(new_n656), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND2_X1  g540(.A1(new_n714), .A2(new_n717), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n719), .B1(new_n727), .B2(new_n235), .ZN(new_n728));
  AOI211_X1 g542(.A(G902), .B(new_n381), .C1(new_n714), .C2(new_n717), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n632), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(KEYINPUT103), .A3(new_n379), .A4(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT103), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n720), .B2(new_n632), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n679), .A2(new_n669), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  INV_X1    g552(.A(new_n720), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n339), .A2(new_n359), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n330), .A2(new_n347), .A3(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(new_n349), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n742), .A2(new_n626), .A3(new_n252), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n583), .A2(new_n590), .A3(new_n620), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n739), .A2(new_n731), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  NOR2_X1   g560(.A1(new_n742), .A2(new_n626), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n675), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n646), .A2(new_n682), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n735), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  NAND2_X1  g567(.A1(new_n350), .A2(new_n353), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n348), .A2(KEYINPUT32), .A3(new_n349), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n376), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n628), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n513), .A2(new_n523), .A3(new_n448), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n446), .A2(new_n749), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT42), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n441), .A2(new_n445), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n761), .A2(new_n379), .A3(new_n758), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n646), .A2(KEYINPUT42), .A3(new_n682), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n679), .A3(new_n628), .A4(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  INV_X1    g580(.A(KEYINPUT104), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n652), .A2(new_n682), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n377), .A2(new_n767), .A3(new_n768), .A4(new_n762), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n762), .A2(new_n679), .A3(new_n628), .A4(new_n768), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT104), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  OAI211_X1 g587(.A(new_n583), .B(new_n645), .C1(KEYINPUT106), .C2(KEYINPUT43), .ZN(new_n774));
  INV_X1    g588(.A(new_n645), .ZN(new_n775));
  AND2_X1   g589(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n776));
  NOR2_X1   g590(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n777));
  OAI22_X1  g591(.A1(new_n636), .A2(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n675), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(new_n627), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n444), .A2(KEYINPUT45), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n442), .B2(new_n443), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(G469), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(G469), .A2(G902), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT46), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n729), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n788), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT105), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(new_n379), .ZN(new_n796));
  INV_X1    g610(.A(new_n758), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n781), .B2(new_n782), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n783), .A2(new_n796), .A3(new_n798), .A4(new_n687), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  AND2_X1   g614(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n795), .A2(new_n379), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n795), .B2(new_n379), .ZN(new_n806));
  OR4_X1    g620(.A1(new_n679), .A2(new_n750), .A3(new_n628), .A4(new_n797), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n803), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT108), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n188), .ZN(G42));
  AOI22_X1  g624(.A1(new_n735), .A2(new_n736), .B1(new_n377), .B2(new_n622), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n652), .B1(new_n583), .B2(new_n775), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n812), .A2(new_n524), .A3(new_n591), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(new_n628), .A3(new_n627), .A4(new_n446), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n814), .A2(new_n745), .A3(new_n670), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n377), .B(new_n739), .C1(new_n647), .C2(new_n656), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n811), .A2(new_n765), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n676), .B(new_n679), .C1(new_n683), .C2(new_n708), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n448), .A2(new_n702), .A3(new_n631), .A4(new_n630), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n663), .A2(new_n682), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n695), .A2(new_n446), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n752), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n752), .A2(new_n818), .A3(KEYINPUT52), .A4(new_n821), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n817), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n675), .A2(new_n446), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n827), .A2(new_n682), .A3(new_n797), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n679), .A2(new_n620), .A3(new_n583), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n646), .A2(new_n742), .A3(new_n626), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n770), .A2(KEYINPUT104), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n770), .A2(KEYINPUT104), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT110), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT110), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n772), .A2(new_n836), .A3(new_n831), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT53), .B1(new_n826), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n826), .A2(new_n838), .ZN(new_n841));
  XOR2_X1   g655(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n842));
  OAI22_X1  g656(.A1(new_n839), .A2(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n824), .A2(new_n825), .ZN(new_n845));
  INV_X1    g659(.A(new_n817), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n772), .A2(new_n836), .A3(new_n831), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n836), .B1(new_n772), .B2(new_n831), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n844), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(KEYINPUT111), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT54), .B1(new_n843), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n696), .A2(new_n628), .ZN(new_n854));
  INV_X1    g668(.A(new_n585), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n720), .A2(new_n797), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n646), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n584), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n743), .A2(new_n779), .A3(new_n585), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n735), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n861), .B1(new_n735), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n860), .B(KEYINPUT118), .C1(new_n863), .C2(new_n864), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT119), .Z(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n856), .A2(new_n779), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n872), .B1(new_n873), .B2(new_n757), .ZN(new_n874));
  NAND2_X1  g688(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n875));
  INV_X1    g689(.A(new_n757), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n856), .A3(new_n779), .A4(new_n871), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n730), .ZN(new_n879));
  OAI22_X1  g693(.A1(new_n803), .A2(new_n806), .B1(new_n379), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n758), .A3(new_n862), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n636), .A2(new_n645), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n696), .A2(new_n628), .A3(new_n856), .A4(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n883), .B(KEYINPUT51), .C1(new_n748), .C2(new_n873), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n862), .A2(new_n449), .A3(new_n701), .A4(new_n739), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT114), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT50), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT50), .B1(new_n885), .B2(new_n886), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n884), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n878), .B1(new_n881), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n869), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT115), .B1(new_n888), .B2(new_n889), .ZN(new_n893));
  INV_X1    g707(.A(new_n889), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT115), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n895), .A3(new_n887), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n873), .A2(new_n748), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n858), .B2(new_n882), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n893), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT116), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT116), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n893), .A2(new_n896), .A3(new_n901), .A4(new_n898), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n902), .A3(new_n881), .ZN(new_n903));
  XNOR2_X1  g717(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n892), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n826), .A2(new_n838), .A3(KEYINPUT53), .ZN(new_n906));
  INV_X1    g720(.A(new_n842), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n826), .B2(new_n838), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n908), .A3(KEYINPUT54), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n853), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(G952), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n221), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n583), .A2(new_n379), .A3(new_n448), .A4(new_n645), .ZN(new_n915));
  INV_X1    g729(.A(new_n701), .ZN(new_n916));
  AOI211_X1 g730(.A(new_n915), .B(new_n916), .C1(KEYINPUT49), .C2(new_n879), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(KEYINPUT49), .B2(new_n879), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n854), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT109), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n914), .A2(new_n920), .ZN(G75));
  NAND2_X1  g735(.A1(new_n912), .A2(G953), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT123), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n842), .B1(new_n847), .B2(new_n850), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n826), .A2(new_n838), .A3(KEYINPUT53), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n235), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT56), .B1(new_n926), .B2(new_n451), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n515), .A2(new_n516), .A3(new_n514), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(new_n496), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT55), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n923), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(G902), .B1(new_n906), .B2(new_n908), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT121), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n934), .B(G902), .C1(new_n906), .C2(new_n908), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n451), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT122), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(KEYINPUT56), .ZN(new_n938));
  MUX2_X1   g752(.A(new_n937), .B(new_n938), .S(new_n930), .Z(new_n939));
  AOI21_X1  g753(.A(new_n931), .B1(new_n936), .B2(new_n939), .ZN(G51));
  INV_X1    g754(.A(new_n923), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n788), .B(KEYINPUT57), .Z(new_n942));
  INV_X1    g756(.A(KEYINPUT54), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n924), .B2(new_n925), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n909), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n727), .B(KEYINPUT124), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n787), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n933), .A2(new_n948), .A3(new_n935), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n941), .B1(new_n947), .B2(new_n949), .ZN(G54));
  AND2_X1   g764(.A1(KEYINPUT58), .A2(G475), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n933), .A2(new_n935), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n577), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n933), .A2(new_n568), .A3(new_n935), .A4(new_n951), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n941), .B1(new_n953), .B2(new_n954), .ZN(G60));
  NAND2_X1  g769(.A1(new_n640), .A2(new_n642), .ZN(new_n956));
  NAND2_X1  g770(.A1(G478), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT59), .Z(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n909), .B2(new_n944), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n923), .ZN(new_n961));
  INV_X1    g775(.A(new_n958), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n847), .A2(new_n850), .ZN(new_n963));
  AOI22_X1  g777(.A1(new_n851), .A2(KEYINPUT111), .B1(new_n963), .B2(new_n907), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n839), .A2(new_n840), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n943), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n962), .B1(new_n966), .B2(new_n909), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n961), .B1(new_n967), .B2(new_n956), .ZN(G63));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT60), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n924), .B2(new_n925), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n661), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n233), .B(KEYINPUT125), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n923), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n969), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n972), .A2(new_n975), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n978), .A2(KEYINPUT61), .A3(new_n923), .A4(new_n973), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(G66));
  INV_X1    g794(.A(G224), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n589), .A2(new_n981), .A3(new_n221), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n811), .A2(new_n815), .A3(new_n816), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n982), .B1(new_n984), .B2(new_n221), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT126), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n492), .B(new_n495), .C1(G898), .C2(new_n221), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G69));
  NAND2_X1  g802(.A1(new_n368), .A2(new_n326), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n561), .A2(new_n562), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT127), .Z(new_n991));
  XNOR2_X1  g805(.A(new_n989), .B(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n808), .A2(new_n772), .A3(new_n799), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n796), .A2(new_n687), .A3(new_n876), .A4(new_n819), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n752), .A2(new_n818), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n994), .A2(new_n765), .A3(new_n995), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n993), .A2(G953), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n681), .A2(new_n221), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n992), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n705), .A2(new_n995), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n758), .A2(new_n812), .ZN(new_n1002));
  OR3_X1    g816(.A1(new_n711), .A2(new_n688), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n808), .A2(new_n799), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT62), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n705), .B2(new_n995), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n1001), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n992), .A2(G953), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n999), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(G227), .ZN(new_n1010));
  OAI21_X1  g824(.A(G953), .B1(new_n1010), .B2(new_n681), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1009), .B(new_n1011), .ZN(G72));
  AND2_X1   g826(.A1(new_n369), .A2(new_n301), .ZN(new_n1013));
  INV_X1    g827(.A(new_n312), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n993), .A2(new_n983), .A3(new_n996), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1016), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1020), .B1(new_n1007), .B2(new_n984), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n923), .B(new_n1021), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n964), .A2(new_n965), .ZN(new_n1026));
  NOR3_X1   g840(.A1(new_n1016), .A2(new_n1023), .A3(new_n1020), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(G57));
endmodule


