

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735;

  NOR2_X1 U366 ( .A1(n682), .A2(n681), .ZN(n585) );
  INV_X1 U367 ( .A(G953), .ZN(n715) );
  XNOR2_X2 U368 ( .A(n515), .B(n514), .ZN(n537) );
  AND2_X2 U369 ( .A1(n345), .A2(n548), .ZN(n515) );
  XNOR2_X2 U370 ( .A(n558), .B(n557), .ZN(n706) );
  XNOR2_X2 U371 ( .A(n465), .B(n464), .ZN(n510) );
  XNOR2_X2 U372 ( .A(n444), .B(n379), .ZN(n721) );
  XNOR2_X2 U373 ( .A(n479), .B(KEYINPUT4), .ZN(n444) );
  AND2_X1 U374 ( .A1(n385), .A2(n603), .ZN(n384) );
  XNOR2_X2 U375 ( .A(n434), .B(n713), .ZN(n445) );
  XNOR2_X1 U376 ( .A(n540), .B(KEYINPUT32), .ZN(n734) );
  NAND2_X1 U377 ( .A1(n539), .A2(n538), .ZN(n540) );
  AND2_X1 U378 ( .A1(n497), .A2(n549), .ZN(n528) );
  XNOR2_X1 U379 ( .A(n470), .B(G134), .ZN(n379) );
  NOR2_X2 U380 ( .A1(n626), .A2(n705), .ZN(n627) );
  OR2_X1 U381 ( .A1(n683), .A2(KEYINPUT47), .ZN(n559) );
  NOR2_X1 U382 ( .A1(n525), .A2(n526), .ZN(n583) );
  NOR2_X1 U383 ( .A1(n581), .A2(n658), .ZN(n582) );
  XNOR2_X1 U384 ( .A(G113), .B(KEYINPUT5), .ZN(n380) );
  XNOR2_X1 U385 ( .A(G137), .B(G119), .ZN(n417) );
  NOR2_X1 U386 ( .A1(n733), .A2(n542), .ZN(n544) );
  XNOR2_X1 U387 ( .A(G146), .B(G125), .ZN(n446) );
  AND2_X1 U388 ( .A1(n655), .A2(n652), .ZN(n683) );
  NAND2_X1 U389 ( .A1(n623), .A2(n460), .ZN(n424) );
  XNOR2_X1 U390 ( .A(G110), .B(G107), .ZN(n427) );
  XOR2_X1 U391 ( .A(KEYINPUT78), .B(G104), .Z(n428) );
  XNOR2_X1 U392 ( .A(n430), .B(n429), .ZN(n431) );
  INV_X1 U393 ( .A(KEYINPUT94), .ZN(n429) );
  INV_X1 U394 ( .A(KEYINPUT67), .ZN(n423) );
  XNOR2_X1 U395 ( .A(G137), .B(G140), .ZN(n433) );
  NAND2_X1 U396 ( .A1(n372), .A2(KEYINPUT2), .ZN(n370) );
  XNOR2_X1 U397 ( .A(n389), .B(KEYINPUT105), .ZN(n388) );
  NAND2_X1 U398 ( .A1(n574), .A2(n573), .ZN(n389) );
  XNOR2_X1 U399 ( .A(n378), .B(n377), .ZN(n376) );
  INV_X1 U400 ( .A(KEYINPUT34), .ZN(n377) );
  INV_X1 U401 ( .A(KEYINPUT22), .ZN(n514) );
  AND2_X1 U402 ( .A1(n443), .A2(n442), .ZN(n586) );
  NAND2_X1 U403 ( .A1(n361), .A2(n358), .ZN(n500) );
  NAND2_X1 U404 ( .A1(n360), .A2(n359), .ZN(n358) );
  NOR2_X1 U405 ( .A1(n362), .A2(n346), .ZN(n361) );
  INV_X1 U406 ( .A(n500), .ZN(n526) );
  XNOR2_X1 U407 ( .A(n671), .B(KEYINPUT6), .ZN(n574) );
  AND2_X1 U408 ( .A1(n612), .A2(G953), .ZN(n705) );
  XNOR2_X1 U409 ( .A(n398), .B(KEYINPUT21), .ZN(n399) );
  NAND2_X1 U410 ( .A1(n660), .A2(KEYINPUT88), .ZN(n385) );
  NAND2_X1 U411 ( .A1(n551), .A2(n354), .ZN(n553) );
  XNOR2_X1 U412 ( .A(n455), .B(n454), .ZN(n481) );
  INV_X1 U413 ( .A(G122), .ZN(n454) );
  XNOR2_X1 U414 ( .A(G116), .B(G107), .ZN(n455) );
  NAND2_X1 U415 ( .A1(G234), .A2(G237), .ZN(n390) );
  XNOR2_X1 U416 ( .A(n415), .B(n414), .ZN(n493) );
  XNOR2_X1 U417 ( .A(G475), .B(KEYINPUT13), .ZN(n363) );
  AND2_X1 U418 ( .A1(n617), .A2(n363), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n438), .B(n381), .ZN(n623) );
  XOR2_X1 U420 ( .A(G119), .B(G110), .Z(n456) );
  XOR2_X1 U421 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n406) );
  XNOR2_X1 U422 ( .A(KEYINPUT69), .B(KEYINPUT10), .ZN(n409) );
  XNOR2_X1 U423 ( .A(n467), .B(n357), .ZN(n356) );
  INV_X1 U424 ( .A(KEYINPUT11), .ZN(n357) );
  XNOR2_X1 U425 ( .A(G140), .B(KEYINPUT99), .ZN(n467) );
  XNOR2_X1 U426 ( .A(KEYINPUT100), .B(KEYINPUT12), .ZN(n355) );
  XNOR2_X1 U427 ( .A(G143), .B(G122), .ZN(n469) );
  XNOR2_X1 U428 ( .A(n532), .B(KEYINPUT33), .ZN(n677) );
  XNOR2_X1 U429 ( .A(n672), .B(n530), .ZN(n531) );
  INV_X1 U430 ( .A(KEYINPUT41), .ZN(n584) );
  BUF_X1 U431 ( .A(n517), .Z(n545) );
  NAND2_X1 U432 ( .A1(n369), .A2(n494), .ZN(n672) );
  XNOR2_X1 U433 ( .A(n496), .B(n495), .ZN(n549) );
  XNOR2_X1 U434 ( .A(n438), .B(n437), .ZN(n636) );
  AND2_X1 U435 ( .A1(n580), .A2(n369), .ZN(n658) );
  XNOR2_X1 U436 ( .A(n374), .B(n351), .ZN(n733) );
  INV_X1 U437 ( .A(n533), .ZN(n375) );
  NAND2_X1 U438 ( .A1(n586), .A2(n466), .ZN(n648) );
  NAND2_X1 U439 ( .A1(n526), .A2(n486), .ZN(n652) );
  NAND2_X1 U440 ( .A1(n701), .A2(G217), .ZN(n630) );
  OR2_X1 U441 ( .A1(G902), .A2(n703), .ZN(n343) );
  XOR2_X1 U442 ( .A(n356), .B(n355), .Z(n344) );
  XNOR2_X1 U443 ( .A(KEYINPUT101), .B(n513), .ZN(n345) );
  NAND2_X1 U444 ( .A1(n493), .A2(n512), .ZN(n666) );
  AND2_X1 U445 ( .A1(n363), .A2(G902), .ZN(n346) );
  AND2_X1 U446 ( .A1(n576), .A2(n577), .ZN(n347) );
  AND2_X1 U447 ( .A1(n388), .A2(n576), .ZN(n348) );
  AND2_X1 U448 ( .A1(n600), .A2(n602), .ZN(n349) );
  XOR2_X1 U449 ( .A(KEYINPUT65), .B(KEYINPUT1), .Z(n350) );
  XOR2_X1 U450 ( .A(KEYINPUT87), .B(KEYINPUT35), .Z(n351) );
  AND2_X1 U451 ( .A1(n373), .A2(n365), .ZN(n352) );
  INV_X1 U452 ( .A(n604), .ZN(n373) );
  XNOR2_X1 U453 ( .A(G902), .B(KEYINPUT15), .ZN(n604) );
  NAND2_X1 U454 ( .A1(n353), .A2(n373), .ZN(n364) );
  INV_X1 U455 ( .A(n605), .ZN(n353) );
  NAND2_X2 U456 ( .A1(n706), .A2(n724), .ZN(n605) );
  XNOR2_X2 U457 ( .A(n511), .B(KEYINPUT0), .ZN(n548) );
  NAND2_X1 U458 ( .A1(n368), .A2(n367), .ZN(n371) );
  AND2_X2 U459 ( .A1(n371), .A2(n370), .ZN(n629) );
  INV_X1 U460 ( .A(n683), .ZN(n354) );
  NOR2_X1 U461 ( .A1(n363), .A2(G902), .ZN(n359) );
  INV_X1 U462 ( .A(n617), .ZN(n360) );
  NAND2_X1 U463 ( .A1(n364), .A2(KEYINPUT85), .ZN(n367) );
  INV_X1 U464 ( .A(n605), .ZN(n372) );
  NAND2_X1 U465 ( .A1(n605), .A2(n692), .ZN(n366) );
  NAND2_X1 U466 ( .A1(n366), .A2(n352), .ZN(n368) );
  NAND2_X1 U467 ( .A1(KEYINPUT85), .A2(n692), .ZN(n365) );
  XNOR2_X2 U468 ( .A(KEYINPUT3), .B(KEYINPUT73), .ZN(n713) );
  XNOR2_X2 U469 ( .A(n516), .B(n350), .ZN(n369) );
  XNOR2_X2 U470 ( .A(n440), .B(n439), .ZN(n516) );
  INV_X1 U471 ( .A(n369), .ZN(n529) );
  NAND2_X1 U472 ( .A1(n376), .A2(n375), .ZN(n374) );
  NAND2_X1 U473 ( .A1(n677), .A2(n548), .ZN(n378) );
  XNOR2_X2 U474 ( .A(n721), .B(G146), .ZN(n438) );
  XNOR2_X1 U475 ( .A(n380), .B(G116), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n382), .B(n422), .ZN(n381) );
  XNOR2_X1 U477 ( .A(n445), .B(n421), .ZN(n382) );
  NOR2_X2 U478 ( .A1(n387), .A2(n383), .ZN(n724) );
  NAND2_X1 U479 ( .A1(n386), .A2(n384), .ZN(n383) );
  NAND2_X1 U480 ( .A1(n601), .A2(n349), .ZN(n386) );
  NOR2_X1 U481 ( .A1(n601), .A2(n602), .ZN(n387) );
  NAND2_X1 U482 ( .A1(n388), .A2(n347), .ZN(n579) );
  NAND2_X1 U483 ( .A1(n528), .A2(n527), .ZN(n565) );
  AND2_X1 U484 ( .A1(n492), .A2(n491), .ZN(n497) );
  INV_X1 U485 ( .A(KEYINPUT104), .ZN(n530) );
  INV_X1 U486 ( .A(KEYINPUT44), .ZN(n543) );
  XNOR2_X1 U487 ( .A(n400), .B(n399), .ZN(n661) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n436) );
  INV_X1 U489 ( .A(n598), .ZN(n577) );
  XNOR2_X1 U490 ( .A(n598), .B(KEYINPUT38), .ZN(n679) );
  XNOR2_X1 U491 ( .A(n585), .B(n584), .ZN(n693) );
  XNOR2_X1 U492 ( .A(n390), .B(KEYINPUT14), .ZN(n391) );
  XNOR2_X1 U493 ( .A(KEYINPUT76), .B(n391), .ZN(n393) );
  NAND2_X1 U494 ( .A1(n393), .A2(G952), .ZN(n392) );
  XOR2_X1 U495 ( .A(KEYINPUT93), .B(n392), .Z(n691) );
  NOR2_X1 U496 ( .A1(G953), .A2(n691), .ZN(n508) );
  AND2_X1 U497 ( .A1(n393), .A2(G953), .ZN(n394) );
  NAND2_X1 U498 ( .A1(G902), .A2(n394), .ZN(n506) );
  NOR2_X1 U499 ( .A1(G900), .A2(n506), .ZN(n395) );
  OR2_X1 U500 ( .A1(n508), .A2(n395), .ZN(n396) );
  XNOR2_X1 U501 ( .A(n396), .B(KEYINPUT80), .ZN(n491) );
  NAND2_X1 U502 ( .A1(n604), .A2(G234), .ZN(n397) );
  XNOR2_X1 U503 ( .A(n397), .B(KEYINPUT20), .ZN(n412) );
  NAND2_X1 U504 ( .A1(n412), .A2(G221), .ZN(n400) );
  XOR2_X1 U505 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n398) );
  INV_X1 U506 ( .A(n661), .ZN(n401) );
  AND2_X1 U507 ( .A1(n491), .A2(n401), .ZN(n416) );
  XNOR2_X1 U508 ( .A(G128), .B(KEYINPUT24), .ZN(n403) );
  XNOR2_X1 U509 ( .A(KEYINPUT84), .B(KEYINPUT23), .ZN(n402) );
  XNOR2_X1 U510 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U511 ( .A(n456), .B(n404), .ZN(n408) );
  NAND2_X1 U512 ( .A1(G234), .A2(n715), .ZN(n405) );
  XNOR2_X1 U513 ( .A(n406), .B(n405), .ZN(n478) );
  NAND2_X1 U514 ( .A1(n478), .A2(G221), .ZN(n407) );
  XNOR2_X1 U515 ( .A(n408), .B(n407), .ZN(n411) );
  XNOR2_X1 U516 ( .A(n446), .B(n409), .ZN(n474) );
  INV_X1 U517 ( .A(n433), .ZN(n410) );
  XNOR2_X1 U518 ( .A(n474), .B(n410), .ZN(n723) );
  XNOR2_X1 U519 ( .A(n411), .B(n723), .ZN(n631) );
  INV_X1 U520 ( .A(G902), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n631), .A2(n460), .ZN(n415) );
  AND2_X1 U522 ( .A1(n412), .A2(G217), .ZN(n413) );
  XNOR2_X1 U523 ( .A(n413), .B(KEYINPUT25), .ZN(n414) );
  INV_X1 U524 ( .A(n493), .ZN(n521) );
  AND2_X1 U525 ( .A1(n416), .A2(n521), .ZN(n573) );
  XNOR2_X1 U526 ( .A(n418), .B(n417), .ZN(n422) );
  INV_X1 U527 ( .A(G953), .ZN(n448) );
  INV_X1 U528 ( .A(G237), .ZN(n419) );
  NAND2_X1 U529 ( .A1(n448), .A2(n419), .ZN(n420) );
  XNOR2_X1 U530 ( .A(KEYINPUT77), .B(n420), .ZN(n468) );
  NAND2_X1 U531 ( .A1(n468), .A2(G210), .ZN(n421) );
  XNOR2_X2 U532 ( .A(n423), .B(G101), .ZN(n434) );
  XNOR2_X2 U533 ( .A(G143), .B(G128), .ZN(n479) );
  XNOR2_X2 U534 ( .A(KEYINPUT70), .B(G131), .ZN(n470) );
  XNOR2_X2 U535 ( .A(n424), .B(G472), .ZN(n517) );
  NAND2_X1 U536 ( .A1(n573), .A2(n545), .ZN(n426) );
  INV_X1 U537 ( .A(KEYINPUT28), .ZN(n425) );
  XNOR2_X1 U538 ( .A(n426), .B(n425), .ZN(n443) );
  XNOR2_X1 U539 ( .A(n428), .B(n427), .ZN(n432) );
  NAND2_X1 U540 ( .A1(G227), .A2(n715), .ZN(n430) );
  XNOR2_X1 U541 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U542 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U543 ( .A1(n636), .A2(n460), .ZN(n440) );
  XNOR2_X1 U544 ( .A(KEYINPUT72), .B(G469), .ZN(n439) );
  INV_X1 U545 ( .A(KEYINPUT107), .ZN(n441) );
  XNOR2_X1 U546 ( .A(n516), .B(n441), .ZN(n442) );
  XNOR2_X1 U547 ( .A(n445), .B(n444), .ZN(n453) );
  XNOR2_X1 U548 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n447) );
  XNOR2_X1 U549 ( .A(n447), .B(n446), .ZN(n451) );
  NAND2_X1 U550 ( .A1(G224), .A2(n448), .ZN(n449) );
  XNOR2_X1 U551 ( .A(n449), .B(KEYINPUT79), .ZN(n450) );
  XNOR2_X1 U552 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U553 ( .A(n453), .B(n452), .ZN(n459) );
  XOR2_X1 U554 ( .A(G113), .B(G104), .Z(n475) );
  XNOR2_X1 U555 ( .A(n481), .B(n475), .ZN(n458) );
  XNOR2_X1 U556 ( .A(KEYINPUT16), .B(n456), .ZN(n457) );
  XNOR2_X1 U557 ( .A(n458), .B(n457), .ZN(n711) );
  XNOR2_X1 U558 ( .A(n711), .B(n459), .ZN(n606) );
  NAND2_X1 U559 ( .A1(n606), .A2(n604), .ZN(n462) );
  NAND2_X1 U560 ( .A1(n460), .A2(n419), .ZN(n463) );
  NAND2_X1 U561 ( .A1(n463), .A2(G210), .ZN(n461) );
  XNOR2_X2 U562 ( .A(n462), .B(n461), .ZN(n598) );
  NAND2_X1 U563 ( .A1(n463), .A2(G214), .ZN(n678) );
  NAND2_X1 U564 ( .A1(n577), .A2(n678), .ZN(n465) );
  INV_X1 U565 ( .A(KEYINPUT19), .ZN(n464) );
  INV_X1 U566 ( .A(n510), .ZN(n466) );
  NAND2_X1 U567 ( .A1(n468), .A2(G214), .ZN(n472) );
  XNOR2_X1 U568 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U569 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U570 ( .A(n344), .B(n473), .ZN(n477) );
  XNOR2_X1 U571 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U572 ( .A(n477), .B(n476), .ZN(n617) );
  XNOR2_X1 U573 ( .A(G134), .B(KEYINPUT9), .ZN(n485) );
  NAND2_X1 U574 ( .A1(G217), .A2(n478), .ZN(n483) );
  XOR2_X1 U575 ( .A(KEYINPUT7), .B(n479), .Z(n480) );
  XNOR2_X1 U576 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U577 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U578 ( .A(n485), .B(n484), .ZN(n703) );
  XNOR2_X2 U579 ( .A(G478), .B(n343), .ZN(n525) );
  INV_X1 U580 ( .A(n525), .ZN(n486) );
  NOR2_X1 U581 ( .A1(n648), .A2(n652), .ZN(n487) );
  XOR2_X1 U582 ( .A(G146), .B(n487), .Z(G48) );
  NAND2_X1 U583 ( .A1(n517), .A2(n678), .ZN(n490) );
  INV_X1 U584 ( .A(KEYINPUT106), .ZN(n488) );
  XNOR2_X1 U585 ( .A(n488), .B(KEYINPUT30), .ZN(n489) );
  XNOR2_X1 U586 ( .A(n490), .B(n489), .ZN(n492) );
  XNOR2_X1 U587 ( .A(n661), .B(KEYINPUT97), .ZN(n512) );
  INV_X1 U588 ( .A(n666), .ZN(n494) );
  NAND2_X1 U589 ( .A1(n516), .A2(n494), .ZN(n496) );
  INV_X1 U590 ( .A(KEYINPUT98), .ZN(n495) );
  NAND2_X1 U591 ( .A1(n528), .A2(n679), .ZN(n499) );
  INV_X1 U592 ( .A(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U593 ( .A(n499), .B(n498), .ZN(n501) );
  NAND2_X1 U594 ( .A1(n500), .A2(n525), .ZN(n655) );
  OR2_X1 U595 ( .A1(n501), .A2(n655), .ZN(n603) );
  XNOR2_X1 U596 ( .A(n603), .B(G134), .ZN(G36) );
  INV_X1 U597 ( .A(n501), .ZN(n503) );
  INV_X1 U598 ( .A(n652), .ZN(n502) );
  NAND2_X1 U599 ( .A1(n503), .A2(n502), .ZN(n505) );
  XNOR2_X1 U600 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n504) );
  XNOR2_X1 U601 ( .A(n505), .B(n504), .ZN(n590) );
  XNOR2_X1 U602 ( .A(n590), .B(G131), .ZN(G33) );
  NOR2_X1 U603 ( .A1(G898), .A2(n506), .ZN(n507) );
  NOR2_X1 U604 ( .A1(n508), .A2(n507), .ZN(n509) );
  NOR2_X2 U605 ( .A1(n510), .A2(n509), .ZN(n511) );
  NAND2_X1 U606 ( .A1(n512), .A2(n583), .ZN(n513) );
  INV_X1 U607 ( .A(n537), .ZN(n524) );
  INV_X1 U608 ( .A(n517), .ZN(n671) );
  NAND2_X1 U609 ( .A1(n671), .A2(n521), .ZN(n518) );
  NOR2_X1 U610 ( .A1(n369), .A2(n518), .ZN(n519) );
  NAND2_X1 U611 ( .A1(n524), .A2(n519), .ZN(n541) );
  XNOR2_X1 U612 ( .A(G110), .B(KEYINPUT114), .ZN(n520) );
  XNOR2_X1 U613 ( .A(n541), .B(n520), .ZN(G12) );
  XNOR2_X1 U614 ( .A(n521), .B(KEYINPUT102), .ZN(n662) );
  OR2_X1 U615 ( .A1(n369), .A2(n662), .ZN(n522) );
  NOR2_X1 U616 ( .A1(n522), .A2(n574), .ZN(n523) );
  NAND2_X1 U617 ( .A1(n524), .A2(n523), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(G101), .ZN(G3) );
  NAND2_X1 U619 ( .A1(n526), .A2(n525), .ZN(n533) );
  NOR2_X1 U620 ( .A1(n533), .A2(n598), .ZN(n527) );
  XNOR2_X1 U621 ( .A(n565), .B(G143), .ZN(G45) );
  NAND2_X1 U622 ( .A1(n531), .A2(n574), .ZN(n532) );
  INV_X1 U623 ( .A(n662), .ZN(n534) );
  NOR2_X1 U624 ( .A1(n529), .A2(n534), .ZN(n535) );
  XNOR2_X1 U625 ( .A(n535), .B(KEYINPUT103), .ZN(n536) );
  NOR2_X1 U626 ( .A1(n537), .A2(n536), .ZN(n539) );
  INV_X1 U627 ( .A(n574), .ZN(n538) );
  NAND2_X1 U628 ( .A1(n734), .A2(n541), .ZN(n542) );
  XNOR2_X1 U629 ( .A(n544), .B(n543), .ZN(n555) );
  NAND2_X1 U630 ( .A1(n548), .A2(n545), .ZN(n546) );
  NOR2_X1 U631 ( .A1(n546), .A2(n672), .ZN(n547) );
  XNOR2_X1 U632 ( .A(n547), .B(KEYINPUT31), .ZN(n654) );
  AND2_X1 U633 ( .A1(n548), .A2(n671), .ZN(n550) );
  NAND2_X1 U634 ( .A1(n550), .A2(n549), .ZN(n642) );
  NAND2_X1 U635 ( .A1(n654), .A2(n642), .ZN(n551) );
  NAND2_X1 U636 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U637 ( .A1(n555), .A2(n554), .ZN(n558) );
  INV_X1 U638 ( .A(KEYINPUT86), .ZN(n556) );
  XNOR2_X1 U639 ( .A(n556), .B(KEYINPUT45), .ZN(n557) );
  XNOR2_X1 U640 ( .A(n559), .B(KEYINPUT75), .ZN(n561) );
  INV_X1 U641 ( .A(n648), .ZN(n560) );
  NAND2_X1 U642 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U643 ( .A(n562), .B(KEYINPUT74), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n648), .A2(KEYINPUT47), .ZN(n563) );
  XNOR2_X1 U645 ( .A(n563), .B(KEYINPUT82), .ZN(n570) );
  NAND2_X1 U646 ( .A1(n683), .A2(KEYINPUT47), .ZN(n567) );
  INV_X1 U647 ( .A(KEYINPUT83), .ZN(n564) );
  XNOR2_X1 U648 ( .A(n565), .B(n564), .ZN(n566) );
  NAND2_X1 U649 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U650 ( .A(n568), .B(KEYINPUT81), .ZN(n569) );
  AND2_X1 U651 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U652 ( .A1(n572), .A2(n571), .ZN(n581) );
  INV_X1 U653 ( .A(n678), .ZN(n575) );
  NOR2_X1 U654 ( .A1(n652), .A2(n575), .ZN(n576) );
  XNOR2_X1 U655 ( .A(KEYINPUT91), .B(KEYINPUT36), .ZN(n578) );
  XNOR2_X1 U656 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U657 ( .A(n582), .B(KEYINPUT71), .ZN(n594) );
  NAND2_X1 U658 ( .A1(n679), .A2(n678), .ZN(n682) );
  INV_X1 U659 ( .A(n583), .ZN(n681) );
  NAND2_X1 U660 ( .A1(n693), .A2(n586), .ZN(n589) );
  INV_X1 U661 ( .A(KEYINPUT109), .ZN(n587) );
  XNOR2_X1 U662 ( .A(n587), .B(KEYINPUT42), .ZN(n588) );
  XNOR2_X1 U663 ( .A(n589), .B(n588), .ZN(n735) );
  NAND2_X1 U664 ( .A1(n590), .A2(n735), .ZN(n592) );
  XNOR2_X1 U665 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n591) );
  XNOR2_X1 U666 ( .A(n592), .B(n591), .ZN(n593) );
  NOR2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n596) );
  XNOR2_X1 U668 ( .A(KEYINPUT90), .B(KEYINPUT48), .ZN(n595) );
  XNOR2_X1 U669 ( .A(n596), .B(n595), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n348), .A2(n529), .ZN(n597) );
  XNOR2_X1 U671 ( .A(n597), .B(KEYINPUT43), .ZN(n599) );
  AND2_X1 U672 ( .A1(n598), .A2(n599), .ZN(n660) );
  INV_X1 U673 ( .A(n660), .ZN(n600) );
  INV_X1 U674 ( .A(KEYINPUT88), .ZN(n602) );
  INV_X1 U675 ( .A(KEYINPUT2), .ZN(n692) );
  NAND2_X1 U676 ( .A1(n629), .A2(G210), .ZN(n611) );
  XNOR2_X1 U677 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n608) );
  XNOR2_X1 U678 ( .A(KEYINPUT55), .B(KEYINPUT92), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n606), .B(n609), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n611), .B(n610), .ZN(n613) );
  INV_X1 U682 ( .A(G952), .ZN(n612) );
  NOR2_X1 U683 ( .A1(n613), .A2(n705), .ZN(n615) );
  XOR2_X1 U684 ( .A(KEYINPUT89), .B(KEYINPUT56), .Z(n614) );
  XNOR2_X1 U685 ( .A(n615), .B(n614), .ZN(G51) );
  NAND2_X1 U686 ( .A1(n629), .A2(G475), .ZN(n619) );
  XOR2_X1 U687 ( .A(KEYINPUT66), .B(KEYINPUT59), .Z(n616) );
  XNOR2_X1 U688 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X1 U690 ( .A1(n620), .A2(n705), .ZN(n621) );
  XNOR2_X1 U691 ( .A(n621), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U692 ( .A(KEYINPUT63), .ZN(n628) );
  NAND2_X1 U693 ( .A1(n629), .A2(G472), .ZN(n625) );
  XOR2_X1 U694 ( .A(KEYINPUT110), .B(KEYINPUT62), .Z(n622) );
  XNOR2_X1 U695 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U697 ( .A(n628), .B(n627), .ZN(G57) );
  BUF_X2 U698 ( .A(n629), .Z(n701) );
  XOR2_X1 U699 ( .A(n631), .B(n630), .Z(n632) );
  NOR2_X1 U700 ( .A1(n632), .A2(n705), .ZN(G66) );
  NAND2_X1 U701 ( .A1(n701), .A2(G469), .ZN(n638) );
  XOR2_X1 U702 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n634) );
  XNOR2_X1 U703 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n638), .B(n637), .ZN(n639) );
  NOR2_X1 U707 ( .A1(n639), .A2(n705), .ZN(G54) );
  NOR2_X1 U708 ( .A1(n642), .A2(n652), .ZN(n641) );
  XNOR2_X1 U709 ( .A(G104), .B(KEYINPUT111), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n641), .B(n640), .ZN(G6) );
  NOR2_X1 U711 ( .A1(n642), .A2(n655), .ZN(n647) );
  XOR2_X1 U712 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n644) );
  XNOR2_X1 U713 ( .A(G107), .B(KEYINPUT112), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U715 ( .A(KEYINPUT26), .B(n645), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(G9) );
  NOR2_X1 U717 ( .A1(n648), .A2(n655), .ZN(n650) );
  XNOR2_X1 U718 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U720 ( .A(G128), .B(n651), .Z(G30) );
  NOR2_X1 U721 ( .A1(n652), .A2(n654), .ZN(n653) );
  XOR2_X1 U722 ( .A(G113), .B(n653), .Z(G15) );
  NOR2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U724 ( .A(G116), .B(n656), .Z(G18) );
  XNOR2_X1 U725 ( .A(KEYINPUT116), .B(KEYINPUT37), .ZN(n657) );
  XNOR2_X1 U726 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U727 ( .A(G125), .B(n659), .ZN(G27) );
  XOR2_X1 U728 ( .A(G140), .B(n660), .Z(G42) );
  NAND2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U730 ( .A(n663), .B(KEYINPUT49), .ZN(n664) );
  XNOR2_X1 U731 ( .A(KEYINPUT117), .B(n664), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n665), .A2(n671), .ZN(n670) );
  NAND2_X1 U733 ( .A1(n529), .A2(n666), .ZN(n668) );
  XOR2_X1 U734 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n667) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n673) );
  OR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U739 ( .A(KEYINPUT51), .B(n675), .Z(n676) );
  NAND2_X1 U740 ( .A1(n693), .A2(n676), .ZN(n688) );
  NOR2_X1 U741 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U742 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n684) );
  OR2_X1 U744 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U745 ( .A1(n677), .A2(n686), .ZN(n687) );
  NAND2_X1 U746 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U747 ( .A(KEYINPUT52), .B(n689), .Z(n690) );
  NOR2_X1 U748 ( .A1(n691), .A2(n690), .ZN(n697) );
  XNOR2_X1 U749 ( .A(n605), .B(n692), .ZN(n695) );
  NAND2_X1 U750 ( .A1(n693), .A2(n677), .ZN(n694) );
  NAND2_X1 U751 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U752 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n698), .B(KEYINPUT119), .ZN(n699) );
  NOR2_X1 U754 ( .A1(G953), .A2(n699), .ZN(n700) );
  XNOR2_X1 U755 ( .A(KEYINPUT53), .B(n700), .ZN(G75) );
  NAND2_X1 U756 ( .A1(n701), .A2(G478), .ZN(n702) );
  XNOR2_X1 U757 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U758 ( .A1(n705), .A2(n704), .ZN(G63) );
  NAND2_X1 U759 ( .A1(n715), .A2(n706), .ZN(n710) );
  NAND2_X1 U760 ( .A1(G953), .A2(G224), .ZN(n707) );
  XNOR2_X1 U761 ( .A(KEYINPUT61), .B(n707), .ZN(n708) );
  NAND2_X1 U762 ( .A1(n708), .A2(G898), .ZN(n709) );
  NAND2_X1 U763 ( .A1(n710), .A2(n709), .ZN(n719) );
  XOR2_X1 U764 ( .A(n711), .B(KEYINPUT123), .Z(n712) );
  XNOR2_X1 U765 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n714), .B(G101), .ZN(n717) );
  NOR2_X1 U767 ( .A1(n715), .A2(G898), .ZN(n716) );
  NOR2_X1 U768 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U769 ( .A(n719), .B(n718), .ZN(G69) );
  XOR2_X1 U770 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n720) );
  XNOR2_X1 U771 ( .A(n721), .B(n720), .ZN(n722) );
  XOR2_X1 U772 ( .A(n723), .B(n722), .Z(n726) );
  XNOR2_X1 U773 ( .A(n724), .B(n726), .ZN(n725) );
  NOR2_X1 U774 ( .A1(n725), .A2(G953), .ZN(n731) );
  XNOR2_X1 U775 ( .A(n726), .B(G227), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U777 ( .A1(n728), .A2(G953), .ZN(n729) );
  XOR2_X1 U778 ( .A(KEYINPUT126), .B(n729), .Z(n730) );
  NOR2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U780 ( .A(KEYINPUT127), .B(n732), .ZN(G72) );
  XOR2_X1 U781 ( .A(G122), .B(n733), .Z(G24) );
  XNOR2_X1 U782 ( .A(G119), .B(n734), .ZN(G21) );
  XNOR2_X1 U783 ( .A(G137), .B(n735), .ZN(G39) );
endmodule

