

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793;

  NOR2_X1 U380 ( .A1(G953), .A2(G237), .ZN(n561) );
  INV_X1 U381 ( .A(KEYINPUT4), .ZN(n383) );
  XOR2_X1 U382 ( .A(G125), .B(G146), .Z(n575) );
  AND2_X2 U383 ( .A1(n405), .A2(n468), .ZN(n642) );
  XNOR2_X2 U384 ( .A(n651), .B(KEYINPUT31), .ZN(n699) );
  XNOR2_X2 U385 ( .A(n372), .B(n575), .ZN(n778) );
  NOR2_X2 U386 ( .A1(n666), .A2(n504), .ZN(n667) );
  INV_X4 U387 ( .A(G143), .ZN(n486) );
  XNOR2_X1 U388 ( .A(n658), .B(KEYINPUT102), .ZN(n793) );
  INV_X1 U389 ( .A(n456), .ZN(n716) );
  NOR2_X1 U390 ( .A1(n731), .A2(n732), .ZN(n611) );
  INV_X1 U391 ( .A(n408), .ZN(n361) );
  NOR2_X1 U392 ( .A1(n608), .A2(n607), .ZN(n616) );
  AND2_X1 U393 ( .A1(n376), .A2(n713), .ZN(n408) );
  NAND2_X1 U394 ( .A1(n483), .A2(n484), .ZN(n572) );
  BUF_X1 U395 ( .A(n539), .Z(n782) );
  AND2_X1 U396 ( .A1(n780), .A2(n706), .ZN(n709) );
  AND2_X2 U397 ( .A1(n628), .A2(n627), .ZN(n780) );
  XNOR2_X1 U398 ( .A(n435), .B(n445), .ZN(n628) );
  NOR2_X1 U399 ( .A1(n661), .A2(n660), .ZN(n665) );
  XNOR2_X1 U400 ( .A(n646), .B(KEYINPUT72), .ZN(n668) );
  NAND2_X1 U401 ( .A1(n452), .A2(KEYINPUT39), .ZN(n447) );
  XNOR2_X1 U402 ( .A(n639), .B(KEYINPUT32), .ZN(n791) );
  XNOR2_X1 U403 ( .A(n360), .B(KEYINPUT79), .ZN(n386) );
  AND2_X1 U404 ( .A1(n641), .A2(n716), .ZN(n654) );
  XNOR2_X1 U405 ( .A(n637), .B(n636), .ZN(n641) );
  NOR2_X1 U406 ( .A1(n716), .A2(n361), .ZN(n649) );
  NAND2_X1 U407 ( .A1(n716), .A2(n361), .ZN(n717) );
  XNOR2_X1 U408 ( .A(n369), .B(n392), .ZN(n412) );
  NAND2_X1 U409 ( .A1(n370), .A2(n634), .ZN(n369) );
  XNOR2_X1 U410 ( .A(n616), .B(KEYINPUT103), .ZN(n697) );
  INV_X1 U411 ( .A(n376), .ZN(n656) );
  XNOR2_X1 U412 ( .A(n544), .B(n377), .ZN(n376) );
  NOR2_X1 U413 ( .A1(n763), .A2(G902), .ZN(n544) );
  XNOR2_X1 U414 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U415 ( .A(n367), .B(n362), .ZN(n540) );
  XNOR2_X1 U416 ( .A(n366), .B(n363), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n538), .B(n572), .ZN(n366) );
  XNOR2_X1 U418 ( .A(n368), .B(n424), .ZN(n546) );
  XNOR2_X1 U419 ( .A(n592), .B(KEYINPUT88), .ZN(n371) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n363) );
  NAND2_X1 U421 ( .A1(n539), .A2(G234), .ZN(n368) );
  XNOR2_X1 U422 ( .A(G128), .B(G137), .ZN(n365) );
  XNOR2_X1 U423 ( .A(G101), .B(KEYINPUT68), .ZN(n519) );
  XNOR2_X1 U424 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n364) );
  XOR2_X1 U425 ( .A(KEYINPUT64), .B(G953), .Z(n539) );
  NAND2_X1 U426 ( .A1(n358), .A2(n662), .ZN(n663) );
  NAND2_X1 U427 ( .A1(n645), .A2(n358), .ZN(n646) );
  XNOR2_X1 U428 ( .A(n358), .B(G122), .ZN(G24) );
  XNOR2_X2 U429 ( .A(n458), .B(n457), .ZN(n358) );
  XNOR2_X2 U430 ( .A(n359), .B(n392), .ZN(n405) );
  NAND2_X1 U431 ( .A1(n381), .A2(n634), .ZN(n359) );
  XNOR2_X2 U432 ( .A(n374), .B(n592), .ZN(n381) );
  XNOR2_X2 U433 ( .A(n467), .B(KEYINPUT88), .ZN(n374) );
  NAND2_X1 U434 ( .A1(n598), .A2(n597), .ZN(n360) );
  NAND2_X1 U435 ( .A1(n546), .A2(G221), .ZN(n367) );
  XNOR2_X1 U436 ( .A(n467), .B(n371), .ZN(n370) );
  XOR2_X1 U437 ( .A(G140), .B(KEYINPUT10), .Z(n372) );
  INV_X1 U438 ( .A(n452), .ZN(n373) );
  INV_X1 U439 ( .A(n410), .ZN(n409) );
  BUF_X2 U440 ( .A(n586), .Z(n587) );
  XNOR2_X1 U441 ( .A(G475), .B(n570), .ZN(n375) );
  XNOR2_X1 U442 ( .A(G475), .B(n570), .ZN(n608) );
  XOR2_X1 U443 ( .A(n543), .B(n542), .Z(n377) );
  INV_X1 U444 ( .A(n413), .ZN(n378) );
  BUF_X1 U445 ( .A(n647), .Z(n379) );
  NAND2_X1 U446 ( .A1(n448), .A2(n447), .ZN(n380) );
  NAND2_X1 U447 ( .A1(n448), .A2(n447), .ZN(n624) );
  NAND2_X1 U448 ( .A1(n553), .A2(KEYINPUT4), .ZN(n384) );
  NAND2_X1 U449 ( .A1(n382), .A2(n383), .ZN(n385) );
  NAND2_X1 U450 ( .A1(n384), .A2(n385), .ZN(n509) );
  INV_X1 U451 ( .A(n553), .ZN(n382) );
  INV_X1 U452 ( .A(n409), .ZN(n387) );
  INV_X1 U453 ( .A(KEYINPUT33), .ZN(n498) );
  NOR2_X1 U454 ( .A1(n694), .A2(n414), .ZN(n428) );
  NAND2_X1 U455 ( .A1(n652), .A2(n415), .ZN(n414) );
  INV_X1 U456 ( .A(KEYINPUT75), .ZN(n427) );
  XNOR2_X1 U457 ( .A(G902), .B(KEYINPUT15), .ZN(n523) );
  XOR2_X1 U458 ( .A(KEYINPUT4), .B(KEYINPUT18), .Z(n577) );
  OR2_X1 U459 ( .A1(G902), .A2(G237), .ZN(n581) );
  XOR2_X1 U460 ( .A(G119), .B(KEYINPUT5), .Z(n517) );
  XNOR2_X1 U461 ( .A(n515), .B(KEYINPUT3), .ZN(n573) );
  INV_X1 U462 ( .A(n523), .ZN(n676) );
  INV_X1 U463 ( .A(G146), .ZN(n510) );
  INV_X1 U464 ( .A(KEYINPUT1), .ZN(n455) );
  XOR2_X1 U465 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n526) );
  INV_X1 U466 ( .A(KEYINPUT8), .ZN(n424) );
  XNOR2_X1 U467 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U468 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n549) );
  INV_X1 U469 ( .A(KEYINPUT36), .ZN(n430) );
  XNOR2_X1 U470 ( .A(n642), .B(KEYINPUT34), .ZN(n459) );
  NOR2_X1 U471 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U472 ( .A1(n792), .A2(n444), .ZN(n442) );
  NAND2_X1 U473 ( .A1(n440), .A2(n439), .ZN(n438) );
  XOR2_X1 U474 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n563) );
  XOR2_X1 U475 ( .A(G113), .B(G104), .Z(n558) );
  XNOR2_X1 U476 ( .A(n413), .B(G122), .ZN(n557) );
  NAND2_X1 U477 ( .A1(n676), .A2(n496), .ZN(n495) );
  INV_X1 U478 ( .A(KEYINPUT65), .ZN(n496) );
  XOR2_X1 U479 ( .A(G110), .B(G140), .Z(n512) );
  NAND2_X1 U480 ( .A1(n782), .A2(G224), .ZN(n477) );
  XNOR2_X1 U481 ( .A(KEYINPUT81), .B(KEYINPUT17), .ZN(n576) );
  XNOR2_X1 U482 ( .A(n473), .B(n765), .ZN(n574) );
  XNOR2_X1 U483 ( .A(n519), .B(n474), .ZN(n473) );
  INV_X1 U484 ( .A(KEYINPUT71), .ZN(n474) );
  NAND2_X1 U485 ( .A1(G237), .A2(G234), .ZN(n528) );
  INV_X1 U486 ( .A(KEYINPUT48), .ZN(n445) );
  XNOR2_X1 U487 ( .A(KEYINPUT91), .B(n582), .ZN(n618) );
  XNOR2_X1 U488 ( .A(n521), .B(n573), .ZN(n501) );
  XOR2_X1 U489 ( .A(G107), .B(G104), .Z(n765) );
  NAND2_X1 U490 ( .A1(n523), .A2(KEYINPUT65), .ZN(n490) );
  NAND2_X1 U491 ( .A1(n493), .A2(n492), .ZN(n491) );
  XNOR2_X1 U492 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n636) );
  NAND2_X1 U493 ( .A1(n409), .A2(n408), .ZN(n647) );
  INV_X1 U494 ( .A(KEYINPUT6), .ZN(n500) );
  XNOR2_X1 U495 ( .A(n552), .B(n551), .ZN(n554) );
  XNOR2_X1 U496 ( .A(n681), .B(n680), .ZN(n682) );
  INV_X1 U497 ( .A(G953), .ZN(n772) );
  XNOR2_X1 U498 ( .A(n621), .B(n425), .ZN(n622) );
  XNOR2_X1 U499 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n425) );
  XNOR2_X1 U500 ( .A(n584), .B(n429), .ZN(n585) );
  XNOR2_X1 U501 ( .A(n430), .B(KEYINPUT87), .ZN(n429) );
  XNOR2_X1 U502 ( .A(KEYINPUT85), .B(KEYINPUT35), .ZN(n457) );
  NAND2_X1 U503 ( .A1(n459), .A2(n644), .ZN(n458) );
  INV_X1 U504 ( .A(n721), .ZN(n469) );
  BUF_X1 U505 ( .A(G143), .Z(n413) );
  INV_X1 U506 ( .A(KEYINPUT124), .ZN(n432) );
  INV_X1 U507 ( .A(KEYINPUT60), .ZN(n418) );
  AND2_X1 U508 ( .A1(n713), .A2(n635), .ZN(n388) );
  AND2_X1 U509 ( .A1(n675), .A2(KEYINPUT65), .ZN(n389) );
  OR2_X1 U510 ( .A1(n415), .A2(n594), .ZN(n390) );
  XOR2_X1 U511 ( .A(n579), .B(KEYINPUT90), .Z(n391) );
  XNOR2_X1 U512 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n392) );
  XOR2_X1 U513 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n393) );
  NOR2_X1 U514 ( .A1(n782), .A2(G952), .ZN(n764) );
  INV_X1 U515 ( .A(n764), .ZN(n463) );
  XOR2_X1 U516 ( .A(n677), .B(n503), .Z(n394) );
  INV_X1 U517 ( .A(KEYINPUT47), .ZN(n415) );
  XNOR2_X1 U518 ( .A(n760), .B(KEYINPUT59), .ZN(n395) );
  XOR2_X1 U519 ( .A(KEYINPUT63), .B(KEYINPUT111), .Z(n396) );
  XOR2_X1 U520 ( .A(KEYINPUT86), .B(KEYINPUT56), .Z(n397) );
  XNOR2_X1 U521 ( .A(n779), .B(n510), .ZN(n398) );
  XNOR2_X1 U522 ( .A(n779), .B(n510), .ZN(n407) );
  AND2_X1 U523 ( .A1(n456), .A2(n408), .ZN(n426) );
  INV_X1 U524 ( .A(n729), .ZN(n615) );
  XNOR2_X1 U525 ( .A(n410), .B(n455), .ZN(n456) );
  BUF_X1 U526 ( .A(n773), .Z(n399) );
  AND2_X1 U527 ( .A1(n656), .A2(n400), .ZN(n629) );
  NOR2_X1 U528 ( .A1(n716), .A2(n655), .ZN(n400) );
  NAND2_X1 U529 ( .A1(n654), .A2(n657), .ZN(n658) );
  BUF_X1 U530 ( .A(n753), .Z(n401) );
  BUF_X1 U531 ( .A(n553), .Z(n402) );
  XNOR2_X1 U532 ( .A(n407), .B(n506), .ZN(n753) );
  AND2_X1 U533 ( .A1(n780), .A2(KEYINPUT2), .ZN(n671) );
  BUF_X1 U534 ( .A(n411), .Z(n403) );
  XNOR2_X1 U535 ( .A(n578), .B(n477), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n478), .B(n573), .ZN(n411) );
  XNOR2_X1 U537 ( .A(n378), .B(G128), .ZN(n404) );
  NAND2_X1 U538 ( .A1(n426), .A2(n655), .ZN(n499) );
  NAND2_X1 U539 ( .A1(n441), .A2(n438), .ZN(n436) );
  XNOR2_X1 U540 ( .A(n411), .B(n476), .ZN(n475) );
  BUF_X1 U541 ( .A(n679), .Z(n406) );
  XNOR2_X1 U542 ( .A(n475), .B(n471), .ZN(n679) );
  AND2_X1 U543 ( .A1(n780), .A2(KEYINPUT78), .ZN(n669) );
  XNOR2_X1 U544 ( .A(n482), .B(n481), .ZN(n480) );
  XNOR2_X1 U545 ( .A(n454), .B(n682), .ZN(n453) );
  XNOR2_X1 U546 ( .A(n485), .B(n572), .ZN(n478) );
  XNOR2_X1 U547 ( .A(n502), .B(G122), .ZN(n485) );
  NAND2_X1 U548 ( .A1(n453), .A2(n463), .ZN(n431) );
  NAND2_X1 U549 ( .A1(n756), .A2(G217), .ZN(n482) );
  NAND2_X1 U550 ( .A1(n756), .A2(G210), .ZN(n454) );
  XNOR2_X1 U551 ( .A(n398), .B(n501), .ZN(n677) );
  NOR2_X1 U552 ( .A1(n591), .A2(n387), .ZN(n606) );
  XNOR2_X2 U553 ( .A(n514), .B(G469), .ZN(n410) );
  XNOR2_X1 U554 ( .A(n403), .B(n766), .ZN(n768) );
  NAND2_X1 U555 ( .A1(n412), .A2(n388), .ZN(n637) );
  AND2_X1 U556 ( .A1(n405), .A2(n469), .ZN(n651) );
  AND2_X1 U557 ( .A1(n405), .A2(n470), .ZN(n648) );
  NAND2_X1 U558 ( .A1(n654), .A2(n640), .ZN(n690) );
  NAND2_X1 U559 ( .A1(n791), .A2(n690), .ZN(n479) );
  AND2_X2 U560 ( .A1(n416), .A2(n450), .ZN(n448) );
  NAND2_X1 U561 ( .A1(n446), .A2(n386), .ZN(n416) );
  XNOR2_X2 U562 ( .A(n417), .B(KEYINPUT30), .ZN(n599) );
  NOR2_X2 U563 ( .A1(n587), .A2(n618), .ZN(n417) );
  XNOR2_X1 U564 ( .A(n419), .B(n418), .ZN(G60) );
  NAND2_X1 U565 ( .A1(n421), .A2(n463), .ZN(n419) );
  XNOR2_X1 U566 ( .A(n420), .B(n396), .ZN(G57) );
  NAND2_X1 U567 ( .A1(n422), .A2(n463), .ZN(n420) );
  XNOR2_X1 U568 ( .A(n761), .B(n395), .ZN(n421) );
  XNOR2_X1 U569 ( .A(n678), .B(n394), .ZN(n422) );
  XNOR2_X1 U570 ( .A(KEYINPUT41), .B(n611), .ZN(n727) );
  NAND2_X1 U571 ( .A1(n729), .A2(n728), .ZN(n732) );
  XNOR2_X2 U572 ( .A(n423), .B(KEYINPUT45), .ZN(n773) );
  NAND2_X1 U573 ( .A1(n667), .A2(n668), .ZN(n423) );
  NAND2_X1 U574 ( .A1(n571), .A2(n655), .ZN(n617) );
  XNOR2_X1 U575 ( .A(n580), .B(n391), .ZN(n505) );
  NAND2_X1 U576 ( .A1(n479), .A2(KEYINPUT66), .ZN(n662) );
  NOR2_X2 U577 ( .A1(n753), .A2(G902), .ZN(n514) );
  NAND2_X1 U578 ( .A1(n793), .A2(n659), .ZN(n661) );
  XNOR2_X1 U579 ( .A(n428), .B(n427), .ZN(n603) );
  XNOR2_X1 U580 ( .A(n617), .B(KEYINPUT109), .ZN(n583) );
  NOR2_X1 U581 ( .A1(n497), .A2(n495), .ZN(n494) );
  XNOR2_X1 U582 ( .A(n431), .B(n397), .ZN(G51) );
  XNOR2_X1 U583 ( .A(n433), .B(n432), .ZN(G66) );
  NAND2_X1 U584 ( .A1(n480), .A2(n463), .ZN(n433) );
  XNOR2_X2 U585 ( .A(n623), .B(n610), .ZN(n729) );
  NAND2_X1 U586 ( .A1(n756), .A2(G475), .ZN(n761) );
  NAND2_X1 U587 ( .A1(n756), .A2(G472), .ZN(n678) );
  NAND2_X1 U588 ( .A1(n756), .A2(G478), .ZN(n466) );
  NAND2_X2 U589 ( .A1(n488), .A2(n487), .ZN(n756) );
  NOR2_X1 U590 ( .A1(n702), .A2(n434), .ZN(n437) );
  NAND2_X1 U591 ( .A1(n605), .A2(n390), .ZN(n434) );
  NAND2_X1 U592 ( .A1(n789), .A2(n444), .ZN(n443) );
  NAND2_X1 U593 ( .A1(n436), .A2(n437), .ZN(n435) );
  INV_X1 U594 ( .A(n789), .ZN(n439) );
  NOR2_X1 U595 ( .A1(n792), .A2(n444), .ZN(n440) );
  AND2_X1 U596 ( .A1(n443), .A2(n442), .ZN(n441) );
  INV_X1 U597 ( .A(KEYINPUT46), .ZN(n444) );
  AND2_X1 U598 ( .A1(n449), .A2(n599), .ZN(n446) );
  INV_X1 U599 ( .A(n386), .ZN(n452) );
  NAND2_X1 U600 ( .A1(n373), .A2(n599), .ZN(n614) );
  NOR2_X1 U601 ( .A1(n615), .A2(KEYINPUT39), .ZN(n449) );
  NAND2_X1 U602 ( .A1(n451), .A2(KEYINPUT39), .ZN(n450) );
  NAND2_X1 U603 ( .A1(n599), .A2(n729), .ZN(n451) );
  XNOR2_X2 U604 ( .A(n460), .B(n507), .ZN(n553) );
  XNOR2_X1 U605 ( .A(n404), .B(n575), .ZN(n472) );
  XNOR2_X2 U606 ( .A(n486), .B(G128), .ZN(n460) );
  XNOR2_X2 U607 ( .A(n461), .B(n393), .ZN(n789) );
  NAND2_X1 U608 ( .A1(n624), .A2(n616), .ZN(n461) );
  XNOR2_X1 U609 ( .A(n462), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U610 ( .A1(n464), .A2(n463), .ZN(n462) );
  XNOR2_X1 U611 ( .A(n466), .B(n465), .ZN(n464) );
  INV_X1 U612 ( .A(n762), .ZN(n465) );
  NOR2_X2 U613 ( .A1(n505), .A2(n618), .ZN(n467) );
  INV_X1 U614 ( .A(n737), .ZN(n468) );
  INV_X1 U615 ( .A(n379), .ZN(n470) );
  XNOR2_X1 U616 ( .A(n574), .B(n472), .ZN(n471) );
  NOR2_X1 U617 ( .A1(n479), .A2(KEYINPUT66), .ZN(n660) );
  NOR2_X1 U618 ( .A1(n479), .A2(KEYINPUT44), .ZN(n645) );
  INV_X1 U619 ( .A(n763), .ZN(n481) );
  NAND2_X1 U620 ( .A1(n537), .A2(G110), .ZN(n484) );
  NAND2_X1 U621 ( .A1(n536), .A2(G119), .ZN(n483) );
  INV_X1 U622 ( .A(n675), .ZN(n493) );
  NAND2_X1 U623 ( .A1(n491), .A2(n490), .ZN(n489) );
  NOR2_X1 U624 ( .A1(n494), .A2(n489), .ZN(n488) );
  NAND2_X1 U625 ( .A1(n497), .A2(n389), .ZN(n487) );
  INV_X1 U626 ( .A(n495), .ZN(n492) );
  NAND2_X1 U627 ( .A1(n673), .A2(n672), .ZN(n497) );
  XNOR2_X2 U628 ( .A(n499), .B(n498), .ZN(n737) );
  XNOR2_X2 U629 ( .A(n650), .B(n500), .ZN(n655) );
  XNOR2_X2 U630 ( .A(n509), .B(n508), .ZN(n779) );
  XNOR2_X2 U631 ( .A(KEYINPUT16), .B(KEYINPUT74), .ZN(n502) );
  XNOR2_X1 U632 ( .A(KEYINPUT62), .B(KEYINPUT110), .ZN(n503) );
  NOR2_X1 U633 ( .A1(KEYINPUT44), .A2(KEYINPUT66), .ZN(n504) );
  XOR2_X1 U634 ( .A(n574), .B(n513), .Z(n506) );
  INV_X1 U635 ( .A(KEYINPUT106), .ZN(n596) );
  INV_X1 U636 ( .A(n704), .ZN(n626) );
  XNOR2_X1 U637 ( .A(n647), .B(n596), .ZN(n598) );
  INV_X1 U638 ( .A(G134), .ZN(n507) );
  XNOR2_X1 U639 ( .A(n522), .B(G472), .ZN(n586) );
  INV_X1 U640 ( .A(KEYINPUT19), .ZN(n592) );
  XOR2_X1 U641 ( .A(KEYINPUT69), .B(G131), .Z(n560) );
  XOR2_X1 U642 ( .A(G137), .B(n560), .Z(n508) );
  NAND2_X1 U643 ( .A1(G227), .A2(n782), .ZN(n511) );
  XNOR2_X1 U644 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U645 ( .A(G116), .B(G113), .ZN(n515) );
  NAND2_X1 U646 ( .A1(n561), .A2(G210), .ZN(n516) );
  XNOR2_X1 U647 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U648 ( .A(KEYINPUT97), .B(n518), .ZN(n520) );
  XNOR2_X1 U649 ( .A(n520), .B(n519), .ZN(n521) );
  NOR2_X1 U650 ( .A1(n677), .A2(G902), .ZN(n522) );
  INV_X1 U651 ( .A(n586), .ZN(n650) );
  NAND2_X1 U652 ( .A1(G234), .A2(n523), .ZN(n524) );
  XNOR2_X1 U653 ( .A(KEYINPUT20), .B(n524), .ZN(n541) );
  NAND2_X1 U654 ( .A1(G221), .A2(n541), .ZN(n525) );
  XNOR2_X1 U655 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U656 ( .A(KEYINPUT95), .B(n527), .Z(n713) );
  XNOR2_X1 U657 ( .A(n528), .B(KEYINPUT14), .ZN(n529) );
  XNOR2_X1 U658 ( .A(KEYINPUT76), .B(n529), .ZN(n531) );
  NAND2_X1 U659 ( .A1(G952), .A2(n531), .ZN(n744) );
  NOR2_X1 U660 ( .A1(G953), .A2(n744), .ZN(n530) );
  XOR2_X1 U661 ( .A(KEYINPUT92), .B(n530), .Z(n632) );
  NAND2_X1 U662 ( .A1(G902), .A2(n531), .ZN(n630) );
  NOR2_X1 U663 ( .A1(G900), .A2(n630), .ZN(n533) );
  INV_X1 U664 ( .A(n782), .ZN(n532) );
  NAND2_X1 U665 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U666 ( .A1(n632), .A2(n534), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n713), .A2(n597), .ZN(n535) );
  XOR2_X1 U668 ( .A(KEYINPUT70), .B(n535), .Z(n545) );
  INV_X1 U669 ( .A(G110), .ZN(n536) );
  INV_X1 U670 ( .A(G119), .ZN(n537) );
  XNOR2_X1 U671 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n538) );
  XNOR2_X1 U672 ( .A(n540), .B(n778), .ZN(n763) );
  XOR2_X1 U673 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n543) );
  NAND2_X1 U674 ( .A1(n541), .A2(G217), .ZN(n542) );
  NAND2_X1 U675 ( .A1(n545), .A2(n656), .ZN(n588) );
  NAND2_X1 U676 ( .A1(G217), .A2(n546), .ZN(n552) );
  XOR2_X1 U677 ( .A(KEYINPUT7), .B(G122), .Z(n548) );
  XNOR2_X1 U678 ( .A(G107), .B(G116), .ZN(n547) );
  XNOR2_X1 U679 ( .A(n548), .B(n547), .ZN(n550) );
  XNOR2_X1 U680 ( .A(n402), .B(n554), .ZN(n762) );
  NOR2_X1 U681 ( .A1(n762), .A2(G902), .ZN(n555) );
  XNOR2_X1 U682 ( .A(G478), .B(n555), .ZN(n556) );
  XNOR2_X1 U683 ( .A(n556), .B(KEYINPUT101), .ZN(n607) );
  XNOR2_X1 U684 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n569) );
  XNOR2_X1 U685 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U686 ( .A(n778), .B(n559), .Z(n567) );
  XNOR2_X1 U687 ( .A(n560), .B(KEYINPUT98), .ZN(n565) );
  NAND2_X1 U688 ( .A1(n561), .A2(G214), .ZN(n562) );
  XNOR2_X1 U689 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U690 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U691 ( .A(n567), .B(n566), .ZN(n760) );
  NOR2_X1 U692 ( .A1(G902), .A2(n760), .ZN(n568) );
  NOR2_X1 U693 ( .A1(n588), .A2(n697), .ZN(n571) );
  XNOR2_X1 U694 ( .A(n577), .B(n576), .ZN(n578) );
  NOR2_X1 U695 ( .A1(n679), .A2(n676), .ZN(n580) );
  NAND2_X1 U696 ( .A1(n581), .A2(G210), .ZN(n579) );
  NAND2_X1 U697 ( .A1(G214), .A2(n581), .ZN(n582) );
  NAND2_X1 U698 ( .A1(n583), .A2(n374), .ZN(n584) );
  NOR2_X2 U699 ( .A1(n716), .A2(n585), .ZN(n702) );
  XOR2_X1 U700 ( .A(KEYINPUT28), .B(KEYINPUT107), .Z(n590) );
  OR2_X1 U701 ( .A1(n588), .A2(n586), .ZN(n589) );
  XNOR2_X1 U702 ( .A(n590), .B(n589), .ZN(n591) );
  NAND2_X1 U703 ( .A1(n606), .A2(n381), .ZN(n694) );
  NAND2_X1 U704 ( .A1(n607), .A2(n375), .ZN(n700) );
  INV_X1 U705 ( .A(n700), .ZN(n625) );
  NOR2_X1 U706 ( .A1(n625), .A2(n616), .ZN(n733) );
  INV_X1 U707 ( .A(n733), .ZN(n652) );
  NOR2_X1 U708 ( .A1(KEYINPUT83), .A2(n652), .ZN(n593) );
  NOR2_X1 U709 ( .A1(n694), .A2(n593), .ZN(n594) );
  NAND2_X1 U710 ( .A1(KEYINPUT47), .A2(n733), .ZN(n595) );
  NAND2_X1 U711 ( .A1(n595), .A2(KEYINPUT83), .ZN(n602) );
  INV_X1 U712 ( .A(n375), .ZN(n600) );
  NAND2_X1 U713 ( .A1(n607), .A2(n600), .ZN(n643) );
  NOR2_X1 U714 ( .A1(n614), .A2(n643), .ZN(n601) );
  INV_X1 U715 ( .A(n505), .ZN(n623) );
  NAND2_X1 U716 ( .A1(n601), .A2(n623), .ZN(n693) );
  NAND2_X1 U717 ( .A1(n602), .A2(n693), .ZN(n604) );
  INV_X1 U718 ( .A(n606), .ZN(n612) );
  INV_X1 U719 ( .A(n607), .ZN(n609) );
  NAND2_X1 U720 ( .A1(n609), .A2(n375), .ZN(n731) );
  XNOR2_X1 U721 ( .A(KEYINPUT38), .B(KEYINPUT77), .ZN(n610) );
  INV_X1 U722 ( .A(n618), .ZN(n728) );
  NOR2_X1 U723 ( .A1(n612), .A2(n727), .ZN(n613) );
  XNOR2_X1 U724 ( .A(n613), .B(KEYINPUT42), .ZN(n792) );
  NOR2_X1 U725 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U726 ( .A(KEYINPUT104), .B(n619), .ZN(n620) );
  NAND2_X1 U727 ( .A1(n620), .A2(n716), .ZN(n621) );
  NOR2_X1 U728 ( .A1(n623), .A2(n622), .ZN(n705) );
  NAND2_X1 U729 ( .A1(n625), .A2(n380), .ZN(n704) );
  NOR2_X1 U730 ( .A1(n705), .A2(n626), .ZN(n627) );
  XNOR2_X1 U731 ( .A(KEYINPUT82), .B(n629), .ZN(n638) );
  INV_X1 U732 ( .A(n630), .ZN(n631) );
  NOR2_X1 U733 ( .A1(G898), .A2(n772), .ZN(n767) );
  NAND2_X1 U734 ( .A1(n631), .A2(n767), .ZN(n633) );
  NAND2_X1 U735 ( .A1(n633), .A2(n632), .ZN(n634) );
  INV_X1 U736 ( .A(n731), .ZN(n635) );
  NAND2_X1 U737 ( .A1(n641), .A2(n638), .ZN(n639) );
  AND2_X1 U738 ( .A1(n656), .A2(n587), .ZN(n640) );
  INV_X1 U739 ( .A(n643), .ZN(n644) );
  NAND2_X1 U740 ( .A1(n648), .A2(n587), .ZN(n685) );
  NAND2_X1 U741 ( .A1(n650), .A2(n649), .ZN(n721) );
  NAND2_X1 U742 ( .A1(n685), .A2(n699), .ZN(n653) );
  NAND2_X1 U743 ( .A1(n653), .A2(n652), .ZN(n659) );
  NOR2_X1 U744 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U745 ( .A1(n663), .A2(KEYINPUT44), .ZN(n664) );
  NAND2_X1 U746 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n773), .A2(n669), .ZN(n670) );
  INV_X1 U748 ( .A(KEYINPUT2), .ZN(n706) );
  NAND2_X1 U749 ( .A1(n670), .A2(n706), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n671), .A2(n773), .ZN(n672) );
  NOR2_X1 U751 ( .A1(n780), .A2(KEYINPUT78), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n773), .A2(n674), .ZN(n675) );
  XOR2_X1 U753 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n681) );
  XNOR2_X1 U754 ( .A(n406), .B(KEYINPUT89), .ZN(n680) );
  NOR2_X1 U755 ( .A1(n697), .A2(n685), .ZN(n683) );
  XOR2_X1 U756 ( .A(KEYINPUT112), .B(n683), .Z(n684) );
  XNOR2_X1 U757 ( .A(G104), .B(n684), .ZN(G6) );
  NOR2_X1 U758 ( .A1(n685), .A2(n700), .ZN(n689) );
  XOR2_X1 U759 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n687) );
  XNOR2_X1 U760 ( .A(G107), .B(KEYINPUT113), .ZN(n686) );
  XNOR2_X1 U761 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U762 ( .A(n689), .B(n688), .ZN(G9) );
  XNOR2_X1 U763 ( .A(n690), .B(G110), .ZN(G12) );
  NOR2_X1 U764 ( .A1(n700), .A2(n694), .ZN(n692) );
  XNOR2_X1 U765 ( .A(G128), .B(KEYINPUT29), .ZN(n691) );
  XNOR2_X1 U766 ( .A(n692), .B(n691), .ZN(G30) );
  XNOR2_X1 U767 ( .A(n413), .B(n693), .ZN(G45) );
  NOR2_X1 U768 ( .A1(n697), .A2(n694), .ZN(n695) );
  XOR2_X1 U769 ( .A(KEYINPUT114), .B(n695), .Z(n696) );
  XNOR2_X1 U770 ( .A(G146), .B(n696), .ZN(G48) );
  NOR2_X1 U771 ( .A1(n697), .A2(n699), .ZN(n698) );
  XOR2_X1 U772 ( .A(G113), .B(n698), .Z(G15) );
  NOR2_X1 U773 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U774 ( .A(G116), .B(n701), .Z(G18) );
  XNOR2_X1 U775 ( .A(G125), .B(n702), .ZN(n703) );
  XNOR2_X1 U776 ( .A(n703), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U777 ( .A(G134), .B(n704), .ZN(G36) );
  XOR2_X1 U778 ( .A(G140), .B(n705), .Z(G42) );
  AND2_X1 U779 ( .A1(n399), .A2(n780), .ZN(n707) );
  NOR2_X1 U780 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U781 ( .A1(n709), .A2(n708), .ZN(n712) );
  NOR2_X1 U782 ( .A1(KEYINPUT2), .A2(n399), .ZN(n710) );
  XNOR2_X1 U783 ( .A(n710), .B(KEYINPUT84), .ZN(n711) );
  NOR2_X1 U784 ( .A1(n712), .A2(n711), .ZN(n750) );
  NOR2_X1 U785 ( .A1(n727), .A2(n737), .ZN(n747) );
  XOR2_X1 U786 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n743) );
  NOR2_X1 U787 ( .A1(n376), .A2(n713), .ZN(n714) );
  XNOR2_X1 U788 ( .A(n714), .B(KEYINPUT49), .ZN(n715) );
  NAND2_X1 U789 ( .A1(n587), .A2(n715), .ZN(n719) );
  XOR2_X1 U790 ( .A(KEYINPUT50), .B(n717), .Z(n718) );
  NOR2_X1 U791 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U792 ( .A(KEYINPUT115), .B(n720), .ZN(n722) );
  NAND2_X1 U793 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U794 ( .A(n723), .B(KEYINPUT117), .ZN(n725) );
  XOR2_X1 U795 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n724) );
  XNOR2_X1 U796 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U797 ( .A1(n727), .A2(n726), .ZN(n740) );
  NOR2_X1 U798 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U799 ( .A1(n731), .A2(n730), .ZN(n736) );
  NOR2_X1 U800 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U801 ( .A(n734), .B(KEYINPUT118), .ZN(n735) );
  NOR2_X1 U802 ( .A1(n736), .A2(n735), .ZN(n738) );
  NOR2_X1 U803 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U804 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U805 ( .A(n741), .B(KEYINPUT52), .ZN(n742) );
  XNOR2_X1 U806 ( .A(n743), .B(n742), .ZN(n745) );
  NOR2_X1 U807 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U808 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U809 ( .A(n748), .B(KEYINPUT121), .ZN(n749) );
  NOR2_X1 U810 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U811 ( .A1(n772), .A2(n751), .ZN(n752) );
  XOR2_X1 U812 ( .A(KEYINPUT53), .B(n752), .Z(G75) );
  XNOR2_X1 U813 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n755) );
  XNOR2_X1 U814 ( .A(n401), .B(KEYINPUT57), .ZN(n754) );
  XNOR2_X1 U815 ( .A(n755), .B(n754), .ZN(n758) );
  NAND2_X1 U816 ( .A1(n756), .A2(G469), .ZN(n757) );
  XOR2_X1 U817 ( .A(n758), .B(n757), .Z(n759) );
  NOR2_X1 U818 ( .A1(n764), .A2(n759), .ZN(G54) );
  XNOR2_X1 U819 ( .A(n765), .B(G101), .ZN(n766) );
  NOR2_X1 U820 ( .A1(n768), .A2(n767), .ZN(n777) );
  XOR2_X1 U821 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n770) );
  NAND2_X1 U822 ( .A1(G224), .A2(G953), .ZN(n769) );
  XNOR2_X1 U823 ( .A(n770), .B(n769), .ZN(n771) );
  NAND2_X1 U824 ( .A1(n771), .A2(G898), .ZN(n775) );
  NAND2_X1 U825 ( .A1(n399), .A2(n772), .ZN(n774) );
  NAND2_X1 U826 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U827 ( .A(n777), .B(n776), .ZN(G69) );
  XOR2_X1 U828 ( .A(n778), .B(n779), .Z(n783) );
  XNOR2_X1 U829 ( .A(n780), .B(n783), .ZN(n781) );
  NAND2_X1 U830 ( .A1(n782), .A2(n781), .ZN(n788) );
  XOR2_X1 U831 ( .A(G227), .B(n783), .Z(n784) );
  XNOR2_X1 U832 ( .A(n784), .B(KEYINPUT126), .ZN(n785) );
  NAND2_X1 U833 ( .A1(n785), .A2(G900), .ZN(n786) );
  NAND2_X1 U834 ( .A1(G953), .A2(n786), .ZN(n787) );
  NAND2_X1 U835 ( .A1(n788), .A2(n787), .ZN(G72) );
  XNOR2_X1 U836 ( .A(G131), .B(n789), .ZN(n790) );
  XNOR2_X1 U837 ( .A(n790), .B(KEYINPUT127), .ZN(G33) );
  XNOR2_X1 U838 ( .A(n791), .B(G119), .ZN(G21) );
  XOR2_X1 U839 ( .A(G137), .B(n792), .Z(G39) );
  XNOR2_X1 U840 ( .A(G101), .B(n793), .ZN(G3) );
endmodule

