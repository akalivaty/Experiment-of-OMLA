

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U546 ( .A(KEYINPUT28), .ZN(n719) );
  NOR2_X1 U547 ( .A1(n697), .A2(n696), .ZN(n698) );
  AND2_X1 U548 ( .A1(G137), .A2(n873), .ZN(n513) );
  XOR2_X1 U549 ( .A(KEYINPUT23), .B(n518), .Z(n514) );
  NOR2_X1 U550 ( .A1(n771), .A2(n752), .ZN(n515) );
  BUF_X1 U551 ( .A(n692), .Z(n730) );
  NOR2_X1 U552 ( .A1(G1966), .A2(n771), .ZN(n741) );
  XNOR2_X1 U553 ( .A(n689), .B(KEYINPUT64), .ZN(n692) );
  OR2_X1 U554 ( .A1(n761), .A2(n760), .ZN(n767) );
  NOR2_X2 U555 ( .A1(G2105), .A2(n517), .ZN(n875) );
  NOR2_X1 U556 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  AND2_X1 U557 ( .A1(n808), .A2(n816), .ZN(n809) );
  NOR2_X1 U558 ( .A1(G651), .A2(n634), .ZN(n646) );
  NAND2_X1 U559 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U560 ( .A(n524), .B(KEYINPUT65), .ZN(n687) );
  BUF_X1 U561 ( .A(n687), .Z(G160) );
  INV_X1 U562 ( .A(G2105), .ZN(n516) );
  NOR2_X1 U563 ( .A1(G2104), .A2(n516), .ZN(n870) );
  NAND2_X1 U564 ( .A1(G125), .A2(n870), .ZN(n523) );
  INV_X1 U565 ( .A(G2104), .ZN(n517) );
  NOR2_X1 U566 ( .A1(n516), .A2(n517), .ZN(n869) );
  NAND2_X1 U567 ( .A1(G113), .A2(n869), .ZN(n519) );
  NAND2_X1 U568 ( .A1(G101), .A2(n875), .ZN(n518) );
  NAND2_X1 U569 ( .A1(n519), .A2(n514), .ZN(n521) );
  XOR2_X2 U570 ( .A(KEYINPUT17), .B(n520), .Z(n873) );
  NOR2_X1 U571 ( .A1(n521), .A2(n513), .ZN(n522) );
  INV_X1 U572 ( .A(G651), .ZN(n532) );
  XOR2_X1 U573 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  OR2_X1 U574 ( .A1(n532), .A2(n634), .ZN(n525) );
  XOR2_X1 U575 ( .A(KEYINPUT66), .B(n525), .Z(n644) );
  NAND2_X1 U576 ( .A1(G76), .A2(n644), .ZN(n526) );
  XNOR2_X1 U577 ( .A(KEYINPUT73), .B(n526), .ZN(n529) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n639) );
  NAND2_X1 U579 ( .A1(n639), .A2(G89), .ZN(n527) );
  XOR2_X1 U580 ( .A(n527), .B(KEYINPUT4), .Z(n528) );
  NOR2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U582 ( .A(KEYINPUT74), .B(n530), .Z(n531) );
  XNOR2_X1 U583 ( .A(KEYINPUT5), .B(n531), .ZN(n540) );
  XNOR2_X1 U584 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n538) );
  NOR2_X1 U585 ( .A1(G543), .A2(n532), .ZN(n534) );
  XNOR2_X1 U586 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n533) );
  XNOR2_X1 U587 ( .A(n534), .B(n533), .ZN(n640) );
  NAND2_X1 U588 ( .A1(G63), .A2(n640), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G51), .A2(n646), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U591 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U593 ( .A(n541), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U594 ( .A(G168), .B(KEYINPUT8), .Z(n542) );
  XNOR2_X1 U595 ( .A(KEYINPUT76), .B(n542), .ZN(G286) );
  NAND2_X1 U596 ( .A1(G64), .A2(n640), .ZN(n544) );
  NAND2_X1 U597 ( .A1(G52), .A2(n646), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n544), .A2(n543), .ZN(n549) );
  NAND2_X1 U599 ( .A1(G90), .A2(n639), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G77), .A2(n644), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U602 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U603 ( .A1(n549), .A2(n548), .ZN(G171) );
  XOR2_X1 U604 ( .A(KEYINPUT106), .B(G2438), .Z(n551) );
  XNOR2_X1 U605 ( .A(G1341), .B(G2454), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U607 ( .A(n552), .B(G2446), .Z(n554) );
  XNOR2_X1 U608 ( .A(G1348), .B(G2451), .ZN(n553) );
  XNOR2_X1 U609 ( .A(n554), .B(n553), .ZN(n558) );
  XOR2_X1 U610 ( .A(G2430), .B(G2435), .Z(n556) );
  XNOR2_X1 U611 ( .A(G2443), .B(G2427), .ZN(n555) );
  XNOR2_X1 U612 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U613 ( .A(n558), .B(n557), .Z(n559) );
  AND2_X1 U614 ( .A1(G14), .A2(n559), .ZN(G401) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U616 ( .A(G57), .ZN(G237) );
  INV_X1 U617 ( .A(G132), .ZN(G219) );
  INV_X1 U618 ( .A(G82), .ZN(G220) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n560) );
  XNOR2_X1 U620 ( .A(n560), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U621 ( .A(G223), .ZN(n825) );
  NAND2_X1 U622 ( .A1(n825), .A2(G567), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT11), .B(n561), .Z(G234) );
  INV_X1 U624 ( .A(G860), .ZN(n609) );
  NAND2_X1 U625 ( .A1(n639), .A2(G81), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G68), .A2(n644), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U629 ( .A(KEYINPUT13), .B(n565), .ZN(n571) );
  NAND2_X1 U630 ( .A1(G56), .A2(n640), .ZN(n566) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n566), .Z(n569) );
  NAND2_X1 U632 ( .A1(n646), .A2(G43), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT70), .B(n567), .Z(n568) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n992) );
  NOR2_X1 U636 ( .A1(n609), .A2(n992), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(KEYINPUT71), .ZN(G153) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U640 ( .A1(G54), .A2(n646), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G92), .A2(n639), .ZN(n574) );
  NAND2_X1 U642 ( .A1(G66), .A2(n640), .ZN(n573) );
  NAND2_X1 U643 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n644), .A2(G79), .ZN(n575) );
  XOR2_X1 U645 ( .A(KEYINPUT72), .B(n575), .Z(n576) );
  NOR2_X1 U646 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT15), .ZN(n985) );
  OR2_X1 U649 ( .A1(n985), .A2(G868), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U651 ( .A1(G91), .A2(n639), .ZN(n584) );
  NAND2_X1 U652 ( .A1(G53), .A2(n646), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n584), .A2(n583), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G65), .A2(n640), .ZN(n585) );
  XNOR2_X1 U655 ( .A(n585), .B(KEYINPUT68), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G78), .A2(n644), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n991) );
  XNOR2_X1 U659 ( .A(n991), .B(KEYINPUT69), .ZN(G299) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n590) );
  XOR2_X1 U661 ( .A(KEYINPUT77), .B(n590), .Z(n592) );
  INV_X1 U662 ( .A(G868), .ZN(n660) );
  NOR2_X1 U663 ( .A1(G286), .A2(n660), .ZN(n591) );
  NOR2_X1 U664 ( .A1(n592), .A2(n591), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n609), .A2(G559), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n593), .A2(n985), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U668 ( .A1(G868), .A2(n992), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G868), .A2(n985), .ZN(n595) );
  NOR2_X1 U670 ( .A1(G559), .A2(n595), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(G282) );
  NAND2_X1 U672 ( .A1(n870), .A2(G123), .ZN(n598) );
  XNOR2_X1 U673 ( .A(n598), .B(KEYINPUT18), .ZN(n600) );
  NAND2_X1 U674 ( .A1(G135), .A2(n873), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U676 ( .A(KEYINPUT78), .B(n601), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G99), .A2(n875), .ZN(n603) );
  NAND2_X1 U678 ( .A1(G111), .A2(n869), .ZN(n602) );
  NAND2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n968) );
  XOR2_X1 U681 ( .A(n968), .B(G2096), .Z(n606) );
  NOR2_X1 U682 ( .A1(G2100), .A2(n606), .ZN(n607) );
  XNOR2_X1 U683 ( .A(KEYINPUT79), .B(n607), .ZN(G156) );
  NAND2_X1 U684 ( .A1(G559), .A2(n985), .ZN(n608) );
  XOR2_X1 U685 ( .A(n992), .B(n608), .Z(n658) );
  NAND2_X1 U686 ( .A1(n609), .A2(n658), .ZN(n617) );
  NAND2_X1 U687 ( .A1(n640), .A2(G67), .ZN(n611) );
  NAND2_X1 U688 ( .A1(G80), .A2(n644), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n639), .A2(G93), .ZN(n612) );
  XOR2_X1 U691 ( .A(KEYINPUT80), .B(n612), .Z(n613) );
  NOR2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n646), .A2(G55), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n661) );
  XNOR2_X1 U695 ( .A(n617), .B(n661), .ZN(G145) );
  AND2_X1 U696 ( .A1(G72), .A2(n644), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G85), .A2(n639), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G60), .A2(n640), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n646), .A2(G47), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(G290) );
  NAND2_X1 U703 ( .A1(G88), .A2(n639), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G75), .A2(n644), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G62), .A2(n640), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G50), .A2(n646), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U710 ( .A(KEYINPUT85), .B(n630), .Z(G166) );
  NAND2_X1 U711 ( .A1(G49), .A2(n646), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U714 ( .A(KEYINPUT81), .B(n633), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G87), .A2(n634), .ZN(n635) );
  XOR2_X1 U716 ( .A(KEYINPUT82), .B(n635), .Z(n636) );
  NOR2_X1 U717 ( .A1(n640), .A2(n636), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(G288) );
  NAND2_X1 U719 ( .A1(G86), .A2(n639), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G61), .A2(n640), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U722 ( .A(KEYINPUT83), .B(n643), .ZN(n651) );
  NAND2_X1 U723 ( .A1(n644), .A2(G73), .ZN(n645) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n645), .Z(n649) );
  NAND2_X1 U725 ( .A1(n646), .A2(G48), .ZN(n647) );
  XOR2_X1 U726 ( .A(KEYINPUT84), .B(n647), .Z(n648) );
  NOR2_X1 U727 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n651), .A2(n650), .ZN(G305) );
  XNOR2_X1 U729 ( .A(KEYINPUT86), .B(KEYINPUT19), .ZN(n653) );
  XNOR2_X1 U730 ( .A(G290), .B(G166), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(G288), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n655), .B(n661), .ZN(n656) );
  XNOR2_X1 U734 ( .A(n656), .B(G305), .ZN(n657) );
  XNOR2_X1 U735 ( .A(n657), .B(G299), .ZN(n893) );
  XOR2_X1 U736 ( .A(n893), .B(n658), .Z(n659) );
  NOR2_X1 U737 ( .A1(n660), .A2(n659), .ZN(n663) );
  NOR2_X1 U738 ( .A1(G868), .A2(n661), .ZN(n662) );
  NOR2_X1 U739 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2084), .A2(G2078), .ZN(n664) );
  XNOR2_X1 U741 ( .A(n664), .B(KEYINPUT20), .ZN(n665) );
  XNOR2_X1 U742 ( .A(KEYINPUT87), .B(n665), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n666), .A2(G2090), .ZN(n667) );
  XNOR2_X1 U744 ( .A(n667), .B(KEYINPUT88), .ZN(n668) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n670) );
  XNOR2_X1 U749 ( .A(KEYINPUT22), .B(n670), .ZN(n671) );
  NAND2_X1 U750 ( .A1(n671), .A2(G96), .ZN(n672) );
  NOR2_X1 U751 ( .A1(n672), .A2(G218), .ZN(n673) );
  XNOR2_X1 U752 ( .A(n673), .B(KEYINPUT89), .ZN(n1013) );
  NAND2_X1 U753 ( .A1(n1013), .A2(G2106), .ZN(n677) );
  NAND2_X1 U754 ( .A1(G108), .A2(G120), .ZN(n674) );
  NOR2_X1 U755 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U756 ( .A1(G69), .A2(n675), .ZN(n1014) );
  NAND2_X1 U757 ( .A1(n1014), .A2(G567), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n677), .A2(n676), .ZN(n829) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n678) );
  XNOR2_X1 U760 ( .A(KEYINPUT90), .B(n678), .ZN(n679) );
  NOR2_X1 U761 ( .A1(n829), .A2(n679), .ZN(n828) );
  NAND2_X1 U762 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U763 ( .A1(n873), .A2(G138), .ZN(n682) );
  NAND2_X1 U764 ( .A1(G102), .A2(n875), .ZN(n680) );
  XOR2_X1 U765 ( .A(KEYINPUT91), .B(n680), .Z(n681) );
  NAND2_X1 U766 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U767 ( .A1(G114), .A2(n869), .ZN(n684) );
  NAND2_X1 U768 ( .A1(G126), .A2(n870), .ZN(n683) );
  NAND2_X1 U769 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U770 ( .A1(n686), .A2(n685), .ZN(G164) );
  INV_X1 U771 ( .A(G166), .ZN(G303) );
  NAND2_X1 U772 ( .A1(n687), .A2(G40), .ZN(n776) );
  INV_X1 U773 ( .A(n776), .ZN(n688) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n777) );
  NAND2_X1 U775 ( .A1(n688), .A2(n777), .ZN(n689) );
  INV_X1 U776 ( .A(n692), .ZN(n712) );
  XNOR2_X1 U777 ( .A(G2078), .B(KEYINPUT25), .ZN(n905) );
  NAND2_X1 U778 ( .A1(n712), .A2(n905), .ZN(n691) );
  OR2_X1 U779 ( .A1(n712), .A2(G1961), .ZN(n690) );
  NAND2_X1 U780 ( .A1(n691), .A2(n690), .ZN(n725) );
  NOR2_X1 U781 ( .A1(G171), .A2(n725), .ZN(n697) );
  NAND2_X1 U782 ( .A1(n692), .A2(G8), .ZN(n771) );
  NOR2_X1 U783 ( .A1(n730), .A2(G2084), .ZN(n740) );
  NOR2_X1 U784 ( .A1(n741), .A2(n740), .ZN(n693) );
  NAND2_X1 U785 ( .A1(G8), .A2(n693), .ZN(n694) );
  XNOR2_X1 U786 ( .A(KEYINPUT30), .B(n694), .ZN(n695) );
  NOR2_X1 U787 ( .A1(G168), .A2(n695), .ZN(n696) );
  XOR2_X1 U788 ( .A(KEYINPUT31), .B(n698), .Z(n729) );
  NAND2_X1 U789 ( .A1(n712), .A2(G1996), .ZN(n699) );
  XNOR2_X1 U790 ( .A(n699), .B(KEYINPUT26), .ZN(n703) );
  NAND2_X1 U791 ( .A1(n730), .A2(G1341), .ZN(n701) );
  INV_X1 U792 ( .A(n992), .ZN(n700) );
  AND2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n702) );
  AND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n704) );
  OR2_X1 U795 ( .A1(n704), .A2(n985), .ZN(n711) );
  NAND2_X1 U796 ( .A1(n985), .A2(n704), .ZN(n709) );
  AND2_X1 U797 ( .A1(n730), .A2(G1348), .ZN(n705) );
  XNOR2_X1 U798 ( .A(n705), .B(KEYINPUT99), .ZN(n707) );
  NAND2_X1 U799 ( .A1(n712), .A2(G2067), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n717) );
  NAND2_X1 U803 ( .A1(G2072), .A2(n712), .ZN(n713) );
  XNOR2_X1 U804 ( .A(n713), .B(KEYINPUT27), .ZN(n715) );
  INV_X1 U805 ( .A(G1956), .ZN(n936) );
  NOR2_X1 U806 ( .A1(n712), .A2(n936), .ZN(n714) );
  NOR2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U808 ( .A1(n991), .A2(n718), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n722) );
  NOR2_X1 U810 ( .A1(n991), .A2(n718), .ZN(n720) );
  XNOR2_X1 U811 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n724) );
  XOR2_X1 U813 ( .A(KEYINPUT100), .B(KEYINPUT29), .Z(n723) );
  XNOR2_X1 U814 ( .A(n724), .B(n723), .ZN(n727) );
  NAND2_X1 U815 ( .A1(n725), .A2(G171), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U817 ( .A1(n729), .A2(n728), .ZN(n739) );
  NAND2_X1 U818 ( .A1(n739), .A2(G286), .ZN(n735) );
  NOR2_X1 U819 ( .A1(n730), .A2(G2090), .ZN(n732) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n771), .ZN(n731) );
  NOR2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U822 ( .A1(n733), .A2(G303), .ZN(n734) );
  NAND2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U824 ( .A1(n736), .A2(G8), .ZN(n738) );
  XOR2_X1 U825 ( .A(KEYINPUT32), .B(KEYINPUT102), .Z(n737) );
  XNOR2_X1 U826 ( .A(n738), .B(n737), .ZN(n747) );
  XNOR2_X1 U827 ( .A(KEYINPUT101), .B(n739), .ZN(n745) );
  NAND2_X1 U828 ( .A1(n740), .A2(G8), .ZN(n743) );
  INV_X1 U829 ( .A(n741), .ZN(n742) );
  NAND2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U832 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U833 ( .A(n748), .B(KEYINPUT103), .ZN(n764) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U836 ( .A1(n756), .A2(n749), .ZN(n998) );
  INV_X1 U837 ( .A(KEYINPUT33), .ZN(n750) );
  AND2_X1 U838 ( .A1(n998), .A2(n750), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n764), .A2(n751), .ZN(n754) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n997) );
  INV_X1 U841 ( .A(n997), .ZN(n752) );
  OR2_X1 U842 ( .A1(KEYINPUT33), .A2(n515), .ZN(n753) );
  NAND2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n761) );
  XOR2_X1 U844 ( .A(G1981), .B(KEYINPUT104), .Z(n755) );
  XNOR2_X1 U845 ( .A(G305), .B(n755), .ZN(n988) );
  INV_X1 U846 ( .A(n988), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n757), .A2(n771), .ZN(n758) );
  OR2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U851 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n765), .A2(n771), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U855 ( .A(n768), .B(KEYINPUT105), .ZN(n775) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XNOR2_X1 U857 ( .A(n769), .B(KEYINPUT24), .ZN(n770) );
  XNOR2_X1 U858 ( .A(n770), .B(KEYINPUT98), .ZN(n773) );
  INV_X1 U859 ( .A(n771), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n810) );
  NOR2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n820) );
  XNOR2_X1 U863 ( .A(G1991), .B(KEYINPUT94), .ZN(n904) );
  NAND2_X1 U864 ( .A1(G131), .A2(n873), .ZN(n779) );
  NAND2_X1 U865 ( .A1(G119), .A2(n870), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n783) );
  NAND2_X1 U867 ( .A1(G95), .A2(n875), .ZN(n781) );
  NAND2_X1 U868 ( .A1(G107), .A2(n869), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n782) );
  OR2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n881) );
  NAND2_X1 U871 ( .A1(n904), .A2(n881), .ZN(n794) );
  NAND2_X1 U872 ( .A1(n875), .A2(G105), .ZN(n785) );
  XNOR2_X1 U873 ( .A(KEYINPUT38), .B(KEYINPUT96), .ZN(n784) );
  XNOR2_X1 U874 ( .A(n785), .B(n784), .ZN(n792) );
  NAND2_X1 U875 ( .A1(G141), .A2(n873), .ZN(n787) );
  NAND2_X1 U876 ( .A1(G129), .A2(n870), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U878 ( .A1(G117), .A2(n869), .ZN(n788) );
  XNOR2_X1 U879 ( .A(KEYINPUT95), .B(n788), .ZN(n789) );
  NOR2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n886) );
  NAND2_X1 U882 ( .A1(G1996), .A2(n886), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n969) );
  AND2_X1 U884 ( .A1(n820), .A2(n969), .ZN(n813) );
  XNOR2_X1 U885 ( .A(KEYINPUT97), .B(n813), .ZN(n797) );
  XNOR2_X1 U886 ( .A(G1986), .B(G290), .ZN(n994) );
  NAND2_X1 U887 ( .A1(n994), .A2(n820), .ZN(n795) );
  XNOR2_X1 U888 ( .A(n795), .B(KEYINPUT92), .ZN(n796) );
  AND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n808) );
  NAND2_X1 U890 ( .A1(G104), .A2(n875), .ZN(n799) );
  NAND2_X1 U891 ( .A1(G140), .A2(n873), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U893 ( .A(KEYINPUT34), .B(n800), .ZN(n805) );
  NAND2_X1 U894 ( .A1(G116), .A2(n869), .ZN(n802) );
  NAND2_X1 U895 ( .A1(G128), .A2(n870), .ZN(n801) );
  NAND2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U897 ( .A(KEYINPUT35), .B(n803), .Z(n804) );
  NOR2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U899 ( .A(KEYINPUT36), .B(n806), .ZN(n867) );
  XOR2_X1 U900 ( .A(G2067), .B(KEYINPUT37), .Z(n807) );
  XNOR2_X1 U901 ( .A(KEYINPUT93), .B(n807), .ZN(n818) );
  NOR2_X1 U902 ( .A1(n867), .A2(n818), .ZN(n978) );
  NAND2_X1 U903 ( .A1(n820), .A2(n978), .ZN(n816) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n823) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n886), .ZN(n959) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n881), .A2(n904), .ZN(n970) );
  NOR2_X1 U908 ( .A1(n811), .A2(n970), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n959), .A2(n814), .ZN(n815) );
  XNOR2_X1 U911 ( .A(KEYINPUT39), .B(n815), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n867), .A2(n818), .ZN(n965) );
  NAND2_X1 U914 ( .A1(n819), .A2(n965), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U917 ( .A(n824), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n825), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U920 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(G188) );
  XNOR2_X1 U923 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  INV_X1 U924 ( .A(n829), .ZN(G319) );
  XOR2_X1 U925 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n831) );
  XNOR2_X1 U926 ( .A(KEYINPUT110), .B(G2678), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U928 ( .A(n832), .B(G2100), .Z(n834) );
  XNOR2_X1 U929 ( .A(G2072), .B(G2084), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U931 ( .A(KEYINPUT43), .B(G2096), .Z(n836) );
  XNOR2_X1 U932 ( .A(G2090), .B(KEYINPUT109), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U934 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2078), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(G227) );
  XOR2_X1 U937 ( .A(G1966), .B(G1956), .Z(n842) );
  XNOR2_X1 U938 ( .A(G1971), .B(G1961), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U940 ( .A(n843), .B(G2474), .Z(n845) );
  XNOR2_X1 U941 ( .A(G1981), .B(G1976), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U943 ( .A(KEYINPUT41), .B(G1986), .Z(n847) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(G229) );
  NAND2_X1 U947 ( .A1(G112), .A2(n869), .ZN(n856) );
  NAND2_X1 U948 ( .A1(G100), .A2(n875), .ZN(n851) );
  NAND2_X1 U949 ( .A1(G136), .A2(n873), .ZN(n850) );
  NAND2_X1 U950 ( .A1(n851), .A2(n850), .ZN(n854) );
  NAND2_X1 U951 ( .A1(n870), .A2(G124), .ZN(n852) );
  XOR2_X1 U952 ( .A(KEYINPUT44), .B(n852), .Z(n853) );
  NOR2_X1 U953 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n857), .B(KEYINPUT111), .ZN(G162) );
  NAND2_X1 U956 ( .A1(G103), .A2(n875), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G139), .A2(n873), .ZN(n858) );
  NAND2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n865) );
  NAND2_X1 U959 ( .A1(G115), .A2(n869), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G127), .A2(n870), .ZN(n860) );
  NAND2_X1 U961 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U962 ( .A(KEYINPUT113), .B(n862), .ZN(n863) );
  XNOR2_X1 U963 ( .A(KEYINPUT47), .B(n863), .ZN(n864) );
  NOR2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n961) );
  XNOR2_X1 U965 ( .A(G164), .B(n961), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n866), .B(n968), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n891) );
  NAND2_X1 U968 ( .A1(G118), .A2(n869), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G130), .A2(n870), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n880) );
  NAND2_X1 U971 ( .A1(n873), .A2(G142), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n874), .B(KEYINPUT112), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G106), .A2(n875), .ZN(n876) );
  NAND2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U975 ( .A(KEYINPUT45), .B(n878), .Z(n879) );
  NOR2_X1 U976 ( .A1(n880), .A2(n879), .ZN(n885) );
  XNOR2_X1 U977 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n883) );
  XNOR2_X1 U978 ( .A(n881), .B(KEYINPUT114), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U980 ( .A(n885), .B(n884), .ZN(n889) );
  XNOR2_X1 U981 ( .A(G160), .B(G162), .ZN(n887) );
  XNOR2_X1 U982 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U983 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U984 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U985 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U986 ( .A(n992), .B(n893), .ZN(n895) );
  XNOR2_X1 U987 ( .A(G171), .B(n985), .ZN(n894) );
  XNOR2_X1 U988 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U989 ( .A(n896), .B(G286), .Z(n897) );
  NOR2_X1 U990 ( .A1(G37), .A2(n897), .ZN(G397) );
  NOR2_X1 U991 ( .A1(G227), .A2(G229), .ZN(n898) );
  XNOR2_X1 U992 ( .A(n898), .B(KEYINPUT49), .ZN(n899) );
  NOR2_X1 U993 ( .A1(G401), .A2(n899), .ZN(n900) );
  NAND2_X1 U994 ( .A1(G319), .A2(n900), .ZN(n901) );
  XNOR2_X1 U995 ( .A(KEYINPUT115), .B(n901), .ZN(n903) );
  NOR2_X1 U996 ( .A1(G395), .A2(G397), .ZN(n902) );
  NAND2_X1 U997 ( .A1(n903), .A2(n902), .ZN(G225) );
  XOR2_X1 U998 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  XOR2_X1 U1000 ( .A(n904), .B(G25), .Z(n911) );
  XNOR2_X1 U1001 ( .A(G27), .B(KEYINPUT119), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(G32), .B(G1996), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(KEYINPUT120), .B(n909), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(n918) );
  XOR2_X1 U1007 ( .A(G2067), .B(G26), .Z(n912) );
  XNOR2_X1 U1008 ( .A(KEYINPUT117), .B(n912), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(G33), .B(G2072), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(KEYINPUT118), .B(n915), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n916), .A2(G28), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1014 ( .A(KEYINPUT53), .B(n919), .Z(n923) );
  XNOR2_X1 U1015 ( .A(KEYINPUT54), .B(G34), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(n920), .B(KEYINPUT121), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(G2084), .B(n921), .ZN(n922) );
  NAND2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n925) );
  XNOR2_X1 U1019 ( .A(G35), .B(G2090), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(KEYINPUT55), .B(n926), .ZN(n928) );
  INV_X1 U1022 ( .A(G29), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n929), .A2(G11), .ZN(n930) );
  XNOR2_X1 U1025 ( .A(n930), .B(KEYINPUT122), .ZN(n957) );
  XNOR2_X1 U1026 ( .A(G1961), .B(G5), .ZN(n945) );
  XNOR2_X1 U1027 ( .A(G1348), .B(KEYINPUT59), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n931), .B(G4), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(G1981), .B(G6), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(G19), .B(G1341), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n939) );
  XOR2_X1 U1033 ( .A(KEYINPUT124), .B(n936), .Z(n937) );
  XNOR2_X1 U1034 ( .A(G20), .B(n937), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1036 ( .A(KEYINPUT60), .B(n940), .Z(n942) );
  XNOR2_X1 U1037 ( .A(G1966), .B(G21), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(KEYINPUT125), .B(n943), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n953) );
  XOR2_X1 U1041 ( .A(G1986), .B(KEYINPUT126), .Z(n946) );
  XNOR2_X1 U1042 ( .A(G24), .B(n946), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(G1976), .B(G23), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G1971), .B(G22), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1047 ( .A(KEYINPUT58), .B(n951), .Z(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(KEYINPUT61), .B(n954), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n955), .A2(G16), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n984) );
  XOR2_X1 U1052 ( .A(G2090), .B(G162), .Z(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1054 ( .A(KEYINPUT51), .B(n960), .Z(n976) );
  XOR2_X1 U1055 ( .A(G2072), .B(n961), .Z(n963) );
  XOR2_X1 U1056 ( .A(G164), .B(G2078), .Z(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n964), .B(KEYINPUT50), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n974) );
  XOR2_X1 U1060 ( .A(G2084), .B(G160), .Z(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n972) );
  NOR2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1066 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(KEYINPUT52), .B(n979), .ZN(n981) );
  INV_X1 U1068 ( .A(KEYINPUT55), .ZN(n980) );
  NAND2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1070 ( .A1(n982), .A2(G29), .ZN(n983) );
  NAND2_X1 U1071 ( .A1(n984), .A2(n983), .ZN(n1011) );
  XOR2_X1 U1072 ( .A(KEYINPUT56), .B(G16), .Z(n1009) );
  XNOR2_X1 U1073 ( .A(n985), .B(G1348), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(G171), .B(G1961), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n1007) );
  XNOR2_X1 U1076 ( .A(G168), .B(G1966), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(n990), .B(KEYINPUT57), .ZN(n1005) );
  XNOR2_X1 U1079 ( .A(n991), .B(G1956), .ZN(n996) );
  XNOR2_X1 U1080 ( .A(G1341), .B(n992), .ZN(n993) );
  NOR2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1082 ( .A1(n996), .A2(n995), .ZN(n1003) );
  AND2_X1 U1083 ( .A1(G303), .A2(G1971), .ZN(n1000) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(KEYINPUT123), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1087 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1088 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1089 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1090 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1091 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1092 ( .A(KEYINPUT62), .B(n1012), .ZN(G311) );
  XNOR2_X1 U1093 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1094 ( .A(G108), .ZN(G238) );
  INV_X1 U1095 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1096 ( .A1(n1014), .A2(n1013), .ZN(G325) );
  INV_X1 U1097 ( .A(G325), .ZN(G261) );
  INV_X1 U1098 ( .A(G69), .ZN(G235) );
endmodule

