//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT23), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT66), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n215), .A2(new_n216), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n210), .A2(KEYINPUT25), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(new_n211), .A3(new_n212), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n214), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n220), .A2(new_n222), .B1(new_n223), .B2(KEYINPUT64), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n216), .A2(new_n225), .A3(new_n214), .ZN(new_n226));
  NAND3_X1  g025(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n209), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n219), .B1(new_n229), .B2(KEYINPUT25), .ZN(new_n230));
  INV_X1    g029(.A(G120gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G113gat), .ZN(new_n232));
  INV_X1    g031(.A(G113gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G120gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n236));
  INV_X1    g035(.A(G134gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G127gat), .ZN(new_n238));
  INV_X1    g037(.A(G127gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G134gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n235), .A2(new_n236), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(new_n240), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(KEYINPUT1), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n248), .B(new_n212), .C1(new_n211), .C2(KEYINPUT27), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT28), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n212), .B1(new_n211), .B2(KEYINPUT27), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT27), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n252), .A2(G183gat), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n249), .B(new_n250), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(G190gat), .B1(new_n252), .B2(G183gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n255), .B(new_n256), .C1(new_n248), .C2(KEYINPUT28), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n203), .A2(new_n204), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT26), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n259), .A2(new_n260), .A3(new_n208), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n216), .B1(new_n259), .B2(new_n260), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n258), .A2(KEYINPUT68), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT68), .B1(new_n258), .B2(new_n263), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n230), .B(new_n247), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n258), .A2(new_n263), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n258), .A2(KEYINPUT68), .A3(new_n263), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n222), .A2(new_n220), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n223), .A2(KEYINPUT64), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n226), .A2(new_n227), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n210), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT25), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n269), .A2(new_n270), .B1(new_n277), .B2(new_n219), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n245), .B(KEYINPUT69), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n266), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G227gat), .A2(G233gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT32), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT33), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G15gat), .B(G43gat), .Z(new_n287));
  XNOR2_X1  g086(.A(G71gat), .B(G99gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n281), .B(new_n266), .C1(new_n278), .C2(new_n279), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT34), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n289), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n283), .B(KEYINPUT32), .C1(new_n285), .C2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n290), .A2(new_n298), .A3(new_n293), .A4(new_n295), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n293), .B1(new_n290), .B2(new_n295), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n202), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  AOI211_X1 g102(.A(KEYINPUT83), .B(new_n301), .C1(new_n297), .C2(new_n299), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G141gat), .B(G148gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(G155gat), .B2(G162gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n308), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G141gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G148gat), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G141gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G155gat), .B(G162gat), .ZN(new_n318));
  INV_X1    g117(.A(G155gat), .ZN(new_n319));
  INV_X1    g118(.A(G162gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT2), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n312), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n324), .A2(new_n245), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n312), .A2(new_n322), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT73), .B1(new_n326), .B2(KEYINPUT3), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n328));
  AOI211_X1 g127(.A(new_n328), .B(new_n323), .C1(new_n312), .C2(new_n322), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n325), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n331));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n312), .A2(new_n322), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT4), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n334), .A2(new_n335), .A3(new_n241), .A4(new_n244), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n241), .A2(new_n244), .A3(new_n312), .A4(new_n322), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(KEYINPUT77), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n337), .A2(new_n340), .A3(KEYINPUT4), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n333), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n245), .A2(new_n326), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n337), .ZN(new_n346));
  INV_X1    g145(.A(new_n332), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT74), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n349));
  AOI211_X1 g148(.A(new_n349), .B(new_n332), .C1(new_n345), .C2(new_n337), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT5), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n338), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n330), .A2(new_n352), .A3(new_n332), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n344), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n337), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n241), .A2(new_n244), .B1(new_n312), .B2(new_n322), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n347), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n349), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n346), .A2(KEYINPUT74), .A3(new_n347), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n330), .A2(new_n352), .A3(new_n332), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n360), .A2(KEYINPUT75), .A3(KEYINPUT5), .A4(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n343), .B1(new_n354), .B2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(G1gat), .B(G29gat), .Z(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G57gat), .B(G85gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT6), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT6), .ZN(new_n371));
  INV_X1    g170(.A(new_n343), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n351), .A2(new_n353), .A3(new_n344), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n331), .B1(new_n358), .B2(new_n359), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT75), .B1(new_n374), .B2(new_n361), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n372), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n368), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n371), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n370), .B1(new_n378), .B2(new_n369), .ZN(new_n379));
  NAND2_X1  g178(.A1(G228gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT29), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n324), .A2(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(G211gat), .A2(G218gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(G211gat), .A2(G218gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(G197gat), .A2(G204gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(G197gat), .A2(G204gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G211gat), .B(G218gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G197gat), .B(G204gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n390), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n383), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n396), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT3), .B1(new_n398), .B2(new_n382), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n381), .B(new_n397), .C1(new_n399), .C2(new_n334), .ZN(new_n400));
  INV_X1    g199(.A(new_n397), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT80), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n391), .A2(new_n395), .A3(KEYINPUT79), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n392), .A2(new_n393), .A3(new_n404), .A4(new_n394), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n382), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n402), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n405), .A2(new_n382), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n395), .A3(KEYINPUT79), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT80), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n323), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n401), .B1(new_n411), .B2(new_n326), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n400), .B1(new_n412), .B2(new_n381), .ZN(new_n413));
  INV_X1    g212(.A(G22gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT31), .B(G50gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  NAND2_X1  g218(.A1(new_n410), .A2(new_n323), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT80), .B1(new_n408), .B2(new_n409), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n326), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n397), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n380), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n414), .B1(new_n424), .B2(new_n400), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT81), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n416), .B(new_n419), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n426), .B1(new_n413), .B2(G22gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n419), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT82), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n415), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n427), .A2(new_n430), .A3(new_n415), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n230), .A2(new_n267), .ZN(new_n434));
  INV_X1    g233(.A(G226gat), .ZN(new_n435));
  INV_X1    g234(.A(G233gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(KEYINPUT29), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n230), .B1(new_n264), .B2(new_n265), .ZN(new_n440));
  INV_X1    g239(.A(new_n437), .ZN(new_n441));
  OAI22_X1  g240(.A1(new_n434), .A2(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n398), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n230), .A2(new_n267), .A3(new_n437), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n396), .B(new_n444), .C1(new_n278), .C2(new_n439), .ZN(new_n445));
  XNOR2_X1  g244(.A(G8gat), .B(G36gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(G64gat), .B(G92gat), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n446), .B(new_n447), .Z(new_n448));
  NAND3_X1  g247(.A1(new_n443), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n449), .A2(KEYINPUT30), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(KEYINPUT30), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n443), .A2(new_n445), .ZN(new_n452));
  INV_X1    g251(.A(new_n448), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT72), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT72), .ZN(new_n455));
  AOI211_X1 g254(.A(new_n455), .B(new_n448), .C1(new_n443), .C2(new_n445), .ZN(new_n456));
  OAI22_X1  g255(.A1(new_n450), .A2(new_n451), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n458));
  AND4_X1   g257(.A1(new_n379), .A2(new_n432), .A3(new_n433), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n305), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n427), .A2(new_n430), .A3(new_n415), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n431), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n376), .A2(new_n463), .A3(new_n377), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT78), .B1(new_n363), .B2(new_n368), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT6), .B1(new_n363), .B2(new_n368), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n457), .B1(new_n467), .B2(new_n370), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n290), .A2(KEYINPUT70), .A3(new_n295), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n290), .A2(new_n295), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT70), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n293), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n469), .A2(new_n472), .B1(new_n297), .B2(new_n299), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n462), .A2(new_n468), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT35), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n339), .A2(new_n330), .A3(new_n341), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n347), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n368), .B1(new_n478), .B2(KEYINPUT39), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT39), .B1(new_n346), .B2(new_n347), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n477), .B2(new_n347), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n376), .A2(new_n377), .B1(new_n482), .B2(KEYINPUT40), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n482), .A2(KEYINPUT40), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n457), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT38), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n442), .A2(new_n396), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n398), .B(new_n444), .C1(new_n278), .C2(new_n439), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(KEYINPUT37), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n448), .B1(new_n443), .B2(new_n445), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n453), .A2(KEYINPUT37), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n486), .B(new_n489), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n452), .A2(new_n453), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n494), .A2(new_n491), .B1(KEYINPUT37), .B2(new_n452), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n449), .B(new_n493), .C1(new_n495), .C2(new_n486), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n485), .B1(new_n379), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n462), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n432), .A2(new_n433), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n468), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n300), .A2(new_n502), .A3(new_n302), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n473), .B2(new_n502), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n476), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G190gat), .B(G218gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT41), .ZN(new_n510));
  INV_X1    g309(.A(G232gat), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n510), .A2(new_n511), .A3(new_n436), .ZN(new_n512));
  INV_X1    g311(.A(G29gat), .ZN(new_n513));
  INV_X1    g312(.A(G36gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT14), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT14), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(G29gat), .A2(G36gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n520));
  INV_X1    g319(.A(G43gat), .ZN(new_n521));
  INV_X1    g320(.A(G50gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G43gat), .A2(G50gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT85), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n523), .A2(new_n524), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(KEYINPUT15), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n523), .A2(KEYINPUT86), .A3(new_n520), .A4(new_n524), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539));
  INV_X1    g338(.A(G85gat), .ZN(new_n540));
  INV_X1    g339(.A(G92gat), .ZN(new_n541));
  AOI22_X1  g340(.A1(KEYINPUT8), .A2(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G99gat), .B(G106gat), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n544), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(new_n538), .A3(new_n542), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n512), .B1(new_n536), .B2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n548), .B(KEYINPUT93), .Z(new_n551));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT85), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n526), .B(new_n553), .ZN(new_n554));
  AOI211_X1 g353(.A(new_n525), .B(new_n519), .C1(new_n530), .C2(new_n531), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n527), .A2(new_n535), .A3(KEYINPUT17), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n509), .B(new_n550), .C1(new_n551), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT94), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT92), .B(G134gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G162gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n510), .B1(new_n511), .B2(new_n436), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n550), .B1(new_n551), .B2(new_n558), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n508), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n559), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT87), .ZN(new_n571));
  INV_X1    g370(.A(G1gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(KEYINPUT87), .A3(G1gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT16), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(G8gat), .ZN(new_n578));
  INV_X1    g377(.A(G8gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n571), .A2(new_n572), .B1(new_n575), .B2(new_n570), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(new_n574), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT21), .ZN(new_n584));
  XOR2_X1   g383(.A(G71gat), .B(G78gat), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  INV_X1    g386(.A(G71gat), .ZN(new_n588));
  INV_X1    g387(.A(G78gat), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G57gat), .B(G64gat), .Z(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n590), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n585), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n577), .B(G8gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n595), .A2(new_n584), .ZN(new_n598));
  OAI21_X1  g397(.A(KEYINPUT91), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G127gat), .B(G155gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT20), .ZN(new_n602));
  INV_X1    g401(.A(G231gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(new_n436), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n595), .B2(new_n584), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n595), .A2(new_n584), .A3(new_n605), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n602), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n607), .A2(new_n602), .A3(new_n608), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n600), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n599), .B(new_n596), .C1(new_n613), .C2(new_n609), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n612), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n617), .B1(new_n612), .B2(new_n614), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n548), .A2(new_n595), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n545), .A2(new_n547), .A3(new_n594), .A4(new_n592), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n623), .A2(new_n622), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT95), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n621), .A2(new_n623), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n632), .A2(KEYINPUT96), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n632), .A2(KEYINPUT96), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n639), .A2(new_n630), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n565), .A2(new_n568), .ZN(new_n644));
  AND4_X1   g443(.A1(new_n569), .A2(new_n620), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n556), .A2(new_n582), .A3(new_n557), .ZN(new_n646));
  NAND2_X1  g445(.A1(G229gat), .A2(G233gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n597), .A2(new_n536), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT88), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT18), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT18), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(KEYINPUT88), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n597), .B(new_n536), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n647), .B(KEYINPUT13), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G113gat), .B(G141gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT84), .B(G197gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT11), .B(G169gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT12), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n651), .A2(new_n653), .A3(new_n656), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT89), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n650), .A2(KEYINPUT18), .B1(new_n654), .B2(new_n655), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT89), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n665), .A2(new_n666), .A3(new_n653), .A4(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n653), .ZN(new_n669));
  INV_X1    g468(.A(new_n662), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n645), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n507), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n467), .A2(new_n370), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n572), .ZN(G1324gat));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n678));
  INV_X1    g477(.A(new_n674), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n457), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT97), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n679), .A2(new_n457), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT98), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n686), .A3(G8gat), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n686), .B1(new_n685), .B2(G8gat), .ZN(new_n689));
  OAI22_X1  g488(.A1(new_n688), .A2(new_n689), .B1(new_n682), .B2(new_n681), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n678), .B1(new_n684), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT97), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n683), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n681), .A2(new_n682), .ZN(new_n694));
  INV_X1    g493(.A(new_n689), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n687), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n696), .A3(KEYINPUT99), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n691), .A2(new_n697), .ZN(G1325gat));
  NAND2_X1  g497(.A1(new_n470), .A2(new_n471), .ZN(new_n699));
  INV_X1    g498(.A(new_n293), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n700), .A3(new_n469), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n502), .B1(new_n300), .B2(new_n701), .ZN(new_n702));
  AOI211_X1 g501(.A(KEYINPUT36), .B(new_n301), .C1(new_n297), .C2(new_n299), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT100), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT100), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n503), .B(new_n705), .C1(new_n473), .C2(new_n502), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(G15gat), .B1(new_n674), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n305), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(G15gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n674), .B2(new_n712), .ZN(G1326gat));
  NOR2_X1   g512(.A1(new_n674), .A2(new_n462), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  AOI22_X1  g515(.A1(new_n664), .A2(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n717), .A2(new_n620), .A3(new_n642), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n707), .A2(new_n501), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(new_n476), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n704), .A2(new_n706), .B1(new_n498), .B2(new_n500), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n305), .A2(new_n459), .B1(new_n474), .B2(KEYINPUT35), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT102), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n569), .A2(new_n644), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(KEYINPUT44), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n722), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n504), .B1(new_n498), .B2(new_n500), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n731), .B2(new_n727), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n719), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G29gat), .B1(new_n734), .B2(new_n675), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n726), .B(new_n718), .C1(new_n724), .C2(new_n730), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n675), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n737), .A2(new_n513), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT45), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n735), .A2(new_n740), .ZN(G1328gat));
  INV_X1    g540(.A(new_n457), .ZN(new_n742));
  OAI21_X1  g541(.A(G36gat), .B1(new_n734), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n736), .A2(G36gat), .A3(new_n742), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT46), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(G1329gat));
  NOR2_X1   g545(.A1(new_n711), .A2(G43gat), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT103), .B1(new_n736), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n727), .B1(new_n476), .B2(new_n506), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n750), .A2(new_n751), .A3(new_n718), .A4(new_n747), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT47), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  AOI211_X1 g552(.A(new_n709), .B(new_n719), .C1(new_n729), .C2(new_n732), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(new_n521), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n749), .A2(new_n752), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n729), .A2(new_n732), .ZN(new_n758));
  INV_X1    g557(.A(new_n707), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(new_n759), .A3(new_n718), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n757), .B1(new_n760), .B2(G43gat), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n755), .B(new_n756), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n521), .B1(new_n733), .B2(new_n759), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT47), .B1(new_n765), .B2(new_n757), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n756), .B1(new_n766), .B2(new_n755), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n764), .A2(new_n767), .ZN(G1330gat));
  AOI21_X1  g567(.A(G50gat), .B1(new_n737), .B2(new_n499), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n462), .A2(new_n522), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n733), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT105), .B(KEYINPUT48), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n771), .B(new_n772), .Z(G1331gat));
  INV_X1    g572(.A(new_n620), .ZN(new_n774));
  NOR4_X1   g573(.A1(new_n672), .A2(new_n726), .A3(new_n774), .A4(new_n643), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n722), .A2(new_n725), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n722), .A2(new_n725), .A3(KEYINPUT106), .A4(new_n775), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(new_n738), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G57gat), .ZN(G1332gat));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n742), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n784), .A2(KEYINPUT107), .ZN(new_n785));
  INV_X1    g584(.A(G64gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(KEYINPUT107), .ZN(new_n787));
  AND4_X1   g586(.A1(new_n782), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n785), .A2(new_n787), .B1(new_n782), .B2(new_n786), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(G1333gat));
  NOR2_X1   g589(.A1(new_n709), .A2(new_n588), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n778), .A2(new_n779), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n778), .A2(KEYINPUT108), .A3(new_n779), .A4(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n778), .A2(new_n305), .A3(new_n779), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n588), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT50), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n796), .A2(new_n801), .A3(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1334gat));
  NAND3_X1  g602(.A1(new_n778), .A2(new_n499), .A3(new_n779), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g604(.A(new_n727), .B1(new_n720), .B2(new_n476), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n806), .A2(KEYINPUT109), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n672), .A2(new_n620), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n806), .B2(KEYINPUT109), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n807), .A2(KEYINPUT51), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n815), .A2(new_n540), .A3(new_n738), .A4(new_n642), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n809), .A2(new_n643), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n758), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G85gat), .B1(new_n818), .B2(new_n675), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n819), .ZN(G1336gat));
  INV_X1    g619(.A(new_n818), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n541), .B1(new_n821), .B2(new_n457), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n742), .A2(G92gat), .A3(new_n643), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n813), .B2(new_n814), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  XNOR2_X1  g626(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n823), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n828), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n822), .B2(new_n826), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(G1337gat));
  NOR3_X1   g631(.A1(new_n711), .A2(G99gat), .A3(new_n643), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT111), .Z(new_n834));
  NAND2_X1  g633(.A1(new_n815), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(G99gat), .B1(new_n818), .B2(new_n709), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1338gat));
  INV_X1    g636(.A(G106gat), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n821), .B2(new_n499), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n462), .A2(G106gat), .A3(new_n643), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT112), .Z(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(new_n813), .B2(new_n814), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT53), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n839), .A2(KEYINPUT53), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n815), .A2(new_n840), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(G1339gat));
  INV_X1    g645(.A(KEYINPUT113), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n654), .A2(new_n655), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n647), .B1(new_n646), .B2(new_n648), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n661), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n668), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n624), .A2(new_n625), .A3(new_n628), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n630), .A2(KEYINPUT54), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n628), .B1(new_n624), .B2(new_n625), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n636), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT55), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n853), .A2(KEYINPUT55), .A3(new_n856), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n641), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n861), .B1(new_n569), .B2(new_n644), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n847), .B1(new_n851), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n668), .A2(new_n850), .ZN(new_n864));
  INV_X1    g663(.A(new_n861), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n726), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT113), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n668), .A2(new_n642), .A3(new_n850), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n717), .B2(new_n861), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n727), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n620), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n645), .A2(new_n717), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n462), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n675), .A2(new_n457), .ZN(new_n878));
  OAI211_X1 g677(.A(KEYINPUT114), .B(new_n462), .C1(new_n872), .C2(new_n874), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n877), .A2(new_n305), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n711), .B1(new_n875), .B2(new_n876), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n883), .A2(KEYINPUT115), .A3(new_n878), .A4(new_n879), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n882), .A2(G113gat), .A3(new_n672), .A4(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n872), .A2(new_n874), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n675), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n887), .A2(new_n473), .A3(new_n742), .A4(new_n462), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n233), .B1(new_n888), .B2(new_n717), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n885), .A2(new_n889), .ZN(G1340gat));
  NAND3_X1  g689(.A1(new_n882), .A2(new_n642), .A3(new_n884), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n891), .A2(new_n892), .A3(G120gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n891), .B2(G120gat), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n642), .A2(new_n231), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n893), .A2(new_n894), .B1(new_n888), .B2(new_n895), .ZN(G1341gat));
  AND3_X1   g695(.A1(new_n882), .A2(new_n620), .A3(new_n884), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n620), .A2(new_n239), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n897), .A2(new_n239), .B1(new_n888), .B2(new_n898), .ZN(G1342gat));
  NOR3_X1   g698(.A1(new_n888), .A2(G134gat), .A3(new_n727), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT56), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n882), .A2(new_n726), .A3(new_n884), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n237), .B2(new_n902), .ZN(G1343gat));
  NAND2_X1  g702(.A1(new_n707), .A2(new_n878), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n462), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT55), .B1(new_n857), .B2(KEYINPUT117), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(KEYINPUT117), .B2(new_n857), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n641), .A3(new_n860), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n869), .B1(new_n910), .B2(new_n717), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n727), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n868), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n774), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n907), .B1(new_n914), .B2(new_n873), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n905), .B1(new_n886), .B2(new_n462), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n904), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n313), .B1(new_n918), .B2(new_n672), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n887), .A2(new_n742), .A3(new_n499), .A4(new_n709), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n920), .A2(G141gat), .A3(new_n717), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(G1344gat));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n925));
  INV_X1    g724(.A(new_n918), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n925), .B(G148gat), .C1(new_n926), .C2(new_n643), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n904), .B(KEYINPUT118), .Z(new_n928));
  INV_X1    g727(.A(KEYINPUT119), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n645), .A2(new_n929), .A3(new_n717), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n645), .B2(new_n717), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n864), .A2(new_n866), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n933), .B1(new_n911), .B2(new_n727), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n932), .B1(new_n934), .B2(new_n620), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n462), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n932), .B(KEYINPUT120), .C1(new_n934), .C2(new_n620), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT57), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n886), .A2(new_n907), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n642), .B(new_n928), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G148gat), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT121), .B1(new_n942), .B2(KEYINPUT59), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n944));
  AOI211_X1 g743(.A(new_n944), .B(new_n925), .C1(new_n941), .C2(G148gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n927), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OR3_X1    g745(.A1(new_n920), .A2(G148gat), .A3(new_n643), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1345gat));
  OAI21_X1  g747(.A(G155gat), .B1(new_n926), .B2(new_n774), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n620), .A2(new_n319), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n920), .B2(new_n950), .ZN(G1346gat));
  NAND3_X1  g750(.A1(new_n918), .A2(G162gat), .A3(new_n726), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n320), .B1(new_n920), .B2(new_n727), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n738), .A2(new_n742), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n883), .A2(new_n879), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(G169gat), .B1(new_n957), .B2(new_n717), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n956), .A2(new_n473), .A3(new_n462), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n886), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n203), .A3(new_n672), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n962), .B(new_n963), .ZN(G1348gat));
  OAI21_X1  g763(.A(G176gat), .B1(new_n957), .B2(new_n643), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n960), .A2(new_n204), .A3(new_n642), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1349gat));
  OAI21_X1  g766(.A(G183gat), .B1(new_n957), .B2(new_n774), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n774), .A2(new_n969), .A3(new_n253), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT124), .B1(new_n960), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n883), .A2(new_n726), .A3(new_n879), .A4(new_n956), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n974), .B1(new_n975), .B2(G190gat), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(new_n974), .A3(G190gat), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n976), .A2(new_n977), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n960), .A2(new_n212), .A3(new_n726), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(G1351gat));
  NOR2_X1   g782(.A1(new_n939), .A2(new_n940), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n709), .A2(new_n956), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n984), .A2(new_n986), .A3(new_n717), .ZN(new_n987));
  INV_X1    g786(.A(G197gat), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n886), .A2(new_n462), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n672), .A2(new_n988), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(KEYINPUT126), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT126), .ZN(new_n995));
  OAI221_X1 g794(.A(new_n995), .B1(new_n991), .B2(new_n992), .C1(new_n987), .C2(new_n988), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n996), .ZN(G1352gat));
  NOR3_X1   g796(.A1(new_n991), .A2(G204gat), .A3(new_n643), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n999));
  OR2_X1    g798(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n984), .A2(new_n986), .A3(new_n643), .ZN(new_n1002));
  INV_X1    g801(.A(G204gat), .ZN(new_n1003));
  OAI211_X1 g802(.A(new_n1000), .B(new_n1001), .C1(new_n1002), .C2(new_n1003), .ZN(G1353gat));
  NOR2_X1   g803(.A1(new_n984), .A2(new_n986), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(new_n620), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n1006), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(KEYINPUT63), .B1(new_n1006), .B2(G211gat), .ZN(new_n1008));
  OR2_X1    g807(.A1(new_n774), .A2(G211gat), .ZN(new_n1009));
  OAI22_X1  g808(.A1(new_n1007), .A2(new_n1008), .B1(new_n991), .B2(new_n1009), .ZN(G1354gat));
  INV_X1    g809(.A(G218gat), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1011), .B1(new_n991), .B2(new_n727), .ZN(new_n1012));
  XNOR2_X1  g811(.A(new_n1012), .B(KEYINPUT127), .ZN(new_n1013));
  NOR2_X1   g812(.A1(new_n727), .A2(new_n1011), .ZN(new_n1014));
  AOI21_X1  g813(.A(new_n1013), .B1(new_n1005), .B2(new_n1014), .ZN(G1355gat));
endmodule


