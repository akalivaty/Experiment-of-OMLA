

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U554 ( .A1(n771), .A2(n769), .ZN(n718) );
  OR2_X1 U555 ( .A1(n764), .A2(n753), .ZN(n519) );
  XNOR2_X1 U556 ( .A(n727), .B(KEYINPUT99), .ZN(n728) );
  XNOR2_X1 U557 ( .A(n729), .B(n728), .ZN(n730) );
  INV_X1 U558 ( .A(KEYINPUT101), .ZN(n734) );
  XNOR2_X1 U559 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U560 ( .A(n739), .B(KEYINPUT32), .ZN(n747) );
  NAND2_X1 U561 ( .A1(n519), .A2(n912), .ZN(n755) );
  NOR2_X1 U562 ( .A1(G651), .A2(n645), .ZN(n644) );
  NOR2_X1 U563 ( .A1(G2104), .A2(n540), .ZN(n881) );
  NOR2_X1 U564 ( .A1(n571), .A2(n570), .ZN(n924) );
  XOR2_X1 U565 ( .A(KEYINPUT0), .B(G543), .Z(n645) );
  NAND2_X1 U566 ( .A1(n644), .A2(G51), .ZN(n520) );
  XOR2_X1 U567 ( .A(KEYINPUT77), .B(n520), .Z(n523) );
  INV_X1 U568 ( .A(G651), .ZN(n526) );
  NOR2_X1 U569 ( .A1(G543), .A2(n526), .ZN(n521) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n521), .Z(n649) );
  NAND2_X1 U571 ( .A1(n649), .A2(G63), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U573 ( .A(KEYINPUT6), .B(n524), .ZN(n532) );
  NOR2_X1 U574 ( .A1(G651), .A2(G543), .ZN(n634) );
  NAND2_X1 U575 ( .A1(n634), .A2(G89), .ZN(n525) );
  XNOR2_X1 U576 ( .A(n525), .B(KEYINPUT4), .ZN(n528) );
  NOR2_X2 U577 ( .A1(n645), .A2(n526), .ZN(n637) );
  NAND2_X1 U578 ( .A1(G76), .A2(n637), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U580 ( .A(KEYINPUT76), .B(n529), .Z(n530) );
  XNOR2_X1 U581 ( .A(KEYINPUT5), .B(n530), .ZN(n531) );
  NOR2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U583 ( .A(KEYINPUT7), .B(n533), .Z(G168) );
  XOR2_X1 U584 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U585 ( .A(KEYINPUT64), .B(KEYINPUT23), .Z(n535) );
  INV_X1 U586 ( .A(G2105), .ZN(n540) );
  AND2_X1 U587 ( .A1(n540), .A2(G2104), .ZN(n877) );
  NAND2_X1 U588 ( .A1(G101), .A2(n877), .ZN(n534) );
  XNOR2_X1 U589 ( .A(n535), .B(n534), .ZN(n539) );
  XNOR2_X1 U590 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n537) );
  NOR2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  XNOR2_X2 U592 ( .A(n537), .B(n536), .ZN(n878) );
  NAND2_X1 U593 ( .A1(n878), .A2(G137), .ZN(n538) );
  AND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n683) );
  NAND2_X1 U595 ( .A1(G125), .A2(n881), .ZN(n542) );
  AND2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n882) );
  NAND2_X1 U597 ( .A1(G113), .A2(n882), .ZN(n541) );
  AND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n681) );
  AND2_X1 U599 ( .A1(n683), .A2(n681), .ZN(G160) );
  NAND2_X1 U600 ( .A1(G138), .A2(n878), .ZN(n548) );
  AND2_X1 U601 ( .A1(G102), .A2(n877), .ZN(n546) );
  NAND2_X1 U602 ( .A1(G126), .A2(n881), .ZN(n544) );
  NAND2_X1 U603 ( .A1(G114), .A2(n882), .ZN(n543) );
  NAND2_X1 U604 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U605 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(G164) );
  INV_X1 U607 ( .A(G132), .ZN(G219) );
  INV_X1 U608 ( .A(G82), .ZN(G220) );
  NAND2_X1 U609 ( .A1(n644), .A2(G52), .ZN(n549) );
  XNOR2_X1 U610 ( .A(KEYINPUT67), .B(n549), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G77), .A2(n637), .ZN(n551) );
  NAND2_X1 U612 ( .A1(G90), .A2(n634), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U614 ( .A(n552), .B(KEYINPUT9), .ZN(n553) );
  XNOR2_X1 U615 ( .A(n553), .B(KEYINPUT68), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n649), .A2(G64), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U618 ( .A1(n557), .A2(n556), .ZN(G171) );
  NAND2_X1 U619 ( .A1(G94), .A2(G452), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n558), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U623 ( .A(G223), .ZN(n829) );
  NAND2_X1 U624 ( .A1(n829), .A2(G567), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  XOR2_X1 U626 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n562) );
  NAND2_X1 U627 ( .A1(G56), .A2(n649), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n634), .A2(G81), .ZN(n563) );
  XNOR2_X1 U630 ( .A(KEYINPUT12), .B(n563), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n637), .A2(G68), .ZN(n564) );
  XOR2_X1 U632 ( .A(KEYINPUT73), .B(n564), .Z(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT13), .ZN(n569) );
  NAND2_X1 U635 ( .A1(G43), .A2(n644), .ZN(n568) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U637 ( .A1(G860), .A2(n924), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT74), .ZN(G153) );
  INV_X1 U639 ( .A(G171), .ZN(G301) );
  NAND2_X1 U640 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U641 ( .A1(n644), .A2(G54), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G79), .A2(n637), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G66), .A2(n649), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U645 ( .A1(G92), .A2(n634), .ZN(n575) );
  XNOR2_X1 U646 ( .A(KEYINPUT75), .B(n575), .ZN(n576) );
  NOR2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U649 ( .A(KEYINPUT15), .B(n580), .Z(n919) );
  INV_X1 U650 ( .A(G868), .ZN(n664) );
  NAND2_X1 U651 ( .A1(n919), .A2(n664), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U653 ( .A1(G78), .A2(n637), .ZN(n584) );
  NAND2_X1 U654 ( .A1(G91), .A2(n634), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U656 ( .A(KEYINPUT70), .B(n585), .Z(n589) );
  NAND2_X1 U657 ( .A1(G65), .A2(n649), .ZN(n587) );
  NAND2_X1 U658 ( .A1(G53), .A2(n644), .ZN(n586) );
  AND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(G299) );
  NOR2_X1 U661 ( .A1(G286), .A2(n664), .ZN(n591) );
  NOR2_X1 U662 ( .A1(G868), .A2(G299), .ZN(n590) );
  NOR2_X1 U663 ( .A1(n591), .A2(n590), .ZN(G297) );
  INV_X1 U664 ( .A(G860), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n592), .A2(G559), .ZN(n593) );
  INV_X1 U666 ( .A(n919), .ZN(n616) );
  NAND2_X1 U667 ( .A1(n593), .A2(n616), .ZN(n594) );
  XNOR2_X1 U668 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U669 ( .A1(G559), .A2(n664), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n616), .A2(n595), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n924), .A2(n664), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U673 ( .A(KEYINPUT78), .B(n598), .Z(G282) );
  XNOR2_X1 U674 ( .A(G2100), .B(KEYINPUT81), .ZN(n609) );
  NAND2_X1 U675 ( .A1(n881), .A2(G123), .ZN(n599) );
  XNOR2_X1 U676 ( .A(n599), .B(KEYINPUT18), .ZN(n601) );
  NAND2_X1 U677 ( .A1(G135), .A2(n878), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U679 ( .A(n602), .B(KEYINPUT79), .ZN(n604) );
  NAND2_X1 U680 ( .A1(G99), .A2(n877), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n882), .A2(G111), .ZN(n605) );
  XOR2_X1 U683 ( .A(KEYINPUT80), .B(n605), .Z(n606) );
  NOR2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n973) );
  XNOR2_X1 U685 ( .A(n973), .B(G2096), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(G156) );
  NAND2_X1 U687 ( .A1(G80), .A2(n637), .ZN(n611) );
  NAND2_X1 U688 ( .A1(G67), .A2(n649), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U690 ( .A1(G93), .A2(n634), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G55), .A2(n644), .ZN(n612) );
  NAND2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n614) );
  OR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n663) );
  NAND2_X1 U694 ( .A1(n616), .A2(G559), .ZN(n661) );
  XOR2_X1 U695 ( .A(n924), .B(n661), .Z(n617) );
  NOR2_X1 U696 ( .A1(G860), .A2(n617), .ZN(n618) );
  XOR2_X1 U697 ( .A(n663), .B(n618), .Z(G145) );
  NAND2_X1 U698 ( .A1(G72), .A2(n637), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G85), .A2(n634), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U701 ( .A(KEYINPUT66), .B(n621), .Z(n625) );
  NAND2_X1 U702 ( .A1(G60), .A2(n649), .ZN(n623) );
  NAND2_X1 U703 ( .A1(G47), .A2(n644), .ZN(n622) );
  AND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(G290) );
  NAND2_X1 U706 ( .A1(G75), .A2(n637), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G88), .A2(n634), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U709 ( .A(KEYINPUT85), .B(n628), .ZN(n632) );
  NAND2_X1 U710 ( .A1(G62), .A2(n649), .ZN(n630) );
  NAND2_X1 U711 ( .A1(G50), .A2(n644), .ZN(n629) );
  AND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(G303) );
  INV_X1 U714 ( .A(G303), .ZN(G166) );
  NAND2_X1 U715 ( .A1(G61), .A2(n649), .ZN(n633) );
  XNOR2_X1 U716 ( .A(n633), .B(KEYINPUT84), .ZN(n642) );
  NAND2_X1 U717 ( .A1(G86), .A2(n634), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G48), .A2(n644), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n637), .A2(G73), .ZN(n638) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(n638), .Z(n639) );
  NOR2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(G305) );
  NAND2_X1 U724 ( .A1(G74), .A2(G651), .ZN(n643) );
  XNOR2_X1 U725 ( .A(n643), .B(KEYINPUT82), .ZN(n651) );
  NAND2_X1 U726 ( .A1(G49), .A2(n644), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G87), .A2(n645), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U731 ( .A(KEYINPUT83), .B(n652), .Z(G288) );
  INV_X1 U732 ( .A(G299), .ZN(n915) );
  XNOR2_X1 U733 ( .A(n915), .B(G290), .ZN(n658) );
  XOR2_X1 U734 ( .A(KEYINPUT19), .B(KEYINPUT87), .Z(n654) );
  XNOR2_X1 U735 ( .A(G166), .B(KEYINPUT86), .ZN(n653) );
  XNOR2_X1 U736 ( .A(n654), .B(n653), .ZN(n656) );
  XNOR2_X1 U737 ( .A(n924), .B(n663), .ZN(n655) );
  XNOR2_X1 U738 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U739 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n659), .B(G305), .ZN(n660) );
  XNOR2_X1 U741 ( .A(n660), .B(G288), .ZN(n856) );
  XNOR2_X1 U742 ( .A(n661), .B(n856), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n662), .A2(G868), .ZN(n666) );
  NAND2_X1 U744 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U745 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U753 ( .A1(G108), .A2(G120), .ZN(n671) );
  NOR2_X1 U754 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U755 ( .A1(G69), .A2(n672), .ZN(n833) );
  NAND2_X1 U756 ( .A1(n833), .A2(G567), .ZN(n677) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U759 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U760 ( .A1(G96), .A2(n675), .ZN(n834) );
  NAND2_X1 U761 ( .A1(n834), .A2(G2106), .ZN(n676) );
  NAND2_X1 U762 ( .A1(n677), .A2(n676), .ZN(n860) );
  NAND2_X1 U763 ( .A1(G661), .A2(G483), .ZN(n678) );
  XNOR2_X1 U764 ( .A(KEYINPUT88), .B(n678), .ZN(n679) );
  NOR2_X1 U765 ( .A1(n860), .A2(n679), .ZN(n832) );
  NAND2_X1 U766 ( .A1(n832), .A2(G36), .ZN(G176) );
  NOR2_X2 U767 ( .A1(G164), .A2(G1384), .ZN(n771) );
  AND2_X1 U768 ( .A1(n681), .A2(G40), .ZN(n682) );
  AND2_X1 U769 ( .A1(n683), .A2(n682), .ZN(n769) );
  NAND2_X1 U770 ( .A1(G8), .A2(n718), .ZN(n764) );
  NOR2_X1 U771 ( .A1(G1971), .A2(n764), .ZN(n685) );
  NOR2_X1 U772 ( .A1(G2090), .A2(n718), .ZN(n684) );
  NOR2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U774 ( .A1(n686), .A2(G303), .ZN(n687) );
  XNOR2_X1 U775 ( .A(KEYINPUT102), .B(n687), .ZN(n737) );
  XNOR2_X1 U776 ( .A(G1996), .B(KEYINPUT95), .ZN(n1002) );
  NOR2_X1 U777 ( .A1(n718), .A2(n1002), .ZN(n689) );
  XOR2_X1 U778 ( .A(KEYINPUT26), .B(KEYINPUT96), .Z(n688) );
  XNOR2_X1 U779 ( .A(n689), .B(n688), .ZN(n691) );
  NAND2_X1 U780 ( .A1(n718), .A2(G1341), .ZN(n690) );
  NAND2_X1 U781 ( .A1(n691), .A2(n690), .ZN(n696) );
  NAND2_X1 U782 ( .A1(G1348), .A2(n718), .ZN(n693) );
  INV_X1 U783 ( .A(n718), .ZN(n712) );
  NAND2_X1 U784 ( .A1(n712), .A2(G2067), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U786 ( .A1(n919), .A2(n697), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n924), .A2(n694), .ZN(n695) );
  NOR2_X1 U788 ( .A1(n696), .A2(n695), .ZN(n699) );
  NOR2_X1 U789 ( .A1(n697), .A2(n919), .ZN(n698) );
  NOR2_X1 U790 ( .A1(n699), .A2(n698), .ZN(n704) );
  NAND2_X1 U791 ( .A1(n712), .A2(G2072), .ZN(n700) );
  XNOR2_X1 U792 ( .A(n700), .B(KEYINPUT27), .ZN(n702) );
  INV_X1 U793 ( .A(G1956), .ZN(n942) );
  NOR2_X1 U794 ( .A1(n942), .A2(n712), .ZN(n701) );
  NOR2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U796 ( .A1(n915), .A2(n705), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n709) );
  NOR2_X1 U798 ( .A1(n915), .A2(n705), .ZN(n707) );
  XOR2_X1 U799 ( .A(KEYINPUT28), .B(KEYINPUT94), .Z(n706) );
  XNOR2_X1 U800 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n711) );
  XOR2_X1 U802 ( .A(KEYINPUT29), .B(KEYINPUT97), .Z(n710) );
  XNOR2_X1 U803 ( .A(n711), .B(n710), .ZN(n716) );
  NAND2_X1 U804 ( .A1(G1961), .A2(n718), .ZN(n714) );
  XOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .Z(n1003) );
  NAND2_X1 U806 ( .A1(n712), .A2(n1003), .ZN(n713) );
  NAND2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n717) );
  NOR2_X1 U808 ( .A1(G301), .A2(n717), .ZN(n715) );
  NOR2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n731) );
  AND2_X1 U810 ( .A1(G301), .A2(n717), .ZN(n726) );
  INV_X1 U811 ( .A(KEYINPUT93), .ZN(n720) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n718), .ZN(n719) );
  XNOR2_X1 U813 ( .A(n720), .B(n719), .ZN(n740) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n764), .ZN(n743) );
  NOR2_X1 U815 ( .A1(n740), .A2(n743), .ZN(n721) );
  XNOR2_X1 U816 ( .A(n721), .B(KEYINPUT98), .ZN(n722) );
  NAND2_X1 U817 ( .A1(n722), .A2(G8), .ZN(n723) );
  XNOR2_X1 U818 ( .A(n723), .B(KEYINPUT30), .ZN(n724) );
  NOR2_X1 U819 ( .A1(G168), .A2(n724), .ZN(n725) );
  NOR2_X1 U820 ( .A1(n726), .A2(n725), .ZN(n729) );
  INV_X1 U821 ( .A(KEYINPUT31), .ZN(n727) );
  NOR2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n733) );
  INV_X1 U823 ( .A(KEYINPUT100), .ZN(n732) );
  XNOR2_X1 U824 ( .A(n733), .B(n732), .ZN(n741) );
  NAND2_X1 U825 ( .A1(n741), .A2(G286), .ZN(n735) );
  NAND2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U827 ( .A1(n738), .A2(G8), .ZN(n739) );
  NAND2_X1 U828 ( .A1(G8), .A2(n740), .ZN(n745) );
  INV_X1 U829 ( .A(n741), .ZN(n742) );
  NOR2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U832 ( .A1(n747), .A2(n746), .ZN(n759) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n752) );
  NOR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U835 ( .A1(n752), .A2(n748), .ZN(n917) );
  NAND2_X1 U836 ( .A1(n759), .A2(n917), .ZN(n749) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n926) );
  NAND2_X1 U838 ( .A1(n749), .A2(n926), .ZN(n750) );
  NOR2_X1 U839 ( .A1(n750), .A2(n764), .ZN(n751) );
  NOR2_X1 U840 ( .A1(KEYINPUT33), .A2(n751), .ZN(n756) );
  NAND2_X1 U841 ( .A1(n752), .A2(KEYINPUT33), .ZN(n753) );
  XNOR2_X1 U842 ( .A(G1981), .B(KEYINPUT103), .ZN(n754) );
  XNOR2_X1 U843 ( .A(n754), .B(G305), .ZN(n912) );
  NOR2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n768) );
  NOR2_X1 U845 ( .A1(G2090), .A2(G303), .ZN(n757) );
  NAND2_X1 U846 ( .A1(G8), .A2(n757), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n760), .A2(n764), .ZN(n766) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n761) );
  XOR2_X1 U850 ( .A(n761), .B(KEYINPUT92), .Z(n762) );
  XNOR2_X1 U851 ( .A(KEYINPUT24), .B(n762), .ZN(n763) );
  OR2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n793) );
  INV_X1 U855 ( .A(n769), .ZN(n770) );
  NOR2_X1 U856 ( .A1(n771), .A2(n770), .ZN(n813) );
  INV_X1 U857 ( .A(n813), .ZN(n791) );
  XNOR2_X1 U858 ( .A(G1986), .B(G290), .ZN(n928) );
  XOR2_X1 U859 ( .A(KEYINPUT90), .B(KEYINPUT38), .Z(n773) );
  NAND2_X1 U860 ( .A1(G105), .A2(n877), .ZN(n772) );
  XNOR2_X1 U861 ( .A(n773), .B(n772), .ZN(n777) );
  NAND2_X1 U862 ( .A1(G129), .A2(n881), .ZN(n775) );
  NAND2_X1 U863 ( .A1(G117), .A2(n882), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U866 ( .A(KEYINPUT91), .B(n778), .Z(n780) );
  NAND2_X1 U867 ( .A1(n878), .A2(G141), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n890) );
  NAND2_X1 U869 ( .A1(G1996), .A2(n890), .ZN(n789) );
  NAND2_X1 U870 ( .A1(G119), .A2(n881), .ZN(n782) );
  NAND2_X1 U871 ( .A1(G131), .A2(n878), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G107), .A2(n882), .ZN(n783) );
  XNOR2_X1 U874 ( .A(KEYINPUT89), .B(n783), .ZN(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n877), .A2(G95), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n889) );
  NAND2_X1 U878 ( .A1(G1991), .A2(n889), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n972) );
  NOR2_X1 U880 ( .A1(n928), .A2(n972), .ZN(n790) );
  NOR2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n803) );
  XNOR2_X1 U883 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NAND2_X1 U884 ( .A1(G104), .A2(n877), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G140), .A2(n878), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U887 ( .A(KEYINPUT34), .B(n796), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G128), .A2(n881), .ZN(n798) );
  NAND2_X1 U889 ( .A1(G116), .A2(n882), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U891 ( .A(KEYINPUT35), .B(n799), .Z(n800) );
  NOR2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n802), .ZN(n901) );
  NOR2_X1 U894 ( .A1(n810), .A2(n901), .ZN(n977) );
  NAND2_X1 U895 ( .A1(n977), .A2(n813), .ZN(n808) );
  NAND2_X1 U896 ( .A1(n803), .A2(n808), .ZN(n816) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n890), .ZN(n967) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U899 ( .A1(G1991), .A2(n889), .ZN(n971) );
  NOR2_X1 U900 ( .A1(n804), .A2(n971), .ZN(n805) );
  NOR2_X1 U901 ( .A1(n972), .A2(n805), .ZN(n806) );
  NOR2_X1 U902 ( .A1(n967), .A2(n806), .ZN(n807) );
  XNOR2_X1 U903 ( .A(n807), .B(KEYINPUT39), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n810), .A2(n901), .ZN(n985) );
  NAND2_X1 U906 ( .A1(n811), .A2(n985), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U908 ( .A(n814), .B(KEYINPUT104), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U910 ( .A(n817), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U911 ( .A(G2446), .B(G2451), .ZN(n827) );
  XOR2_X1 U912 ( .A(G2430), .B(KEYINPUT106), .Z(n819) );
  XNOR2_X1 U913 ( .A(G2454), .B(G2435), .ZN(n818) );
  XNOR2_X1 U914 ( .A(n819), .B(n818), .ZN(n823) );
  XOR2_X1 U915 ( .A(G2438), .B(KEYINPUT105), .Z(n821) );
  XNOR2_X1 U916 ( .A(G1348), .B(G1341), .ZN(n820) );
  XNOR2_X1 U917 ( .A(n821), .B(n820), .ZN(n822) );
  XOR2_X1 U918 ( .A(n823), .B(n822), .Z(n825) );
  XNOR2_X1 U919 ( .A(G2427), .B(G2443), .ZN(n824) );
  XNOR2_X1 U920 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U921 ( .A(n827), .B(n826), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n828), .A2(G14), .ZN(n906) );
  XNOR2_X1 U923 ( .A(KEYINPUT107), .B(n906), .ZN(G401) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U926 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(KEYINPUT41), .B(G1991), .Z(n836) );
  XNOR2_X1 U937 ( .A(G1996), .B(G1961), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U939 ( .A(n837), .B(G2474), .Z(n839) );
  XNOR2_X1 U940 ( .A(G1966), .B(G1981), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U942 ( .A(G1986), .B(G1976), .Z(n841) );
  XNOR2_X1 U943 ( .A(G1956), .B(G1971), .ZN(n840) );
  XNOR2_X1 U944 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U945 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U946 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(G229) );
  XOR2_X1 U948 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n847) );
  XNOR2_X1 U949 ( .A(KEYINPUT108), .B(G2678), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U951 ( .A(KEYINPUT42), .B(G2090), .Z(n849) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U953 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U954 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U955 ( .A(G2096), .B(G2100), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n853), .B(n852), .ZN(n855) );
  XOR2_X1 U957 ( .A(G2078), .B(G2084), .Z(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(G227) );
  XNOR2_X1 U959 ( .A(G286), .B(n856), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n919), .B(G171), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n859) );
  NOR2_X1 U962 ( .A1(G37), .A2(n859), .ZN(G397) );
  INV_X1 U963 ( .A(n860), .ZN(G319) );
  NAND2_X1 U964 ( .A1(n881), .A2(G124), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U966 ( .A1(G112), .A2(n882), .ZN(n862) );
  NAND2_X1 U967 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G100), .A2(n877), .ZN(n865) );
  NAND2_X1 U969 ( .A1(G136), .A2(n878), .ZN(n864) );
  NAND2_X1 U970 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U971 ( .A1(n867), .A2(n866), .ZN(G162) );
  XNOR2_X1 U972 ( .A(KEYINPUT113), .B(KEYINPUT45), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G106), .A2(n877), .ZN(n869) );
  NAND2_X1 U974 ( .A1(G142), .A2(n878), .ZN(n868) );
  NAND2_X1 U975 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U976 ( .A(n871), .B(n870), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n882), .A2(G118), .ZN(n872) );
  XNOR2_X1 U978 ( .A(n872), .B(KEYINPUT112), .ZN(n874) );
  NAND2_X1 U979 ( .A1(G130), .A2(n881), .ZN(n873) );
  NAND2_X1 U980 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U981 ( .A1(n876), .A2(n875), .ZN(n894) );
  NAND2_X1 U982 ( .A1(G103), .A2(n877), .ZN(n880) );
  NAND2_X1 U983 ( .A1(G139), .A2(n878), .ZN(n879) );
  NAND2_X1 U984 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G127), .A2(n881), .ZN(n884) );
  NAND2_X1 U986 ( .A1(G115), .A2(n882), .ZN(n883) );
  NAND2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U990 ( .A(KEYINPUT114), .B(n888), .Z(n981) );
  XNOR2_X1 U991 ( .A(G162), .B(n889), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n981), .B(n892), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n898) );
  XOR2_X1 U995 ( .A(KEYINPUT115), .B(KEYINPUT48), .Z(n896) );
  XNOR2_X1 U996 ( .A(n973), .B(KEYINPUT46), .ZN(n895) );
  XNOR2_X1 U997 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U998 ( .A(n898), .B(n897), .Z(n900) );
  XNOR2_X1 U999 ( .A(G160), .B(G164), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n903), .ZN(G395) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n904) );
  XOR2_X1 U1004 ( .A(KEYINPUT116), .B(n904), .Z(n905) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n905), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n906), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(G397), .A2(n907), .ZN(n908) );
  NAND2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n910) );
  NOR2_X1 U1009 ( .A1(n910), .A2(G395), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n911), .B(KEYINPUT117), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1012 ( .A(G16), .B(KEYINPUT56), .ZN(n936) );
  XNOR2_X1 U1013 ( .A(G1966), .B(G168), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(n914), .B(KEYINPUT57), .ZN(n934) );
  XNOR2_X1 U1016 ( .A(n942), .B(n915), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(KEYINPUT123), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(G171), .B(G1961), .ZN(n918) );
  NAND2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(G1348), .B(n919), .ZN(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n932) );
  XNOR2_X1 U1023 ( .A(n924), .B(G1341), .ZN(n930) );
  NAND2_X1 U1024 ( .A1(G1971), .A2(G303), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(n964) );
  INV_X1 U1031 ( .A(G16), .ZN(n962) );
  XOR2_X1 U1032 ( .A(G1976), .B(G23), .Z(n938) );
  XOR2_X1 U1033 ( .A(G1971), .B(G22), .Z(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G24), .B(G1986), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1037 ( .A(KEYINPUT58), .B(n941), .Z(n958) );
  XOR2_X1 U1038 ( .A(G1961), .B(G5), .Z(n952) );
  XNOR2_X1 U1039 ( .A(G20), .B(n942), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G1341), .B(G19), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(G6), .B(G1981), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n949) );
  XOR2_X1 U1044 ( .A(KEYINPUT59), .B(G1348), .Z(n947) );
  XNOR2_X1 U1045 ( .A(G4), .B(n947), .ZN(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(KEYINPUT60), .B(n950), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(KEYINPUT124), .B(G1966), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(G21), .B(n953), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT125), .B(n956), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(n959), .B(KEYINPUT61), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n960), .B(KEYINPUT126), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(n965), .B(KEYINPUT127), .ZN(n994) );
  XOR2_X1 U1059 ( .A(G2090), .B(G162), .Z(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1061 ( .A(KEYINPUT51), .B(n968), .Z(n969) );
  XNOR2_X1 U1062 ( .A(KEYINPUT118), .B(n969), .ZN(n979) );
  XOR2_X1 U1063 ( .A(G2084), .B(G160), .Z(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n975) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n988) );
  XNOR2_X1 U1069 ( .A(G164), .B(G2078), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n980), .B(KEYINPUT119), .ZN(n983) );
  XNOR2_X1 U1071 ( .A(n981), .B(G2072), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(n984), .B(KEYINPUT50), .ZN(n986) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(KEYINPUT52), .B(n989), .ZN(n991) );
  INV_X1 U1077 ( .A(KEYINPUT55), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n992), .A2(G29), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n1020) );
  XOR2_X1 U1081 ( .A(G1991), .B(G25), .Z(n995) );
  NAND2_X1 U1082 ( .A1(n995), .A2(G28), .ZN(n1001) );
  XNOR2_X1 U1083 ( .A(G2072), .B(G33), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(n996), .B(KEYINPUT120), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(G26), .B(G2067), .ZN(n997) );
  NOR2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(n999), .B(KEYINPUT121), .ZN(n1000) );
  NOR2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1007) );
  XOR2_X1 U1089 ( .A(n1002), .B(G32), .Z(n1005) );
  XNOR2_X1 U1090 ( .A(n1003), .B(G27), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(n1008), .B(KEYINPUT53), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(G2084), .B(G34), .Z(n1009) );
  XNOR2_X1 U1095 ( .A(KEYINPUT54), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G35), .B(G2090), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(n1014), .B(KEYINPUT55), .ZN(n1016) );
  INV_X1 U1100 ( .A(G29), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(G11), .A2(n1017), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(KEYINPUT122), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1021), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

