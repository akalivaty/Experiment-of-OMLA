//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(G122), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G122), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n188), .A2(new_n190), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G128), .B(G143), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G128), .ZN(new_n201));
  OAI21_X1  g015(.A(G134), .B1(new_n201), .B2(KEYINPUT13), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n202), .B1(KEYINPUT13), .B2(new_n196), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT92), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n196), .A2(KEYINPUT13), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT92), .B1(new_n206), .B2(new_n202), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n199), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n201), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G134), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT93), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n213), .A2(new_n198), .B1(new_n214), .B2(new_n194), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n188), .B1(new_n190), .B2(KEYINPUT14), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n190), .A2(KEYINPUT14), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n217), .A2(KEYINPUT94), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(KEYINPUT94), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OAI221_X1 g034(.A(new_n215), .B1(new_n214), .B2(new_n194), .C1(new_n220), .C2(new_n193), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n209), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(KEYINPUT9), .B(G234), .Z(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(KEYINPUT78), .ZN(new_n224));
  INV_X1    g038(.A(G217), .ZN(new_n225));
  OR3_X1    g039(.A1(new_n224), .A2(new_n225), .A3(G953), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n224), .A2(new_n225), .A3(G953), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n209), .A2(new_n221), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT72), .B(G902), .Z(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G478), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(KEYINPUT15), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n234), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n230), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(KEYINPUT95), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT95), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n236), .B1(new_n230), .B2(new_n231), .ZN(new_n240));
  INV_X1    g054(.A(new_n231), .ZN(new_n241));
  AOI211_X1 g055(.A(new_n241), .B(new_n234), .C1(new_n227), .C2(new_n229), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G953), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n245), .A2(G952), .ZN(new_n246));
  INV_X1    g060(.A(G234), .ZN(new_n247));
  INV_X1    g061(.A(G237), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AOI211_X1 g064(.A(new_n245), .B(new_n231), .C1(G234), .C2(G237), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT21), .B(G898), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G902), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n248), .A2(new_n245), .A3(G214), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n255), .B(G143), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT18), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n255), .B(new_n200), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT18), .A3(G131), .ZN(new_n261));
  XNOR2_X1  g075(.A(G125), .B(G140), .ZN(new_n262));
  INV_X1    g076(.A(G146), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n259), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n260), .A2(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n256), .A2(new_n258), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT17), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n262), .A2(KEYINPUT16), .ZN(new_n270));
  INV_X1    g084(.A(G125), .ZN(new_n271));
  OR3_X1    g085(.A1(new_n271), .A2(KEYINPUT16), .A3(G140), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n263), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n270), .A2(G146), .A3(new_n272), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n274), .B(new_n275), .C1(new_n266), .C2(new_n268), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n265), .B1(new_n269), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(G113), .B(G122), .ZN(new_n278));
  INV_X1    g092(.A(G104), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n280), .B(new_n265), .C1(new_n269), .C2(new_n276), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n254), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G475), .ZN(new_n286));
  NOR2_X1   g100(.A1(G475), .A2(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n266), .A2(new_n267), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n262), .B(KEYINPUT19), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n263), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n275), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n265), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n281), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n288), .B1(new_n294), .B2(new_n283), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT20), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n295), .A2(new_n296), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n286), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n244), .A2(new_n253), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G214), .B1(G237), .B2(G902), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G210), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT68), .B1(new_n189), .B2(G119), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n308));
  INV_X1    g122(.A(G119), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(G116), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n307), .A2(new_n310), .B1(new_n189), .B2(G119), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT5), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(G116), .ZN(new_n313));
  OAI21_X1  g127(.A(G113), .B1(new_n313), .B2(KEYINPUT5), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT2), .B(G113), .Z(new_n317));
  NAND2_X1  g131(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n193), .A2(G104), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n279), .A2(G107), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G101), .ZN(new_n324));
  INV_X1    g138(.A(new_n322), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n321), .A2(G101), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n316), .A2(new_n318), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n326), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n331), .A2(new_n322), .B1(G104), .B2(new_n193), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n325), .B1(new_n319), .B2(new_n320), .ZN(new_n333));
  OAI21_X1  g147(.A(G101), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n334), .A2(new_n328), .A3(KEYINPUT4), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n336), .B(G101), .C1(new_n332), .C2(new_n333), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n311), .A2(new_n317), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n311), .A2(new_n317), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n330), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G122), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT87), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n330), .B(new_n346), .C1(new_n335), .C2(new_n340), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(KEYINPUT6), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n263), .A2(G143), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n200), .A2(G146), .ZN(new_n352));
  NAND2_X1  g166(.A1(KEYINPUT0), .A2(G128), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(KEYINPUT0), .B(G128), .Z(new_n355));
  XNOR2_X1  g169(.A(G143), .B(G146), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT88), .B1(new_n357), .B2(new_n271), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n351), .A2(new_n352), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT0), .B(G128), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT88), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n361), .A2(new_n362), .A3(G125), .A4(new_n354), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n200), .B(G146), .C1(new_n210), .C2(KEYINPUT1), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n210), .A2(new_n263), .A3(G143), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n351), .A3(new_n352), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n271), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n363), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G224), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(G953), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n371), .B(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n341), .A2(new_n375), .A3(new_n347), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n350), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT89), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n350), .A2(KEYINPUT89), .A3(new_n374), .A4(new_n376), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT7), .B1(new_n372), .B2(G953), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n371), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n382), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n358), .A2(new_n363), .A3(new_n370), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT8), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n344), .A2(new_n387), .A3(new_n345), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n387), .B1(new_n344), .B2(new_n345), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n328), .A2(new_n329), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n314), .B1(new_n311), .B2(KEYINPUT5), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n391), .B1(new_n338), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n390), .B1(new_n393), .B2(new_n330), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT90), .B1(new_n386), .B2(new_n394), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n391), .A2(new_n338), .A3(new_n392), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n316), .A2(new_n318), .B1(new_n328), .B2(new_n329), .ZN(new_n397));
  OAI22_X1  g211(.A1(new_n396), .A2(new_n397), .B1(new_n389), .B2(new_n388), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n398), .A2(new_n399), .A3(new_n383), .A4(new_n385), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n395), .A2(new_n400), .A3(new_n349), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n381), .A2(new_n401), .A3(new_n254), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n306), .B1(new_n380), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n349), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n383), .A3(new_n385), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(KEYINPUT90), .ZN(new_n406));
  AOI21_X1  g220(.A(G902), .B1(new_n406), .B2(new_n400), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n407), .A2(new_n379), .A3(new_n305), .A4(new_n381), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n403), .A2(KEYINPUT91), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT91), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n410), .B(new_n306), .C1(new_n380), .C2(new_n402), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n302), .A2(new_n304), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT23), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n309), .B2(G128), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n309), .A2(G128), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n418), .A2(KEYINPUT75), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(KEYINPUT75), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(G110), .A3(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(KEYINPUT24), .B(G110), .Z(new_n422));
  XNOR2_X1  g236(.A(G119), .B(G128), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT74), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n274), .A2(new_n275), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n262), .A2(new_n263), .ZN(new_n428));
  INV_X1    g242(.A(G110), .ZN(new_n429));
  AND4_X1   g243(.A1(new_n429), .A2(new_n415), .A3(new_n416), .A4(new_n417), .ZN(new_n430));
  OAI22_X1  g244(.A1(new_n430), .A2(KEYINPUT76), .B1(new_n423), .B2(new_n422), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n430), .A2(KEYINPUT76), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n275), .B(new_n428), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT22), .B(G137), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT77), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n245), .A2(G221), .A3(G234), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n434), .B(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT25), .B1(new_n439), .B2(new_n241), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n225), .B1(new_n231), .B2(G234), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n439), .A2(KEYINPUT25), .A3(new_n241), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n441), .A2(G902), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n450));
  INV_X1    g264(.A(G137), .ZN(new_n451));
  AND2_X1   g265(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n452));
  NOR2_X1   g266(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n453));
  OAI211_X1 g267(.A(G134), .B(new_n451), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT65), .B1(new_n451), .B2(G134), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT65), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n197), .A3(G137), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n197), .B2(G137), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n454), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G131), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n454), .A2(new_n458), .A3(new_n258), .A4(new_n460), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n462), .A2(new_n463), .B1(new_n361), .B2(new_n354), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n367), .A2(new_n369), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT66), .B1(new_n197), .B2(G137), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(G134), .B2(new_n451), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n197), .A2(KEYINPUT66), .A3(G137), .ZN(new_n468));
  OAI21_X1  g282(.A(G131), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n465), .A2(new_n469), .A3(new_n463), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n450), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT67), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n338), .A2(new_n339), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT67), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n475), .B(new_n450), .C1(new_n464), .C2(new_n470), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n465), .A2(new_n469), .A3(new_n463), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n357), .A2(KEYINPUT69), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT69), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n361), .A2(new_n479), .A3(new_n354), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n462), .A2(new_n463), .ZN(new_n482));
  OAI211_X1 g296(.A(KEYINPUT30), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n472), .A2(new_n474), .A3(new_n476), .A4(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n473), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n248), .A2(new_n245), .A3(G210), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT26), .B(G101), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n484), .A2(new_n485), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT31), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT28), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n485), .A2(new_n494), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n464), .A2(new_n470), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n474), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n462), .A2(new_n463), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n478), .A2(new_n480), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n470), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT28), .A3(new_n473), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n490), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT31), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n484), .A2(new_n504), .A3(new_n485), .A4(new_n491), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n493), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(G472), .A2(G902), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT71), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT32), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(KEYINPUT71), .A3(new_n507), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n477), .B1(new_n481), .B2(new_n482), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n474), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT29), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n490), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n495), .A2(new_n501), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n231), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT73), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n521), .A3(new_n231), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n516), .B1(new_n502), .B2(new_n490), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n491), .B1(new_n484), .B2(new_n485), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(G472), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n506), .A2(KEYINPUT32), .A3(new_n507), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n449), .B1(new_n513), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(G110), .B(G140), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n245), .A2(G227), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT10), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT80), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n356), .A2(new_n535), .A3(new_n368), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n366), .A2(KEYINPUT81), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT81), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n364), .A2(new_n538), .A3(new_n365), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n369), .A2(KEYINPUT80), .ZN(new_n540));
  AND4_X1   g354(.A1(new_n536), .A2(new_n537), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n534), .B1(new_n541), .B2(new_n391), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n334), .A2(new_n328), .A3(KEYINPUT4), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n499), .A2(new_n543), .A3(new_n337), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n328), .A2(new_n329), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n366), .B1(new_n356), .B2(new_n368), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(new_n534), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n542), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT82), .B1(new_n549), .B2(new_n498), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n537), .A2(new_n540), .A3(new_n536), .A4(new_n539), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n552), .A2(new_n534), .B1(new_n547), .B2(new_n545), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT82), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n553), .A2(new_n554), .A3(new_n482), .A4(new_n544), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n533), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n549), .A2(KEYINPUT83), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT83), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n542), .A2(new_n544), .A3(new_n558), .A4(new_n548), .ZN(new_n559));
  AND4_X1   g373(.A1(KEYINPUT84), .A2(new_n557), .A3(new_n498), .A4(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n482), .B1(new_n549), .B2(KEYINPUT83), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT84), .B1(new_n561), .B2(new_n559), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n556), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n550), .A2(new_n555), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n391), .A2(new_n546), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n482), .B1(new_n552), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT12), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n533), .ZN(new_n569));
  AOI21_X1  g383(.A(G902), .B1(new_n563), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT85), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT85), .ZN(new_n573));
  INV_X1    g387(.A(new_n533), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n564), .B2(new_n567), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n557), .A2(new_n498), .A3(new_n559), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT84), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n561), .A2(KEYINPUT84), .A3(new_n559), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n575), .B1(new_n580), .B2(new_n556), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n573), .B(G469), .C1(new_n581), .C2(G902), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n574), .B1(new_n580), .B2(new_n564), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n564), .A2(new_n567), .A3(new_n574), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n571), .B(new_n231), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n572), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT86), .ZN(new_n587));
  OAI21_X1  g401(.A(G221), .B1(new_n224), .B2(G902), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n413), .B(new_n530), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(G101), .ZN(G3));
  NAND2_X1  g406(.A1(new_n586), .A2(new_n588), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT86), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n304), .B1(new_n403), .B2(new_n408), .ZN(new_n597));
  INV_X1    g411(.A(new_n253), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n300), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n230), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n227), .A2(KEYINPUT33), .A3(new_n229), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n241), .A2(new_n233), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n232), .A2(new_n233), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n599), .A2(new_n600), .A3(new_n608), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n506), .A2(KEYINPUT71), .A3(new_n507), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT71), .B1(new_n506), .B2(new_n507), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n506), .A2(new_n231), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(G472), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n449), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n596), .A2(new_n609), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  NAND3_X1  g433(.A1(new_n295), .A2(KEYINPUT96), .A3(new_n296), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n620), .B1(new_n296), .B2(new_n295), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT96), .B1(new_n295), .B2(new_n296), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n286), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n238), .A2(new_n243), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n599), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n596), .A2(new_n616), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G107), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NOR2_X1   g443(.A1(new_n438), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n434), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n445), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n442), .B2(new_n443), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n612), .A2(new_n614), .A3(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n413), .B(new_n634), .C1(new_n589), .C2(new_n590), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n429), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT97), .B(KEYINPUT37), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G12));
  INV_X1    g452(.A(new_n633), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n513), .B2(new_n529), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n597), .B(new_n640), .C1(new_n589), .C2(new_n590), .ZN(new_n641));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n250), .B1(new_n251), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n625), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n210), .ZN(G30));
  XOR2_X1   g461(.A(new_n643), .B(KEYINPUT39), .Z(new_n648));
  NAND2_X1  g462(.A1(new_n596), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT40), .Z(new_n650));
  NAND2_X1  g464(.A1(new_n484), .A2(new_n485), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n490), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n515), .A2(new_n485), .A3(new_n490), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n254), .ZN(new_n655));
  OAI21_X1  g469(.A(G472), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n513), .A2(new_n528), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n412), .B(KEYINPUT38), .Z(new_n658));
  NOR2_X1   g472(.A1(new_n624), .A2(new_n600), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n660), .A2(new_n304), .A3(new_n633), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n650), .A2(new_n657), .A3(new_n658), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G143), .ZN(G45));
  INV_X1    g477(.A(new_n643), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n300), .A2(new_n607), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n641), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n263), .ZN(G48));
  OAI21_X1  g482(.A(new_n564), .B1(new_n560), .B2(new_n562), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n584), .B1(new_n669), .B2(new_n533), .ZN(new_n670));
  OAI21_X1  g484(.A(G469), .B1(new_n670), .B2(new_n241), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n585), .ZN(new_n672));
  INV_X1    g486(.A(new_n588), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n609), .A2(new_n530), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NAND3_X1  g491(.A1(new_n530), .A2(new_n674), .A3(new_n626), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  AND4_X1   g493(.A1(new_n588), .A2(new_n671), .A3(new_n597), .A4(new_n585), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n640), .A2(new_n680), .A3(new_n301), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G119), .ZN(G21));
  NOR2_X1   g496(.A1(new_n599), .A2(new_n660), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n495), .A2(new_n501), .A3(new_n515), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n493), .B(new_n505), .C1(new_n491), .C2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n507), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n614), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n449), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n674), .A2(new_n683), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G122), .ZN(G24));
  AND4_X1   g504(.A1(new_n614), .A2(new_n665), .A3(new_n633), .A4(new_n686), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n680), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G125), .ZN(G27));
  NOR3_X1   g507(.A1(new_n670), .A2(G469), .A3(new_n241), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n570), .A2(new_n571), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT98), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n666), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT98), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n585), .B(new_n699), .C1(new_n571), .C2(new_n570), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n673), .A2(new_n304), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n409), .B2(new_n411), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n696), .A2(new_n698), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n508), .A2(new_n511), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n449), .B1(new_n529), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n696), .A2(new_n700), .A3(new_n703), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT32), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n527), .A2(new_n528), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n448), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n708), .A2(new_n711), .A3(new_n666), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n707), .B1(new_n712), .B2(KEYINPUT42), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G131), .ZN(G33));
  NOR2_X1   g528(.A1(new_n708), .A2(new_n711), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n644), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT99), .B(G134), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G36));
  NAND2_X1  g532(.A1(new_n581), .A2(KEYINPUT45), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n719), .A2(KEYINPUT100), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(KEYINPUT100), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n581), .A2(KEYINPUT45), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n720), .A2(G469), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(G469), .A2(G902), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n723), .A2(KEYINPUT46), .A3(new_n724), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n585), .A3(new_n728), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n729), .A2(new_n588), .A3(new_n648), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n608), .A2(new_n300), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT43), .B1(new_n608), .B2(new_n300), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n733), .A2(new_n633), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n735), .A2(KEYINPUT44), .A3(new_n615), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT44), .B1(new_n735), .B2(new_n615), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n304), .B1(new_n409), .B2(new_n411), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n730), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G137), .ZN(G39));
  INV_X1    g556(.A(KEYINPUT47), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n729), .A2(new_n743), .A3(new_n588), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n743), .B1(new_n729), .B2(new_n588), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n738), .A2(new_n449), .A3(new_n665), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n709), .A3(new_n710), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G140), .ZN(G42));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n692), .B1(new_n641), .B2(new_n645), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n696), .A2(new_n700), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n659), .A2(new_n597), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n633), .A2(new_n673), .A3(new_n643), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n758), .A3(new_n657), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n641), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(new_n665), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(new_n754), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n759), .B1(new_n641), .B2(new_n666), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n753), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n675), .A2(new_n678), .A3(new_n681), .A4(new_n689), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n755), .A2(new_n530), .A3(new_n665), .A4(new_n703), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n697), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n768), .B1(new_n770), .B2(new_n707), .ZN(new_n771));
  AND4_X1   g585(.A1(new_n691), .A2(new_n696), .A3(new_n700), .A4(new_n703), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n715), .B2(new_n644), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n235), .A2(new_n237), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n623), .A2(new_n774), .A3(new_n643), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n738), .A2(KEYINPUT104), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT104), .B1(new_n738), .B2(new_n775), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n596), .A2(new_n778), .A3(new_n640), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  OAI221_X1 g594(.A(new_n413), .B1(new_n634), .B2(new_n530), .C1(new_n589), .C2(new_n590), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n300), .A2(new_n607), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n774), .B2(new_n600), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n783), .A2(new_n412), .A3(new_n253), .A4(new_n304), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n784), .B(new_n616), .C1(new_n589), .C2(new_n590), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n781), .A2(KEYINPUT103), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT103), .B1(new_n781), .B2(new_n785), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n771), .B(new_n780), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n752), .B1(new_n767), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n754), .A2(new_n762), .A3(KEYINPUT52), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n765), .B1(new_n753), .B2(new_n764), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n675), .A2(new_n678), .A3(new_n681), .A4(new_n689), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n713), .A2(new_n793), .A3(new_n779), .A4(new_n773), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n785), .A2(new_n591), .A3(new_n635), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT103), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n781), .A2(KEYINPUT103), .A3(new_n785), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n792), .A2(new_n799), .A3(KEYINPUT53), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n751), .B1(new_n789), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n801), .A2(KEYINPUT105), .ZN(new_n802));
  INV_X1    g616(.A(new_n800), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT53), .B1(new_n792), .B2(new_n799), .ZN(new_n804));
  OAI211_X1 g618(.A(KEYINPUT105), .B(KEYINPUT54), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT106), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n769), .A2(new_n697), .B1(new_n704), .B2(new_n706), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n806), .B1(new_n807), .B2(new_n768), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n713), .A2(new_n793), .A3(KEYINPUT106), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n773), .A2(new_n779), .A3(KEYINPUT53), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n797), .B2(new_n798), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n810), .B(new_n812), .C1(new_n763), .C2(new_n766), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n788), .B1(new_n791), .B2(new_n790), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n751), .B(new_n813), .C1(new_n814), .C2(KEYINPUT53), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n802), .A2(new_n805), .A3(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n739), .A2(new_n673), .A3(new_n672), .ZN(new_n817));
  INV_X1    g631(.A(new_n657), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n448), .A3(new_n250), .A4(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT112), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(KEYINPUT112), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(new_n782), .ZN(new_n823));
  INV_X1    g637(.A(new_n680), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n733), .A2(new_n250), .A3(new_n734), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n688), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n817), .A2(new_n825), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT110), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n827), .B(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n829), .A2(new_n706), .ZN(new_n830));
  XOR2_X1   g644(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n831));
  OAI221_X1 g645(.A(new_n246), .B1(new_n824), .B2(new_n826), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n823), .B(new_n832), .C1(new_n830), .C2(new_n831), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n671), .A2(new_n585), .A3(new_n673), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n744), .B2(new_n745), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n835), .A2(KEYINPUT115), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n826), .A2(new_n739), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(KEYINPUT115), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n687), .A2(new_n639), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT111), .B1(new_n829), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n829), .A2(KEYINPUT111), .A3(new_n840), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n300), .A2(new_n607), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n672), .A2(new_n673), .A3(new_n303), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n846), .A2(KEYINPUT109), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(KEYINPUT109), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n658), .A2(new_n826), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT50), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n849), .A2(KEYINPUT50), .A3(new_n850), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n822), .A2(new_n845), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n844), .A2(KEYINPUT114), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT114), .B1(new_n844), .B2(new_n855), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n839), .B(KEYINPUT51), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n843), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n841), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n822), .A2(new_n845), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n853), .A2(new_n854), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT113), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n844), .A2(new_n865), .A3(new_n855), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n834), .B(KEYINPUT108), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n837), .B1(new_n746), .B2(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n864), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  XOR2_X1   g683(.A(KEYINPUT107), .B(KEYINPUT51), .Z(new_n870));
  OAI211_X1 g684(.A(new_n833), .B(new_n858), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n816), .A2(new_n871), .B1(G952), .B2(G953), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n672), .A2(KEYINPUT49), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT102), .Z(new_n874));
  NAND3_X1  g688(.A1(new_n448), .A2(new_n731), .A3(new_n701), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT101), .Z(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(KEYINPUT49), .B2(new_n672), .ZN(new_n877));
  INV_X1    g691(.A(new_n658), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n818), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n872), .B1(new_n874), .B2(new_n879), .ZN(G75));
  NAND2_X1  g694(.A1(new_n241), .A2(new_n306), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n789), .B2(new_n813), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n350), .A2(new_n376), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(new_n374), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT55), .Z(new_n885));
  NOR3_X1   g699(.A1(new_n882), .A2(KEYINPUT56), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n245), .A2(G952), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n882), .A2(KEYINPUT117), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n882), .B2(KEYINPUT117), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n885), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT118), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n885), .C1(new_n890), .C2(new_n892), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n888), .B1(new_n894), .B2(new_n896), .ZN(G51));
  INV_X1    g711(.A(new_n813), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT54), .B1(new_n898), .B2(new_n804), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(KEYINPUT119), .A3(new_n815), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n789), .A2(new_n813), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT54), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n724), .B(KEYINPUT57), .Z(new_n904));
  NAND3_X1  g718(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n583), .B2(new_n584), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n901), .A2(new_n241), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n907), .A2(new_n723), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n887), .B1(new_n906), .B2(new_n908), .ZN(G54));
  NAND4_X1  g723(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .A4(new_n241), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n294), .A2(new_n283), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n910), .A2(new_n912), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n887), .ZN(G60));
  XNOR2_X1  g729(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n233), .A2(new_n254), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n815), .B1(new_n801), .B2(KEYINPUT105), .ZN(new_n920));
  INV_X1    g734(.A(new_n805), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n602), .A2(new_n603), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n887), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n918), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n900), .A2(new_n903), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT121), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n900), .A2(new_n928), .A3(new_n903), .A4(new_n925), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n924), .A2(new_n930), .ZN(G63));
  XOR2_X1   g745(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n225), .A2(new_n254), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n898), .B2(new_n804), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n887), .B1(new_n936), .B2(new_n439), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n901), .A2(new_n631), .A3(new_n935), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n937), .B2(new_n938), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n932), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n937), .A2(KEYINPUT61), .A3(new_n940), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(G66));
  NOR3_X1   g758(.A1(new_n252), .A2(new_n372), .A3(new_n245), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n797), .A2(new_n798), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n793), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n945), .B1(new_n948), .B2(new_n245), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n883), .B1(G898), .B2(new_n245), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G69));
  NOR2_X1   g765(.A1(new_n753), .A2(new_n667), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n662), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n955));
  NOR4_X1   g769(.A1(new_n649), .A2(new_n711), .A3(new_n739), .A4(new_n783), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n741), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n959), .A2(G953), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n954), .A2(new_n749), .A3(new_n955), .A4(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n472), .A2(new_n476), .A3(new_n483), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(new_n290), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n807), .B1(new_n746), .B2(new_n748), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n741), .A2(new_n716), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n730), .A2(new_n706), .A3(new_n756), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n952), .ZN(new_n970));
  OR3_X1    g784(.A1(new_n969), .A2(KEYINPUT126), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(KEYINPUT126), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(new_n245), .A3(new_n972), .ZN(new_n973));
  OR3_X1    g787(.A1(new_n642), .A2(KEYINPUT127), .A3(G227), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n245), .B1(KEYINPUT127), .B2(new_n642), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n965), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI22_X1  g790(.A1(new_n963), .A2(new_n965), .B1(new_n973), .B2(new_n976), .ZN(G72));
  NOR2_X1   g791(.A1(new_n959), .A2(new_n947), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n954), .A2(new_n749), .A3(new_n955), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(G472), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT63), .Z(new_n981));
  AOI211_X1 g795(.A(new_n490), .B(new_n652), .C1(new_n979), .C2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n652), .A2(new_n490), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n971), .A2(new_n948), .A3(new_n972), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n981), .ZN(new_n985));
  INV_X1    g799(.A(new_n492), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n981), .B1(new_n986), .B2(new_n525), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n789), .B2(new_n800), .ZN(new_n988));
  NOR4_X1   g802(.A1(new_n982), .A2(new_n985), .A3(new_n887), .A4(new_n988), .ZN(G57));
endmodule


