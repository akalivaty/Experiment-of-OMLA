

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748;

  XNOR2_X1 U374 ( .A(n482), .B(G134), .ZN(n467) );
  INV_X2 U375 ( .A(G128), .ZN(n374) );
  INV_X2 U376 ( .A(G953), .ZN(n736) );
  XNOR2_X1 U377 ( .A(KEYINPUT24), .B(G110), .ZN(n381) );
  AND2_X2 U378 ( .A1(n568), .A2(n567), .ZN(n639) );
  XNOR2_X2 U379 ( .A(n447), .B(n424), .ZN(n695) );
  XNOR2_X2 U380 ( .A(n735), .B(G146), .ZN(n447) );
  XNOR2_X2 U381 ( .A(n544), .B(KEYINPUT114), .ZN(n746) );
  NOR2_X1 U382 ( .A1(n745), .A2(n748), .ZN(n560) );
  XNOR2_X1 U383 ( .A(KEYINPUT23), .B(KEYINPUT81), .ZN(n382) );
  INV_X1 U384 ( .A(KEYINPUT30), .ZN(n451) );
  XNOR2_X1 U385 ( .A(n378), .B(n357), .ZN(n745) );
  NOR2_X1 U386 ( .A1(n554), .A2(n557), .ZN(n556) );
  XNOR2_X1 U387 ( .A(n399), .B(n402), .ZN(n454) );
  XNOR2_X1 U388 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U389 ( .A(n382), .B(n381), .ZN(n380) );
  XNOR2_X1 U390 ( .A(n578), .B(KEYINPUT35), .ZN(n638) );
  NOR2_X2 U391 ( .A1(n640), .A2(n613), .ZN(n617) );
  XNOR2_X1 U392 ( .A(n474), .B(G478), .ZN(n499) );
  NOR2_X1 U393 ( .A1(n719), .A2(G902), .ZN(n474) );
  XNOR2_X1 U394 ( .A(n398), .B(n734), .ZN(n689) );
  XNOR2_X1 U395 ( .A(n384), .B(n379), .ZN(n398) );
  XNOR2_X1 U396 ( .A(n383), .B(n380), .ZN(n379) );
  XNOR2_X1 U397 ( .A(n467), .B(n417), .ZN(n735) );
  XNOR2_X1 U398 ( .A(G146), .B(G125), .ZN(n484) );
  INV_X1 U399 ( .A(G237), .ZN(n434) );
  INV_X1 U400 ( .A(n493), .ZN(n365) );
  XNOR2_X1 U401 ( .A(n526), .B(KEYINPUT1), .ZN(n570) );
  BUF_X1 U402 ( .A(n639), .Z(n641) );
  XNOR2_X1 U403 ( .A(n439), .B(n392), .ZN(n455) );
  INV_X1 U404 ( .A(KEYINPUT75), .ZN(n392) );
  NOR2_X1 U405 ( .A1(G953), .A2(G237), .ZN(n439) );
  XNOR2_X1 U406 ( .A(n484), .B(KEYINPUT10), .ZN(n458) );
  XNOR2_X1 U407 ( .A(n395), .B(n394), .ZN(n393) );
  XNOR2_X1 U408 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n394) );
  XNOR2_X1 U409 ( .A(n456), .B(KEYINPUT105), .ZN(n395) );
  XNOR2_X1 U410 ( .A(G143), .B(G140), .ZN(n456) );
  INV_X1 U411 ( .A(G140), .ZN(n404) );
  NOR2_X1 U412 ( .A1(n589), .A2(KEYINPUT34), .ZN(n373) );
  BUF_X1 U413 ( .A(n570), .Z(n649) );
  XNOR2_X1 U414 ( .A(n502), .B(n501), .ZN(n602) );
  XNOR2_X1 U415 ( .A(n458), .B(n419), .ZN(n734) );
  NAND2_X1 U416 ( .A1(G234), .A2(G237), .ZN(n427) );
  XOR2_X1 U417 ( .A(KEYINPUT38), .B(n553), .Z(n557) );
  INV_X1 U418 ( .A(n509), .ZN(n401) );
  XNOR2_X1 U419 ( .A(n588), .B(KEYINPUT110), .ZN(n400) );
  INV_X1 U420 ( .A(KEYINPUT76), .ZN(n402) );
  XNOR2_X1 U421 ( .A(n450), .B(n449), .ZN(n511) );
  XNOR2_X1 U422 ( .A(n359), .B(n478), .ZN(n723) );
  XNOR2_X1 U423 ( .A(n476), .B(n475), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n407), .B(n385), .ZN(n471) );
  XNOR2_X1 U425 ( .A(n467), .B(n468), .ZN(n469) );
  NAND2_X1 U426 ( .A1(n386), .A2(n641), .ZN(n388) );
  NOR2_X1 U427 ( .A1(n640), .A2(KEYINPUT83), .ZN(n386) );
  NAND2_X1 U428 ( .A1(KEYINPUT2), .A2(n389), .ZN(n387) );
  NAND2_X1 U429 ( .A1(n641), .A2(n642), .ZN(n643) );
  XNOR2_X1 U430 ( .A(n558), .B(KEYINPUT41), .ZN(n678) );
  NAND2_X1 U431 ( .A1(n362), .A2(n355), .ZN(n361) );
  OR2_X1 U432 ( .A1(n662), .A2(n365), .ZN(n364) );
  INV_X1 U433 ( .A(n499), .ZN(n532) );
  BUF_X1 U434 ( .A(n511), .Z(n656) );
  XNOR2_X1 U435 ( .A(n641), .B(n738), .ZN(n737) );
  XNOR2_X1 U436 ( .A(n393), .B(n391), .ZN(n461) );
  NAND2_X1 U437 ( .A1(n455), .A2(G214), .ZN(n391) );
  AND2_X1 U438 ( .A1(n622), .A2(G953), .ZN(n722) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n748) );
  INV_X1 U440 ( .A(KEYINPUT42), .ZN(n376) );
  OR2_X1 U441 ( .A1(n678), .A2(n559), .ZN(n377) );
  NOR2_X1 U442 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U443 ( .A1(n372), .A2(n370), .ZN(n578) );
  NAND2_X1 U444 ( .A1(n371), .A2(n373), .ZN(n370) );
  AND2_X1 U445 ( .A1(n369), .A2(n352), .ZN(n372) );
  NAND2_X1 U446 ( .A1(n602), .A2(n520), .ZN(n358) );
  INV_X1 U447 ( .A(G143), .ZN(n492) );
  XNOR2_X1 U448 ( .A(n464), .B(n463), .ZN(n533) );
  INV_X1 U449 ( .A(n533), .ZN(n396) );
  AND2_X1 U450 ( .A1(n368), .A2(n577), .ZN(n352) );
  INV_X1 U451 ( .A(n553), .ZN(n362) );
  AND2_X1 U452 ( .A1(n606), .A2(n699), .ZN(n353) );
  NOR2_X1 U453 ( .A1(n505), .A2(n522), .ZN(n354) );
  AND2_X1 U454 ( .A1(n662), .A2(n365), .ZN(n355) );
  XNOR2_X1 U455 ( .A(n498), .B(KEYINPUT65), .ZN(n356) );
  XOR2_X1 U456 ( .A(KEYINPUT40), .B(KEYINPUT112), .Z(n357) );
  INV_X1 U457 ( .A(KEYINPUT83), .ZN(n389) );
  INV_X1 U458 ( .A(KEYINPUT2), .ZN(n390) );
  NAND2_X1 U459 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U460 ( .A1(n602), .A2(n354), .ZN(n579) );
  XNOR2_X2 U461 ( .A(n358), .B(KEYINPUT32), .ZN(n580) );
  XNOR2_X2 U462 ( .A(n360), .B(n444), .ZN(n476) );
  XNOR2_X2 U463 ( .A(n443), .B(n442), .ZN(n360) );
  NAND2_X1 U464 ( .A1(n362), .A2(n662), .ZN(n539) );
  NAND2_X1 U465 ( .A1(n363), .A2(n361), .ZN(n529) );
  AND2_X1 U466 ( .A1(n366), .A2(n364), .ZN(n363) );
  NAND2_X1 U467 ( .A1(n553), .A2(n493), .ZN(n366) );
  XNOR2_X2 U468 ( .A(n367), .B(n356), .ZN(n594) );
  OR2_X2 U469 ( .A1(n529), .A2(n497), .ZN(n367) );
  NAND2_X1 U470 ( .A1(n589), .A2(KEYINPUT34), .ZN(n368) );
  NAND2_X1 U471 ( .A1(n661), .A2(KEYINPUT34), .ZN(n369) );
  XNOR2_X1 U472 ( .A(n576), .B(n575), .ZN(n661) );
  INV_X1 U473 ( .A(n661), .ZN(n371) );
  XNOR2_X2 U474 ( .A(n374), .B(G143), .ZN(n482) );
  NOR2_X2 U475 ( .A1(n375), .A2(n526), .ZN(n588) );
  NOR2_X1 U476 ( .A1(n570), .A2(n375), .ZN(n571) );
  NAND2_X1 U477 ( .A1(n649), .A2(n375), .ZN(n650) );
  XNOR2_X2 U478 ( .A(n416), .B(KEYINPUT66), .ZN(n375) );
  NAND2_X1 U479 ( .A1(n565), .A2(n711), .ZN(n378) );
  XNOR2_X1 U480 ( .A(n556), .B(n555), .ZN(n565) );
  XNOR2_X1 U481 ( .A(n406), .B(n405), .ZN(n383) );
  NAND2_X1 U482 ( .A1(n471), .A2(G221), .ZN(n384) );
  NAND2_X1 U483 ( .A1(n736), .A2(G234), .ZN(n385) );
  NAND2_X1 U484 ( .A1(n388), .A2(n387), .ZN(n645) );
  NOR2_X1 U485 ( .A1(n523), .A2(n397), .ZN(n513) );
  NAND2_X1 U486 ( .A1(n396), .A2(n499), .ZN(n397) );
  INV_X1 U487 ( .A(n397), .ZN(n711) );
  NAND2_X1 U488 ( .A1(n400), .A2(n401), .ZN(n399) );
  BUF_X1 U489 ( .A(n688), .Z(n718) );
  XOR2_X1 U490 ( .A(KEYINPUT28), .B(KEYINPUT111), .Z(n403) );
  INV_X1 U491 ( .A(KEYINPUT90), .ZN(n581) );
  INV_X1 U492 ( .A(KEYINPUT44), .ZN(n585) );
  BUF_X1 U493 ( .A(n661), .Z(n679) );
  INV_X1 U494 ( .A(KEYINPUT113), .ZN(n537) );
  XNOR2_X1 U495 ( .A(n538), .B(n537), .ZN(n540) );
  INV_X1 U496 ( .A(G107), .ZN(n468) );
  INV_X1 U497 ( .A(KEYINPUT39), .ZN(n555) );
  XNOR2_X1 U498 ( .A(n404), .B(G137), .ZN(n419) );
  XNOR2_X1 U499 ( .A(KEYINPUT98), .B(KEYINPUT97), .ZN(n405) );
  XNOR2_X1 U500 ( .A(G119), .B(G128), .ZN(n406) );
  XOR2_X1 U501 ( .A(KEYINPUT82), .B(KEYINPUT8), .Z(n407) );
  INV_X1 U502 ( .A(G902), .ZN(n448) );
  NAND2_X1 U503 ( .A1(n689), .A2(n448), .ZN(n413) );
  XOR2_X1 U504 ( .A(KEYINPUT20), .B(KEYINPUT99), .Z(n409) );
  XNOR2_X1 U505 ( .A(G902), .B(KEYINPUT15), .ZN(n614) );
  NAND2_X1 U506 ( .A1(G234), .A2(n614), .ZN(n408) );
  XNOR2_X1 U507 ( .A(n409), .B(n408), .ZN(n414) );
  NAND2_X1 U508 ( .A1(n414), .A2(G217), .ZN(n411) );
  XOR2_X1 U509 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n410) );
  XNOR2_X1 U510 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X2 U511 ( .A(n413), .B(n412), .ZN(n507) );
  NAND2_X1 U512 ( .A1(n414), .A2(G221), .ZN(n415) );
  XNOR2_X1 U513 ( .A(n415), .B(KEYINPUT21), .ZN(n506) );
  INV_X1 U514 ( .A(n506), .ZN(n651) );
  NAND2_X1 U515 ( .A1(n507), .A2(n651), .ZN(n416) );
  XNOR2_X1 U516 ( .A(KEYINPUT4), .B(G131), .ZN(n417) );
  NAND2_X1 U517 ( .A1(G227), .A2(n736), .ZN(n418) );
  XNOR2_X1 U518 ( .A(n418), .B(G104), .ZN(n420) );
  XNOR2_X1 U519 ( .A(n420), .B(n419), .ZN(n423) );
  XNOR2_X1 U520 ( .A(G107), .B(G101), .ZN(n422) );
  XNOR2_X1 U521 ( .A(KEYINPUT94), .B(G110), .ZN(n421) );
  XNOR2_X1 U522 ( .A(n422), .B(n421), .ZN(n477) );
  XNOR2_X1 U523 ( .A(n423), .B(n477), .ZN(n424) );
  NAND2_X1 U524 ( .A1(n695), .A2(n448), .ZN(n426) );
  XOR2_X1 U525 ( .A(KEYINPUT68), .B(G469), .Z(n425) );
  XNOR2_X2 U526 ( .A(n426), .B(n425), .ZN(n526) );
  XOR2_X1 U527 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n428) );
  XNOR2_X1 U528 ( .A(n428), .B(n427), .ZN(n429) );
  NAND2_X1 U529 ( .A1(G952), .A2(n429), .ZN(n677) );
  NOR2_X1 U530 ( .A1(n677), .A2(G953), .ZN(n495) );
  NAND2_X1 U531 ( .A1(G902), .A2(n429), .ZN(n430) );
  XOR2_X1 U532 ( .A(KEYINPUT96), .B(n430), .Z(n431) );
  NAND2_X1 U533 ( .A1(G953), .A2(n431), .ZN(n494) );
  NOR2_X1 U534 ( .A1(G900), .A2(n494), .ZN(n432) );
  XNOR2_X1 U535 ( .A(n432), .B(KEYINPUT108), .ZN(n433) );
  NOR2_X1 U536 ( .A1(n495), .A2(n433), .ZN(n509) );
  NAND2_X1 U537 ( .A1(n448), .A2(n434), .ZN(n488) );
  NAND2_X1 U538 ( .A1(n488), .A2(G214), .ZN(n662) );
  XOR2_X1 U539 ( .A(G113), .B(G137), .Z(n436) );
  XNOR2_X1 U540 ( .A(KEYINPUT100), .B(KEYINPUT5), .ZN(n435) );
  XNOR2_X1 U541 ( .A(n436), .B(n435), .ZN(n438) );
  INV_X1 U542 ( .A(G101), .ZN(n437) );
  XNOR2_X1 U543 ( .A(n438), .B(n437), .ZN(n441) );
  NAND2_X1 U544 ( .A1(n455), .A2(G210), .ZN(n440) );
  XNOR2_X1 U545 ( .A(n441), .B(n440), .ZN(n445) );
  XNOR2_X2 U546 ( .A(KEYINPUT3), .B(G119), .ZN(n443) );
  XNOR2_X2 U547 ( .A(G116), .B(KEYINPUT69), .ZN(n442) );
  XNOR2_X1 U548 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n444) );
  XNOR2_X1 U549 ( .A(n445), .B(n476), .ZN(n446) );
  XNOR2_X1 U550 ( .A(n447), .B(n446), .ZN(n619) );
  NAND2_X1 U551 ( .A1(n619), .A2(n448), .ZN(n450) );
  XOR2_X1 U552 ( .A(G472), .B(KEYINPUT101), .Z(n449) );
  XNOR2_X1 U553 ( .A(n511), .B(KEYINPUT106), .ZN(n522) );
  NAND2_X1 U554 ( .A1(n662), .A2(n522), .ZN(n452) );
  NAND2_X1 U555 ( .A1(n454), .A2(n453), .ZN(n554) );
  XNOR2_X1 U556 ( .A(G122), .B(G113), .ZN(n457) );
  XNOR2_X1 U557 ( .A(n457), .B(G104), .ZN(n475) );
  XNOR2_X1 U558 ( .A(n475), .B(G131), .ZN(n459) );
  XNOR2_X1 U559 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U560 ( .A(n461), .B(n460), .ZN(n633) );
  NOR2_X1 U561 ( .A1(G902), .A2(n633), .ZN(n462) );
  XNOR2_X1 U562 ( .A(G475), .B(n462), .ZN(n464) );
  INV_X1 U563 ( .A(KEYINPUT13), .ZN(n463) );
  XNOR2_X1 U564 ( .A(G116), .B(G122), .ZN(n465) );
  XNOR2_X1 U565 ( .A(n465), .B(KEYINPUT7), .ZN(n466) );
  XOR2_X1 U566 ( .A(n466), .B(KEYINPUT9), .Z(n470) );
  XNOR2_X1 U567 ( .A(n470), .B(n469), .ZN(n473) );
  NAND2_X1 U568 ( .A1(G217), .A2(n471), .ZN(n472) );
  XOR2_X1 U569 ( .A(n473), .B(n472), .Z(n719) );
  AND2_X1 U570 ( .A1(n396), .A2(n532), .ZN(n577) );
  XNOR2_X1 U571 ( .A(n477), .B(KEYINPUT16), .ZN(n478) );
  XNOR2_X1 U572 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n480) );
  NAND2_X1 U573 ( .A1(n736), .A2(G224), .ZN(n479) );
  XNOR2_X1 U574 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U575 ( .A(n482), .B(n481), .ZN(n486) );
  XNOR2_X1 U576 ( .A(KEYINPUT95), .B(KEYINPUT4), .ZN(n483) );
  XNOR2_X1 U577 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U578 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U579 ( .A(n723), .B(n487), .ZN(n627) );
  INV_X1 U580 ( .A(n614), .ZN(n612) );
  OR2_X2 U581 ( .A1(n627), .A2(n612), .ZN(n490) );
  NAND2_X1 U582 ( .A1(n488), .A2(G210), .ZN(n489) );
  XNOR2_X2 U583 ( .A(n490), .B(n489), .ZN(n553) );
  NAND2_X1 U584 ( .A1(n577), .A2(n362), .ZN(n491) );
  NOR2_X1 U585 ( .A1(n554), .A2(n491), .ZN(n547) );
  XNOR2_X1 U586 ( .A(n547), .B(n492), .ZN(G45) );
  XNOR2_X1 U587 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n493) );
  NOR2_X1 U588 ( .A1(n494), .A2(G898), .ZN(n496) );
  NOR2_X1 U589 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U590 ( .A(KEYINPUT92), .B(KEYINPUT0), .ZN(n498) );
  NAND2_X1 U591 ( .A1(n533), .A2(n499), .ZN(n665) );
  NOR2_X1 U592 ( .A1(n665), .A2(n506), .ZN(n500) );
  NAND2_X1 U593 ( .A1(n594), .A2(n500), .ZN(n502) );
  INV_X1 U594 ( .A(KEYINPUT22), .ZN(n501) );
  BUF_X1 U595 ( .A(n507), .Z(n503) );
  INV_X1 U596 ( .A(n503), .ZN(n504) );
  NAND2_X1 U597 ( .A1(n649), .A2(n504), .ZN(n505) );
  XNOR2_X1 U598 ( .A(n579), .B(G110), .ZN(G12) );
  INV_X1 U599 ( .A(n649), .ZN(n542) );
  OR2_X1 U600 ( .A1(n507), .A2(n506), .ZN(n508) );
  NOR2_X1 U601 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U602 ( .A(KEYINPUT67), .B(n510), .ZN(n523) );
  INV_X1 U603 ( .A(KEYINPUT6), .ZN(n512) );
  XNOR2_X1 U604 ( .A(n656), .B(n512), .ZN(n518) );
  NAND2_X1 U605 ( .A1(n513), .A2(n518), .ZN(n538) );
  NOR2_X1 U606 ( .A1(n542), .A2(n538), .ZN(n514) );
  NAND2_X1 U607 ( .A1(n662), .A2(n514), .ZN(n515) );
  XNOR2_X1 U608 ( .A(n515), .B(KEYINPUT43), .ZN(n516) );
  XOR2_X1 U609 ( .A(n516), .B(KEYINPUT109), .Z(n517) );
  NAND2_X1 U610 ( .A1(n517), .A2(n553), .ZN(n566) );
  XNOR2_X1 U611 ( .A(n566), .B(G140), .ZN(G42) );
  XNOR2_X1 U612 ( .A(G119), .B(KEYINPUT127), .ZN(n521) );
  INV_X1 U613 ( .A(n518), .ZN(n601) );
  NOR2_X1 U614 ( .A1(n649), .A2(n503), .ZN(n519) );
  AND2_X1 U615 ( .A1(n601), .A2(n519), .ZN(n520) );
  XOR2_X1 U616 ( .A(n521), .B(n580), .Z(G21) );
  INV_X1 U617 ( .A(n522), .ZN(n524) );
  NOR2_X1 U618 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U619 ( .A(n525), .B(n403), .ZN(n528) );
  INV_X1 U620 ( .A(n526), .ZN(n527) );
  NAND2_X1 U621 ( .A1(n528), .A2(n527), .ZN(n559) );
  NOR2_X1 U622 ( .A1(n559), .A2(n529), .ZN(n708) );
  INV_X1 U623 ( .A(KEYINPUT47), .ZN(n530) );
  NOR2_X1 U624 ( .A1(n708), .A2(n530), .ZN(n531) );
  XOR2_X1 U625 ( .A(n531), .B(KEYINPUT80), .Z(n536) );
  AND2_X1 U626 ( .A1(n533), .A2(n532), .ZN(n713) );
  NOR2_X1 U627 ( .A1(n711), .A2(n713), .ZN(n667) );
  NOR2_X1 U628 ( .A1(n667), .A2(KEYINPUT47), .ZN(n534) );
  NAND2_X1 U629 ( .A1(n708), .A2(n534), .ZN(n535) );
  NAND2_X1 U630 ( .A1(n536), .A2(n535), .ZN(n546) );
  XNOR2_X1 U631 ( .A(n541), .B(KEYINPUT36), .ZN(n543) );
  NAND2_X1 U632 ( .A1(n543), .A2(n542), .ZN(n544) );
  INV_X1 U633 ( .A(n746), .ZN(n545) );
  NOR2_X1 U634 ( .A1(n546), .A2(n545), .ZN(n552) );
  INV_X1 U635 ( .A(n547), .ZN(n549) );
  NAND2_X1 U636 ( .A1(n667), .A2(KEYINPUT47), .ZN(n548) );
  NAND2_X1 U637 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U638 ( .A(n550), .B(KEYINPUT79), .ZN(n551) );
  AND2_X1 U639 ( .A1(n552), .A2(n551), .ZN(n562) );
  INV_X1 U640 ( .A(n557), .ZN(n663) );
  NAND2_X1 U641 ( .A1(n663), .A2(n662), .ZN(n666) );
  NOR2_X1 U642 ( .A1(n665), .A2(n666), .ZN(n558) );
  XNOR2_X1 U643 ( .A(n560), .B(KEYINPUT46), .ZN(n561) );
  NAND2_X1 U644 ( .A1(n562), .A2(n561), .ZN(n564) );
  XOR2_X1 U645 ( .A(KEYINPUT88), .B(KEYINPUT48), .Z(n563) );
  XNOR2_X1 U646 ( .A(n564), .B(n563), .ZN(n568) );
  NAND2_X1 U647 ( .A1(n713), .A2(n565), .ZN(n717) );
  AND2_X1 U648 ( .A1(n566), .A2(n717), .ZN(n567) );
  NAND2_X1 U649 ( .A1(n639), .A2(KEYINPUT2), .ZN(n569) );
  XNOR2_X1 U650 ( .A(n569), .B(KEYINPUT86), .ZN(n611) );
  XNOR2_X1 U651 ( .A(n571), .B(KEYINPUT74), .ZN(n592) );
  XNOR2_X1 U652 ( .A(n592), .B(KEYINPUT107), .ZN(n572) );
  NOR2_X1 U653 ( .A1(n572), .A2(n601), .ZN(n576) );
  XNOR2_X1 U654 ( .A(KEYINPUT93), .B(KEYINPUT33), .ZN(n574) );
  INV_X1 U655 ( .A(KEYINPUT72), .ZN(n573) );
  XNOR2_X1 U656 ( .A(n574), .B(n573), .ZN(n575) );
  INV_X1 U657 ( .A(n594), .ZN(n589) );
  INV_X1 U658 ( .A(n638), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n582), .B(n581), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U661 ( .A(n586), .B(n585), .ZN(n607) );
  INV_X1 U662 ( .A(n656), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n588), .A2(n587), .ZN(n590) );
  NOR2_X1 U664 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U665 ( .A(KEYINPUT102), .B(n591), .ZN(n701) );
  NAND2_X1 U666 ( .A1(n592), .A2(n656), .ZN(n593) );
  XNOR2_X1 U667 ( .A(n593), .B(KEYINPUT103), .ZN(n658) );
  AND2_X1 U668 ( .A1(n658), .A2(n594), .ZN(n596) );
  INV_X1 U669 ( .A(KEYINPUT31), .ZN(n595) );
  XNOR2_X1 U670 ( .A(n596), .B(n595), .ZN(n714) );
  NOR2_X1 U671 ( .A1(n701), .A2(n714), .ZN(n598) );
  INV_X1 U672 ( .A(KEYINPUT104), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n598), .B(n597), .ZN(n600) );
  INV_X1 U674 ( .A(n667), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n606) );
  AND2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n603), .A2(n649), .ZN(n604) );
  XNOR2_X1 U678 ( .A(n604), .B(KEYINPUT89), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n605), .A2(n503), .ZN(n699) );
  NAND2_X1 U680 ( .A1(n607), .A2(n353), .ZN(n610) );
  INV_X1 U681 ( .A(KEYINPUT64), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n608), .B(KEYINPUT45), .ZN(n609) );
  XNOR2_X2 U683 ( .A(n610), .B(n609), .ZN(n640) );
  NOR2_X1 U684 ( .A1(n611), .A2(n640), .ZN(n646) );
  NAND2_X1 U685 ( .A1(n639), .A2(n612), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT85), .ZN(n615) );
  AND2_X1 U687 ( .A1(n615), .A2(KEYINPUT2), .ZN(n616) );
  NOR2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X2 U689 ( .A1(n646), .A2(n618), .ZN(n688) );
  NAND2_X1 U690 ( .A1(n688), .A2(G472), .ZN(n621) );
  XOR2_X1 U691 ( .A(KEYINPUT62), .B(n619), .Z(n620) );
  XNOR2_X1 U692 ( .A(n621), .B(n620), .ZN(n623) );
  INV_X1 U693 ( .A(G952), .ZN(n622) );
  NOR2_X2 U694 ( .A1(n623), .A2(n722), .ZN(n625) );
  XNOR2_X1 U695 ( .A(KEYINPUT91), .B(KEYINPUT63), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(G57) );
  NAND2_X1 U697 ( .A1(n688), .A2(G210), .ZN(n629) );
  XOR2_X1 U698 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n626) );
  XNOR2_X1 U699 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n629), .B(n628), .ZN(n630) );
  NOR2_X2 U701 ( .A1(n630), .A2(n722), .ZN(n632) );
  XOR2_X1 U702 ( .A(KEYINPUT87), .B(KEYINPUT56), .Z(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(G51) );
  NAND2_X1 U704 ( .A1(n688), .A2(G475), .ZN(n635) );
  XOR2_X1 U705 ( .A(KEYINPUT59), .B(n633), .Z(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X2 U707 ( .A1(n636), .A2(n722), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n637), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U709 ( .A(n638), .B(G122), .Z(G24) );
  INV_X1 U710 ( .A(n640), .ZN(n726) );
  AND2_X1 U711 ( .A1(n390), .A2(KEYINPUT83), .ZN(n642) );
  NOR2_X1 U712 ( .A1(n726), .A2(n643), .ZN(n644) );
  NOR2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n647) );
  NOR2_X1 U714 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U715 ( .A(n648), .B(KEYINPUT84), .ZN(n686) );
  XNOR2_X1 U716 ( .A(n650), .B(KEYINPUT50), .ZN(n654) );
  NOR2_X1 U717 ( .A1(n651), .A2(n503), .ZN(n652) );
  XNOR2_X1 U718 ( .A(n652), .B(KEYINPUT49), .ZN(n653) );
  NAND2_X1 U719 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U721 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U722 ( .A(KEYINPUT51), .B(n659), .Z(n660) );
  NOR2_X1 U723 ( .A1(n678), .A2(n660), .ZN(n673) );
  NOR2_X1 U724 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U725 ( .A1(n665), .A2(n664), .ZN(n670) );
  NOR2_X1 U726 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U727 ( .A(n668), .B(KEYINPUT118), .ZN(n669) );
  NOR2_X1 U728 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U729 ( .A1(n679), .A2(n671), .ZN(n672) );
  NOR2_X1 U730 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U731 ( .A(n674), .B(KEYINPUT119), .Z(n675) );
  XNOR2_X1 U732 ( .A(KEYINPUT52), .B(n675), .ZN(n676) );
  NOR2_X1 U733 ( .A1(n677), .A2(n676), .ZN(n682) );
  NOR2_X1 U734 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U735 ( .A(n680), .B(KEYINPUT120), .ZN(n681) );
  OR2_X1 U736 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U737 ( .A(n683), .B(KEYINPUT121), .ZN(n684) );
  NAND2_X1 U738 ( .A1(n684), .A2(n736), .ZN(n685) );
  NOR2_X1 U739 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U740 ( .A(n687), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U741 ( .A1(n718), .A2(G217), .ZN(n692) );
  BUF_X1 U742 ( .A(n689), .Z(n690) );
  XOR2_X1 U743 ( .A(KEYINPUT122), .B(n690), .Z(n691) );
  XNOR2_X1 U744 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U745 ( .A1(n693), .A2(n722), .ZN(G66) );
  NAND2_X1 U746 ( .A1(n718), .A2(G469), .ZN(n697) );
  XNOR2_X1 U747 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n694) );
  XNOR2_X1 U748 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U749 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U750 ( .A1(n698), .A2(n722), .ZN(G54) );
  XNOR2_X1 U751 ( .A(G101), .B(n699), .ZN(G3) );
  NAND2_X1 U752 ( .A1(n701), .A2(n711), .ZN(n700) );
  XNOR2_X1 U753 ( .A(n700), .B(G104), .ZN(G6) );
  XOR2_X1 U754 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n703) );
  NAND2_X1 U755 ( .A1(n713), .A2(n701), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U757 ( .A(G107), .B(n704), .ZN(G9) );
  XOR2_X1 U758 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n706) );
  NAND2_X1 U759 ( .A1(n708), .A2(n713), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(n707) );
  XOR2_X1 U761 ( .A(G128), .B(n707), .Z(G30) );
  NAND2_X1 U762 ( .A1(n708), .A2(n711), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n709), .B(KEYINPUT116), .ZN(n710) );
  XNOR2_X1 U764 ( .A(G146), .B(n710), .ZN(G48) );
  NAND2_X1 U765 ( .A1(n714), .A2(n711), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n712), .B(G113), .ZN(G15) );
  NAND2_X1 U767 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n715), .B(G116), .ZN(G18) );
  XOR2_X1 U769 ( .A(G134), .B(KEYINPUT117), .Z(n716) );
  XNOR2_X1 U770 ( .A(n717), .B(n716), .ZN(G36) );
  NAND2_X1 U771 ( .A1(n718), .A2(G478), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U773 ( .A1(n722), .A2(n721), .ZN(G63) );
  XNOR2_X1 U774 ( .A(n723), .B(KEYINPUT124), .ZN(n725) );
  NOR2_X1 U775 ( .A1(G898), .A2(n736), .ZN(n724) );
  NOR2_X1 U776 ( .A1(n725), .A2(n724), .ZN(n733) );
  NAND2_X1 U777 ( .A1(n726), .A2(n736), .ZN(n731) );
  XOR2_X1 U778 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n728) );
  NAND2_X1 U779 ( .A1(G224), .A2(G953), .ZN(n727) );
  XNOR2_X1 U780 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U781 ( .A1(n729), .A2(G898), .ZN(n730) );
  NAND2_X1 U782 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U783 ( .A(n733), .B(n732), .ZN(G69) );
  XNOR2_X1 U784 ( .A(n735), .B(n734), .ZN(n738) );
  NAND2_X1 U785 ( .A1(n737), .A2(n736), .ZN(n744) );
  XNOR2_X1 U786 ( .A(n738), .B(G227), .ZN(n739) );
  XNOR2_X1 U787 ( .A(n739), .B(KEYINPUT125), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n740), .A2(G900), .ZN(n741) );
  XNOR2_X1 U789 ( .A(KEYINPUT126), .B(n741), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n742), .A2(G953), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n744), .A2(n743), .ZN(G72) );
  XOR2_X1 U792 ( .A(n745), .B(G131), .Z(G33) );
  XOR2_X1 U793 ( .A(G125), .B(n746), .Z(n747) );
  XNOR2_X1 U794 ( .A(KEYINPUT37), .B(n747), .ZN(G27) );
  XOR2_X1 U795 ( .A(n748), .B(G137), .Z(G39) );
endmodule

