

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772;

  XNOR2_X1 U376 ( .A(n511), .B(n752), .ZN(n520) );
  INV_X1 U377 ( .A(G953), .ZN(n766) );
  AND2_X1 U378 ( .A1(n640), .A2(n726), .ZN(n628) );
  XNOR2_X2 U379 ( .A(n632), .B(KEYINPUT42), .ZN(n770) );
  NOR2_X2 U380 ( .A1(n661), .A2(KEYINPUT44), .ZN(n554) );
  NOR2_X2 U381 ( .A1(n638), .A2(n429), .ZN(n428) );
  INV_X2 U382 ( .A(n681), .ZN(n354) );
  XNOR2_X2 U383 ( .A(n382), .B(n480), .ZN(n505) );
  XNOR2_X2 U384 ( .A(G143), .B(G128), .ZN(n382) );
  XNOR2_X2 U385 ( .A(n514), .B(G472), .ZN(n601) );
  NOR2_X2 U386 ( .A1(n729), .A2(n726), .ZN(n695) );
  XNOR2_X2 U387 ( .A(n566), .B(n425), .ZN(n726) );
  AND2_X1 U388 ( .A1(n641), .A2(n434), .ZN(n645) );
  NOR2_X1 U389 ( .A1(KEYINPUT18), .A2(G953), .ZN(n404) );
  NOR2_X2 U390 ( .A1(n677), .A2(n367), .ZN(n431) );
  NAND2_X1 U391 ( .A1(n354), .A2(n544), .ZN(n367) );
  XNOR2_X1 U392 ( .A(n374), .B(KEYINPUT66), .ZN(n647) );
  NOR2_X1 U393 ( .A1(n771), .A2(n770), .ZN(n634) );
  NOR2_X1 U394 ( .A1(n693), .A2(n694), .ZN(n630) );
  XNOR2_X1 U395 ( .A(n545), .B(KEYINPUT33), .ZN(n705) );
  BUF_X1 U396 ( .A(n677), .Z(n420) );
  XNOR2_X1 U397 ( .A(n564), .B(n426), .ZN(n729) );
  XNOR2_X1 U398 ( .A(n602), .B(n603), .ZN(n624) );
  XNOR2_X1 U399 ( .A(n479), .B(n478), .ZN(n565) );
  AND2_X1 U400 ( .A1(n409), .A2(n408), .ZN(n407) );
  XNOR2_X1 U401 ( .A(G902), .B(KEYINPUT15), .ZN(n643) );
  XNOR2_X1 U402 ( .A(n525), .B(n524), .ZN(n569) );
  NAND2_X1 U403 ( .A1(n432), .A2(n635), .ZN(n391) );
  INV_X1 U404 ( .A(G134), .ZN(n480) );
  XNOR2_X1 U405 ( .A(n411), .B(KEYINPUT39), .ZN(n640) );
  NAND2_X1 U406 ( .A1(n627), .A2(n403), .ZN(n411) );
  AND2_X1 U407 ( .A1(n626), .A2(n435), .ZN(n627) );
  NOR2_X1 U408 ( .A1(n624), .A2(n625), .ZN(n403) );
  XNOR2_X1 U409 ( .A(n502), .B(n501), .ZN(n557) );
  XNOR2_X1 U410 ( .A(n492), .B(G478), .ZN(n604) );
  INV_X1 U411 ( .A(G224), .ZN(n405) );
  NAND2_X1 U412 ( .A1(KEYINPUT18), .A2(G953), .ZN(n408) );
  NOR2_X1 U413 ( .A1(n558), .A2(n720), .ZN(n377) );
  INV_X1 U414 ( .A(n643), .ZN(n375) );
  XNOR2_X1 U415 ( .A(G131), .B(G116), .ZN(n508) );
  XOR2_X1 U416 ( .A(KEYINPUT5), .B(G113), .Z(n509) );
  XOR2_X1 U417 ( .A(KEYINPUT3), .B(G119), .Z(n512) );
  XNOR2_X1 U418 ( .A(n424), .B(G122), .ZN(n466) );
  INV_X1 U419 ( .A(G113), .ZN(n424) );
  XNOR2_X1 U420 ( .A(n505), .B(n430), .ZN(n760) );
  XNOR2_X1 U421 ( .A(n391), .B(n390), .ZN(n641) );
  INV_X1 U422 ( .A(KEYINPUT48), .ZN(n390) );
  INV_X1 U423 ( .A(G237), .ZN(n446) );
  XNOR2_X1 U424 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U425 ( .A(n535), .B(KEYINPUT25), .ZN(n536) );
  XOR2_X1 U426 ( .A(G131), .B(G140), .Z(n519) );
  XNOR2_X1 U427 ( .A(n760), .B(G146), .ZN(n522) );
  INV_X1 U428 ( .A(KEYINPUT36), .ZN(n421) );
  NOR2_X1 U429 ( .A1(n358), .A2(n421), .ZN(n418) );
  XNOR2_X1 U430 ( .A(n462), .B(KEYINPUT0), .ZN(n463) );
  AND2_X1 U431 ( .A1(n557), .A2(n516), .ZN(n563) );
  XNOR2_X1 U432 ( .A(n488), .B(n487), .ZN(n491) );
  BUF_X1 U433 ( .A(n380), .Z(n740) );
  INV_X1 U434 ( .A(KEYINPUT89), .ZN(n376) );
  XNOR2_X1 U435 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n438) );
  NAND2_X1 U436 ( .A1(n407), .A2(n406), .ZN(n436) );
  INV_X1 U437 ( .A(G125), .ZN(n439) );
  XNOR2_X1 U438 ( .A(n466), .B(n465), .ZN(n470) );
  XNOR2_X1 U439 ( .A(G143), .B(KEYINPUT103), .ZN(n465) );
  XNOR2_X1 U440 ( .A(KEYINPUT105), .B(KEYINPUT11), .ZN(n467) );
  XOR2_X1 U441 ( .A(KEYINPUT104), .B(KEYINPUT106), .Z(n468) );
  XOR2_X1 U442 ( .A(G104), .B(KEYINPUT12), .Z(n472) );
  NAND2_X1 U443 ( .A1(n371), .A2(n370), .ZN(n374) );
  AND2_X1 U444 ( .A1(n372), .A2(n375), .ZN(n371) );
  NAND2_X1 U445 ( .A1(G234), .A2(G237), .ZN(n451) );
  XOR2_X1 U446 ( .A(KEYINPUT14), .B(KEYINPUT93), .Z(n452) );
  XNOR2_X1 U447 ( .A(n428), .B(n427), .ZN(n388) );
  INV_X1 U448 ( .A(KEYINPUT19), .ZN(n427) );
  INV_X1 U449 ( .A(n691), .ZN(n429) );
  INV_X1 U450 ( .A(G902), .ZN(n523) );
  XNOR2_X1 U451 ( .A(n601), .B(n515), .ZN(n614) );
  XNOR2_X1 U452 ( .A(n569), .B(KEYINPUT1), .ZN(n677) );
  XNOR2_X1 U453 ( .A(n415), .B(n414), .ZN(n413) );
  XNOR2_X1 U454 ( .A(n507), .B(n360), .ZN(n414) );
  XNOR2_X1 U455 ( .A(n510), .B(n513), .ZN(n415) );
  XNOR2_X1 U456 ( .A(n444), .B(n443), .ZN(n749) );
  XNOR2_X1 U457 ( .A(G128), .B(G119), .ZN(n526) );
  XNOR2_X1 U458 ( .A(n369), .B(n368), .ZN(n528) );
  XNOR2_X1 U459 ( .A(KEYINPUT97), .B(KEYINPUT23), .ZN(n369) );
  XNOR2_X1 U460 ( .A(G137), .B(KEYINPUT24), .ZN(n368) );
  XOR2_X1 U461 ( .A(G116), .B(G107), .Z(n486) );
  XOR2_X1 U462 ( .A(KEYINPUT9), .B(G122), .Z(n485) );
  XNOR2_X1 U463 ( .A(KEYINPUT109), .B(KEYINPUT107), .ZN(n482) );
  XOR2_X1 U464 ( .A(KEYINPUT108), .B(KEYINPUT7), .Z(n483) );
  AND2_X1 U465 ( .A1(n595), .A2(n594), .ZN(n631) );
  NOR2_X1 U466 ( .A1(n420), .A2(n354), .ZN(n540) );
  AND2_X1 U467 ( .A1(n601), .A2(n691), .ZN(n602) );
  XNOR2_X1 U468 ( .A(n522), .B(n357), .ZN(n664) );
  NOR2_X1 U469 ( .A1(n416), .A2(n356), .ZN(n733) );
  NAND2_X1 U470 ( .A1(n419), .A2(n417), .ZN(n416) );
  NOR2_X1 U471 ( .A1(n418), .A2(n420), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n568), .B(KEYINPUT31), .ZN(n730) );
  INV_X1 U473 ( .A(KEYINPUT111), .ZN(n426) );
  INV_X1 U474 ( .A(KEYINPUT110), .ZN(n425) );
  AND2_X1 U475 ( .A1(n422), .A2(n354), .ZN(n714) );
  XNOR2_X1 U476 ( .A(n423), .B(KEYINPUT87), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n739), .B(n738), .ZN(n393) );
  INV_X1 U478 ( .A(KEYINPUT60), .ZN(n394) );
  INV_X1 U479 ( .A(KEYINPUT56), .ZN(n396) );
  AND2_X1 U480 ( .A1(n410), .A2(n601), .ZN(n355) );
  NOR2_X1 U481 ( .A1(n616), .A2(n421), .ZN(n356) );
  XOR2_X1 U482 ( .A(n520), .B(n521), .Z(n357) );
  AND2_X1 U483 ( .A1(n450), .A2(n691), .ZN(n358) );
  XOR2_X1 U484 ( .A(G140), .B(G110), .Z(n359) );
  XNOR2_X1 U485 ( .A(KEYINPUT102), .B(KEYINPUT77), .ZN(n360) );
  AND2_X1 U486 ( .A1(n626), .A2(n684), .ZN(n361) );
  AND2_X1 U487 ( .A1(n358), .A2(n421), .ZN(n362) );
  XOR2_X1 U488 ( .A(n650), .B(n649), .Z(n363) );
  XOR2_X1 U489 ( .A(n656), .B(n659), .Z(n364) );
  XNOR2_X1 U490 ( .A(KEYINPUT62), .B(n653), .ZN(n365) );
  XOR2_X1 U491 ( .A(n655), .B(KEYINPUT91), .Z(n366) );
  AND2_X1 U492 ( .A1(n652), .A2(G953), .ZN(n743) );
  INV_X1 U493 ( .A(n743), .ZN(n401) );
  NOR2_X1 U494 ( .A1(n593), .A2(n367), .ZN(n626) );
  NAND2_X1 U495 ( .A1(n420), .A2(n367), .ZN(n679) );
  NOR2_X1 U496 ( .A1(n644), .A2(n669), .ZN(n642) );
  NAND2_X1 U497 ( .A1(n644), .A2(n373), .ZN(n370) );
  NAND2_X1 U498 ( .A1(n669), .A2(n373), .ZN(n372) );
  INV_X1 U499 ( .A(KEYINPUT2), .ZN(n373) );
  XNOR2_X1 U500 ( .A(n695), .B(KEYINPUT82), .ZN(n618) );
  INV_X1 U501 ( .A(n695), .ZN(n598) );
  XNOR2_X1 U502 ( .A(n377), .B(n376), .ZN(n559) );
  XNOR2_X1 U503 ( .A(n503), .B(n504), .ZN(n430) );
  XNOR2_X1 U504 ( .A(n542), .B(n541), .ZN(n378) );
  XNOR2_X1 U505 ( .A(n542), .B(n541), .ZN(n558) );
  XNOR2_X1 U506 ( .A(n431), .B(KEYINPUT76), .ZN(n410) );
  OR2_X1 U507 ( .A1(n378), .A2(n720), .ZN(n379) );
  BUF_X1 U508 ( .A(n669), .Z(n765) );
  NOR2_X1 U509 ( .A1(n733), .A2(n621), .ZN(n622) );
  XNOR2_X1 U510 ( .A(n742), .B(n741), .ZN(n389) );
  XNOR2_X1 U511 ( .A(n539), .B(n538), .ZN(n681) );
  BUF_X1 U512 ( .A(n569), .Z(n593) );
  NOR2_X1 U513 ( .A1(n647), .A2(n675), .ZN(n380) );
  XNOR2_X1 U514 ( .A(n553), .B(KEYINPUT35), .ZN(n381) );
  NOR2_X1 U515 ( .A1(n647), .A2(n675), .ZN(n662) );
  XNOR2_X1 U516 ( .A(n553), .B(KEYINPUT35), .ZN(n661) );
  XNOR2_X1 U517 ( .A(G143), .B(G128), .ZN(n481) );
  NOR2_X1 U518 ( .A1(n642), .A2(KEYINPUT2), .ZN(n383) );
  NAND2_X1 U519 ( .A1(n445), .A2(n749), .ZN(n386) );
  NAND2_X1 U520 ( .A1(n384), .A2(n385), .ZN(n387) );
  NAND2_X1 U521 ( .A1(n386), .A2(n387), .ZN(n656) );
  INV_X1 U522 ( .A(n445), .ZN(n384) );
  INV_X1 U523 ( .A(n749), .ZN(n385) );
  NAND2_X1 U524 ( .A1(n388), .A2(n461), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n631), .A2(n388), .ZN(n617) );
  NOR2_X1 U526 ( .A1(n712), .A2(G953), .ZN(n713) );
  XNOR2_X1 U527 ( .A(n638), .B(KEYINPUT38), .ZN(n435) );
  XNOR2_X2 U528 ( .A(n448), .B(n447), .ZN(n638) );
  NOR2_X1 U529 ( .A1(n389), .A2(n743), .ZN(G66) );
  NAND2_X1 U530 ( .A1(n410), .A2(n614), .ZN(n545) );
  XNOR2_X1 U531 ( .A(n567), .B(KEYINPUT96), .ZN(n392) );
  NAND2_X1 U532 ( .A1(n705), .A2(n392), .ZN(n548) );
  AND2_X1 U533 ( .A1(n392), .A2(n361), .ZN(n716) );
  NOR2_X1 U534 ( .A1(n393), .A2(n743), .ZN(G63) );
  XNOR2_X1 U535 ( .A(n395), .B(n394), .ZN(G60) );
  NAND2_X1 U536 ( .A1(n399), .A2(n401), .ZN(n395) );
  XNOR2_X1 U537 ( .A(n397), .B(n396), .ZN(G51) );
  NAND2_X1 U538 ( .A1(n400), .A2(n401), .ZN(n397) );
  XNOR2_X1 U539 ( .A(n398), .B(n366), .ZN(G57) );
  NAND2_X1 U540 ( .A1(n402), .A2(n401), .ZN(n398) );
  XNOR2_X1 U541 ( .A(n651), .B(n363), .ZN(n399) );
  XNOR2_X1 U542 ( .A(n660), .B(n364), .ZN(n400) );
  XNOR2_X1 U543 ( .A(n654), .B(n365), .ZN(n402) );
  NAND2_X1 U544 ( .A1(n404), .A2(G224), .ZN(n406) );
  XNOR2_X2 U545 ( .A(n585), .B(n584), .ZN(n644) );
  XNOR2_X2 U546 ( .A(n645), .B(KEYINPUT85), .ZN(n669) );
  NAND2_X1 U547 ( .A1(n405), .A2(KEYINPUT18), .ZN(n409) );
  XNOR2_X2 U548 ( .A(KEYINPUT71), .B(G101), .ZN(n511) );
  XNOR2_X2 U549 ( .A(G110), .B(G104), .ZN(n752) );
  INV_X1 U550 ( .A(n625), .ZN(n412) );
  XNOR2_X1 U551 ( .A(n522), .B(n413), .ZN(n653) );
  NAND2_X1 U552 ( .A1(n616), .A2(n362), .ZN(n419) );
  AND2_X1 U553 ( .A1(n616), .A2(n691), .ZN(n636) );
  NAND2_X1 U554 ( .A1(n563), .A2(n420), .ZN(n423) );
  INV_X1 U555 ( .A(n638), .ZN(n450) );
  NOR2_X1 U556 ( .A1(n730), .A2(n716), .ZN(n570) );
  AND2_X1 U557 ( .A1(n623), .A2(n622), .ZN(n432) );
  AND2_X1 U558 ( .A1(n614), .A2(n613), .ZN(n433) );
  AND2_X1 U559 ( .A1(n736), .A2(n735), .ZN(n434) );
  AND2_X1 U560 ( .A1(n726), .A2(n433), .ZN(n615) );
  XNOR2_X1 U561 ( .A(n533), .B(n476), .ZN(n759) );
  XNOR2_X1 U562 ( .A(n505), .B(n484), .ZN(n488) );
  XNOR2_X1 U563 ( .A(n436), .B(n481), .ZN(n437) );
  XNOR2_X1 U564 ( .A(n437), .B(n520), .ZN(n442) );
  XNOR2_X2 U565 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n504), .B(n438), .ZN(n440) );
  XNOR2_X1 U567 ( .A(n439), .B(G146), .ZN(n475) );
  XNOR2_X1 U568 ( .A(n440), .B(n475), .ZN(n441) );
  XNOR2_X1 U569 ( .A(n442), .B(n441), .ZN(n445) );
  XOR2_X1 U570 ( .A(KEYINPUT16), .B(n466), .Z(n444) );
  XNOR2_X1 U571 ( .A(n512), .B(n486), .ZN(n443) );
  NAND2_X1 U572 ( .A1(n656), .A2(n643), .ZN(n448) );
  NAND2_X1 U573 ( .A1(n523), .A2(n446), .ZN(n449) );
  NAND2_X1 U574 ( .A1(n449), .A2(G210), .ZN(n447) );
  NAND2_X1 U575 ( .A1(n449), .A2(G214), .ZN(n691) );
  XNOR2_X1 U576 ( .A(n452), .B(n451), .ZN(n457) );
  NAND2_X1 U577 ( .A1(G902), .A2(n457), .ZN(n453) );
  XNOR2_X1 U578 ( .A(KEYINPUT95), .B(n453), .ZN(n454) );
  NAND2_X1 U579 ( .A1(n454), .A2(G953), .ZN(n586) );
  INV_X1 U580 ( .A(n586), .ZN(n456) );
  INV_X1 U581 ( .A(G898), .ZN(n455) );
  NAND2_X1 U582 ( .A1(n456), .A2(n455), .ZN(n460) );
  NAND2_X1 U583 ( .A1(G952), .A2(n457), .ZN(n702) );
  NOR2_X1 U584 ( .A1(G953), .A2(n702), .ZN(n458) );
  XNOR2_X1 U585 ( .A(KEYINPUT94), .B(n458), .ZN(n588) );
  INV_X1 U586 ( .A(n588), .ZN(n459) );
  NAND2_X1 U587 ( .A1(n460), .A2(n459), .ZN(n461) );
  INV_X1 U588 ( .A(KEYINPUT70), .ZN(n462) );
  XNOR2_X2 U589 ( .A(n464), .B(n463), .ZN(n567) );
  XNOR2_X1 U590 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U591 ( .A(n470), .B(n469), .ZN(n474) );
  NOR2_X1 U592 ( .A1(G953), .A2(G237), .ZN(n506) );
  NAND2_X1 U593 ( .A1(G214), .A2(n506), .ZN(n471) );
  XNOR2_X1 U594 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U595 ( .A(n474), .B(n473), .ZN(n477) );
  XOR2_X1 U596 ( .A(n475), .B(KEYINPUT10), .Z(n533) );
  INV_X1 U597 ( .A(n519), .ZN(n476) );
  XNOR2_X1 U598 ( .A(n477), .B(n759), .ZN(n650) );
  NOR2_X1 U599 ( .A1(G902), .A2(n650), .ZN(n479) );
  XNOR2_X1 U600 ( .A(KEYINPUT13), .B(G475), .ZN(n478) );
  INV_X1 U601 ( .A(n565), .ZN(n493) );
  XNOR2_X1 U602 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U603 ( .A(n486), .B(n485), .ZN(n487) );
  NAND2_X1 U604 ( .A1(G234), .A2(n766), .ZN(n489) );
  XOR2_X1 U605 ( .A(KEYINPUT8), .B(n489), .Z(n529) );
  NAND2_X1 U606 ( .A1(G217), .A2(n529), .ZN(n490) );
  XNOR2_X1 U607 ( .A(n491), .B(n490), .ZN(n738) );
  NOR2_X1 U608 ( .A1(G902), .A2(n738), .ZN(n492) );
  NAND2_X1 U609 ( .A1(n493), .A2(n604), .ZN(n693) );
  XOR2_X1 U610 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n496) );
  NAND2_X1 U611 ( .A1(G234), .A2(n643), .ZN(n494) );
  XNOR2_X1 U612 ( .A(KEYINPUT20), .B(n494), .ZN(n534) );
  NAND2_X1 U613 ( .A1(n534), .A2(G221), .ZN(n495) );
  XNOR2_X1 U614 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U615 ( .A(KEYINPUT21), .B(n497), .ZN(n680) );
  INV_X1 U616 ( .A(KEYINPUT101), .ZN(n498) );
  XNOR2_X1 U617 ( .A(n680), .B(n498), .ZN(n543) );
  NOR2_X1 U618 ( .A1(n693), .A2(n543), .ZN(n499) );
  NAND2_X1 U619 ( .A1(n567), .A2(n499), .ZN(n502) );
  INV_X1 U620 ( .A(KEYINPUT68), .ZN(n500) );
  XNOR2_X1 U621 ( .A(n500), .B(KEYINPUT22), .ZN(n501) );
  XNOR2_X1 U622 ( .A(KEYINPUT73), .B(G137), .ZN(n503) );
  NAND2_X1 U623 ( .A1(n506), .A2(G210), .ZN(n507) );
  XNOR2_X1 U624 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U625 ( .A(n512), .B(n511), .ZN(n513) );
  NAND2_X1 U626 ( .A1(n653), .A2(n523), .ZN(n514) );
  INV_X1 U627 ( .A(KEYINPUT6), .ZN(n515) );
  INV_X1 U628 ( .A(n614), .ZN(n516) );
  NAND2_X1 U629 ( .A1(n766), .A2(G227), .ZN(n517) );
  XNOR2_X1 U630 ( .A(n517), .B(G107), .ZN(n518) );
  XNOR2_X1 U631 ( .A(n519), .B(n518), .ZN(n521) );
  NAND2_X1 U632 ( .A1(n664), .A2(n523), .ZN(n525) );
  INV_X1 U633 ( .A(G469), .ZN(n524) );
  XNOR2_X1 U634 ( .A(n359), .B(n526), .ZN(n527) );
  XNOR2_X1 U635 ( .A(n528), .B(n527), .ZN(n531) );
  NAND2_X1 U636 ( .A1(G221), .A2(n529), .ZN(n530) );
  XNOR2_X1 U637 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U638 ( .A(n532), .B(n533), .ZN(n741) );
  NOR2_X1 U639 ( .A1(n741), .A2(G902), .ZN(n539) );
  NAND2_X1 U640 ( .A1(G217), .A2(n534), .ZN(n537) );
  INV_X1 U641 ( .A(KEYINPUT98), .ZN(n535) );
  NAND2_X1 U642 ( .A1(n563), .A2(n540), .ZN(n542) );
  INV_X1 U643 ( .A(KEYINPUT32), .ZN(n541) );
  XOR2_X1 U644 ( .A(n558), .B(G119), .Z(G21) );
  INV_X1 U645 ( .A(n543), .ZN(n544) );
  INV_X1 U646 ( .A(KEYINPUT79), .ZN(n546) );
  XOR2_X1 U647 ( .A(n546), .B(KEYINPUT34), .Z(n547) );
  XNOR2_X1 U648 ( .A(n548), .B(n547), .ZN(n552) );
  INV_X1 U649 ( .A(n604), .ZN(n549) );
  NAND2_X1 U650 ( .A1(n549), .A2(n565), .ZN(n550) );
  XOR2_X1 U651 ( .A(n550), .B(KEYINPUT78), .Z(n551) );
  NAND2_X1 U652 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U653 ( .A(n554), .B(KEYINPUT72), .ZN(n560) );
  NOR2_X1 U654 ( .A1(n601), .A2(n354), .ZN(n555) );
  AND2_X1 U655 ( .A1(n420), .A2(n555), .ZN(n556) );
  AND2_X1 U656 ( .A1(n557), .A2(n556), .ZN(n720) );
  NAND2_X1 U657 ( .A1(n560), .A2(n559), .ZN(n562) );
  INV_X1 U658 ( .A(KEYINPUT75), .ZN(n561) );
  XNOR2_X1 U659 ( .A(n562), .B(n561), .ZN(n582) );
  NOR2_X1 U660 ( .A1(n565), .A2(n604), .ZN(n564) );
  NAND2_X1 U661 ( .A1(n604), .A2(n565), .ZN(n566) );
  INV_X1 U662 ( .A(n601), .ZN(n684) );
  NAND2_X1 U663 ( .A1(n355), .A2(n567), .ZN(n568) );
  NOR2_X1 U664 ( .A1(n618), .A2(n570), .ZN(n571) );
  XNOR2_X1 U665 ( .A(n571), .B(KEYINPUT112), .ZN(n572) );
  NOR2_X1 U666 ( .A1(n714), .A2(n572), .ZN(n574) );
  NAND2_X1 U667 ( .A1(n381), .A2(KEYINPUT44), .ZN(n573) );
  NAND2_X1 U668 ( .A1(n574), .A2(n573), .ZN(n576) );
  INV_X1 U669 ( .A(KEYINPUT88), .ZN(n575) );
  XNOR2_X1 U670 ( .A(n576), .B(n575), .ZN(n580) );
  NAND2_X1 U671 ( .A1(n379), .A2(KEYINPUT44), .ZN(n578) );
  INV_X1 U672 ( .A(KEYINPUT67), .ZN(n577) );
  XNOR2_X1 U673 ( .A(n578), .B(n577), .ZN(n579) );
  AND2_X1 U674 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U675 ( .A1(n582), .A2(n581), .ZN(n585) );
  INV_X1 U676 ( .A(KEYINPUT64), .ZN(n583) );
  XNOR2_X1 U677 ( .A(n583), .B(KEYINPUT45), .ZN(n584) );
  XOR2_X1 U678 ( .A(KEYINPUT113), .B(n586), .Z(n587) );
  NOR2_X1 U679 ( .A1(G900), .A2(n587), .ZN(n589) );
  NOR2_X1 U680 ( .A1(n589), .A2(n588), .ZN(n625) );
  NOR2_X1 U681 ( .A1(n625), .A2(n680), .ZN(n590) );
  AND2_X1 U682 ( .A1(n681), .A2(n590), .ZN(n591) );
  XNOR2_X1 U683 ( .A(KEYINPUT74), .B(n591), .ZN(n613) );
  AND2_X1 U684 ( .A1(n601), .A2(n613), .ZN(n592) );
  XNOR2_X1 U685 ( .A(KEYINPUT28), .B(n592), .ZN(n595) );
  INV_X1 U686 ( .A(n593), .ZN(n594) );
  INV_X1 U687 ( .A(n617), .ZN(n724) );
  OR2_X1 U688 ( .A1(KEYINPUT81), .A2(n598), .ZN(n596) );
  NAND2_X1 U689 ( .A1(n724), .A2(n596), .ZN(n597) );
  NAND2_X1 U690 ( .A1(n597), .A2(KEYINPUT47), .ZN(n600) );
  NAND2_X1 U691 ( .A1(n598), .A2(KEYINPUT81), .ZN(n599) );
  NAND2_X1 U692 ( .A1(n600), .A2(n599), .ZN(n612) );
  INV_X1 U693 ( .A(KEYINPUT30), .ZN(n603) );
  INV_X1 U694 ( .A(n624), .ZN(n610) );
  NAND2_X1 U695 ( .A1(n565), .A2(n412), .ZN(n605) );
  NOR2_X1 U696 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U697 ( .A1(n606), .A2(n450), .ZN(n608) );
  INV_X1 U698 ( .A(n626), .ZN(n607) );
  NOR2_X1 U699 ( .A1(n608), .A2(n607), .ZN(n609) );
  AND2_X1 U700 ( .A1(n610), .A2(n609), .ZN(n723) );
  XOR2_X1 U701 ( .A(KEYINPUT83), .B(n723), .Z(n611) );
  NOR2_X1 U702 ( .A1(n612), .A2(n611), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n615), .B(KEYINPUT114), .ZN(n616) );
  NOR2_X1 U704 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U705 ( .A1(KEYINPUT81), .A2(n619), .ZN(n620) );
  NOR2_X1 U706 ( .A1(KEYINPUT47), .A2(n620), .ZN(n621) );
  XNOR2_X1 U707 ( .A(n628), .B(KEYINPUT40), .ZN(n771) );
  NAND2_X1 U708 ( .A1(n435), .A2(n691), .ZN(n694) );
  XOR2_X1 U709 ( .A(KEYINPUT41), .B(KEYINPUT115), .Z(n629) );
  XNOR2_X1 U710 ( .A(n630), .B(n629), .ZN(n690) );
  INV_X1 U711 ( .A(n690), .ZN(n706) );
  AND2_X1 U712 ( .A1(n706), .A2(n631), .ZN(n632) );
  XNOR2_X1 U713 ( .A(KEYINPUT46), .B(KEYINPUT86), .ZN(n633) );
  XNOR2_X1 U714 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n420), .ZN(n637) );
  XNOR2_X1 U716 ( .A(n637), .B(KEYINPUT43), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n736) );
  NAND2_X1 U718 ( .A1(n640), .A2(n729), .ZN(n735) );
  NAND2_X1 U719 ( .A1(n645), .A2(KEYINPUT2), .ZN(n646) );
  NOR2_X1 U720 ( .A1(n644), .A2(n646), .ZN(n675) );
  NAND2_X1 U721 ( .A1(n662), .A2(G475), .ZN(n651) );
  XNOR2_X1 U722 ( .A(KEYINPUT69), .B(KEYINPUT122), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n648), .B(KEYINPUT59), .ZN(n649) );
  INV_X1 U724 ( .A(G952), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n380), .A2(G472), .ZN(n654) );
  XNOR2_X1 U726 ( .A(KEYINPUT116), .B(KEYINPUT63), .ZN(n655) );
  NAND2_X1 U727 ( .A1(n662), .A2(G210), .ZN(n660) );
  XOR2_X1 U728 ( .A(KEYINPUT90), .B(KEYINPUT80), .Z(n658) );
  XNOR2_X1 U729 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n657) );
  XOR2_X1 U730 ( .A(n658), .B(n657), .Z(n659) );
  XOR2_X1 U731 ( .A(n381), .B(G122), .Z(G24) );
  NAND2_X1 U732 ( .A1(n740), .A2(G469), .ZN(n666) );
  XNOR2_X1 U733 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n666), .B(n665), .ZN(n667) );
  NOR2_X1 U736 ( .A1(n667), .A2(n743), .ZN(G54) );
  INV_X1 U737 ( .A(KEYINPUT84), .ZN(n668) );
  NOR2_X1 U738 ( .A1(n383), .A2(n668), .ZN(n674) );
  INV_X1 U739 ( .A(n765), .ZN(n671) );
  NOR2_X1 U740 ( .A1(KEYINPUT2), .A2(KEYINPUT84), .ZN(n670) );
  NAND2_X1 U741 ( .A1(n671), .A2(n670), .ZN(n672) );
  INV_X1 U742 ( .A(n644), .ZN(n744) );
  NOR2_X1 U743 ( .A1(n672), .A2(n744), .ZN(n673) );
  NOR2_X1 U744 ( .A1(n674), .A2(n673), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n710) );
  XOR2_X1 U746 ( .A(KEYINPUT120), .B(KEYINPUT50), .Z(n678) );
  XNOR2_X1 U747 ( .A(n679), .B(n678), .ZN(n686) );
  NAND2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U749 ( .A(KEYINPUT49), .B(n682), .Z(n683) );
  NAND2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U752 ( .A1(n355), .A2(n687), .ZN(n688) );
  XOR2_X1 U753 ( .A(KEYINPUT51), .B(n688), .Z(n689) );
  NOR2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n700) );
  NOR2_X1 U755 ( .A1(n435), .A2(n691), .ZN(n692) );
  NOR2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n696) );
  OR2_X1 U758 ( .A1(n697), .A2(n696), .ZN(n698) );
  AND2_X1 U759 ( .A1(n705), .A2(n698), .ZN(n699) );
  OR2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U761 ( .A(n701), .B(KEYINPUT52), .ZN(n704) );
  INV_X1 U762 ( .A(n702), .ZN(n703) );
  NAND2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U764 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U765 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U766 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U767 ( .A(n711), .B(KEYINPUT121), .ZN(n712) );
  XNOR2_X1 U768 ( .A(n713), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U769 ( .A(G101), .B(n714), .Z(G3) );
  NAND2_X1 U770 ( .A1(n726), .A2(n716), .ZN(n715) );
  XNOR2_X1 U771 ( .A(n715), .B(G104), .ZN(G6) );
  XOR2_X1 U772 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n718) );
  NAND2_X1 U773 ( .A1(n716), .A2(n729), .ZN(n717) );
  XNOR2_X1 U774 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U775 ( .A(G107), .B(n719), .ZN(G9) );
  XOR2_X1 U776 ( .A(G110), .B(n720), .Z(G12) );
  XOR2_X1 U777 ( .A(G128), .B(KEYINPUT29), .Z(n722) );
  NAND2_X1 U778 ( .A1(n724), .A2(n729), .ZN(n721) );
  XNOR2_X1 U779 ( .A(n722), .B(n721), .ZN(G30) );
  XOR2_X1 U780 ( .A(G143), .B(n723), .Z(G45) );
  NAND2_X1 U781 ( .A1(n724), .A2(n726), .ZN(n725) );
  XNOR2_X1 U782 ( .A(n725), .B(G146), .ZN(G48) );
  XOR2_X1 U783 ( .A(G113), .B(KEYINPUT117), .Z(n728) );
  NAND2_X1 U784 ( .A1(n730), .A2(n726), .ZN(n727) );
  XNOR2_X1 U785 ( .A(n728), .B(n727), .ZN(G15) );
  NAND2_X1 U786 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U787 ( .A(n731), .B(KEYINPUT118), .ZN(n732) );
  XNOR2_X1 U788 ( .A(G116), .B(n732), .ZN(G18) );
  XNOR2_X1 U789 ( .A(n733), .B(G125), .ZN(n734) );
  XNOR2_X1 U790 ( .A(n734), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U791 ( .A(G134), .B(n735), .ZN(G36) );
  XOR2_X1 U792 ( .A(G140), .B(n736), .Z(n737) );
  XNOR2_X1 U793 ( .A(n737), .B(KEYINPUT119), .ZN(G42) );
  NAND2_X1 U794 ( .A1(n740), .A2(G478), .ZN(n739) );
  NAND2_X1 U795 ( .A1(n740), .A2(G217), .ZN(n742) );
  NAND2_X1 U796 ( .A1(n744), .A2(n766), .ZN(n748) );
  NAND2_X1 U797 ( .A1(G953), .A2(G224), .ZN(n745) );
  XNOR2_X1 U798 ( .A(KEYINPUT61), .B(n745), .ZN(n746) );
  NAND2_X1 U799 ( .A1(n746), .A2(G898), .ZN(n747) );
  NAND2_X1 U800 ( .A1(n748), .A2(n747), .ZN(n757) );
  XOR2_X1 U801 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n751) );
  XNOR2_X1 U802 ( .A(G101), .B(n749), .ZN(n750) );
  XNOR2_X1 U803 ( .A(n751), .B(n750), .ZN(n753) );
  XNOR2_X1 U804 ( .A(n753), .B(n752), .ZN(n755) );
  NOR2_X1 U805 ( .A1(G898), .A2(n766), .ZN(n754) );
  NOR2_X1 U806 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U807 ( .A(n757), .B(n756), .ZN(n758) );
  XOR2_X1 U808 ( .A(KEYINPUT123), .B(n758), .Z(G69) );
  XNOR2_X1 U809 ( .A(n760), .B(n759), .ZN(n764) );
  XNOR2_X1 U810 ( .A(n764), .B(G227), .ZN(n761) );
  NAND2_X1 U811 ( .A1(n761), .A2(G900), .ZN(n762) );
  NAND2_X1 U812 ( .A1(n762), .A2(G953), .ZN(n763) );
  XNOR2_X1 U813 ( .A(n763), .B(KEYINPUT126), .ZN(n769) );
  XNOR2_X1 U814 ( .A(n765), .B(n764), .ZN(n767) );
  NAND2_X1 U815 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U816 ( .A1(n769), .A2(n768), .ZN(G72) );
  XOR2_X1 U817 ( .A(G137), .B(n770), .Z(G39) );
  XNOR2_X1 U818 ( .A(G131), .B(KEYINPUT127), .ZN(n772) );
  XNOR2_X1 U819 ( .A(n772), .B(n771), .ZN(G33) );
endmodule

