//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1299, new_n1300, new_n1301, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(G20), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n212), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  OR2_X1    g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  AOI21_X1  g0048(.A(G1698), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G222), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G223), .A3(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n250), .B(new_n252), .C1(new_n253), .C2(new_n251), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n227), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(new_n227), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n206), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n262), .A2(new_n265), .A3(G274), .A4(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n262), .A2(G226), .A3(new_n263), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n258), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n269), .A2(G179), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n226), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n206), .A2(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G50), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n275), .A2(new_n277), .B1(G50), .B2(new_n274), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT69), .B1(G20), .B2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NOR3_X1   g0081(.A1(KEYINPUT69), .A2(G20), .A3(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n207), .A2(G33), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n283), .A2(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n207), .B1(new_n201), .B2(new_n202), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n288), .A2(KEYINPUT70), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(KEYINPUT70), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n287), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n279), .B1(new_n291), .B2(new_n273), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n269), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n270), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n269), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(G200), .B2(new_n269), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n292), .A2(KEYINPUT9), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n292), .A2(KEYINPUT9), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n299), .B(new_n304), .C1(new_n300), .C2(new_n301), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n296), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT18), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n262), .A2(G232), .A3(new_n263), .ZN(new_n308));
  INV_X1    g0108(.A(G33), .ZN(new_n309));
  INV_X1    g0109(.A(G87), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT75), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT75), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(G33), .A3(G87), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(G223), .A2(G1698), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n215), .B2(G1698), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n314), .B1(new_n251), .B2(new_n316), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n267), .B(new_n308), .C1(new_n317), .C2(new_n256), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G169), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n251), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n257), .B1(new_n321), .B2(new_n314), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n322), .A2(G179), .A3(new_n267), .A4(new_n308), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n247), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n248), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT74), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n330), .A2(KEYINPUT74), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n247), .A2(new_n207), .A3(new_n248), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT7), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n327), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G68), .ZN(new_n336));
  INV_X1    g0136(.A(G58), .ZN(new_n337));
  INV_X1    g0137(.A(G68), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(G20), .B1(new_n339), .B2(new_n202), .ZN(new_n340));
  INV_X1    g0140(.A(G159), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n283), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n336), .A2(KEYINPUT16), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n338), .B1(new_n334), .B2(new_n325), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(new_n342), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(new_n272), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n286), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n276), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n351), .A2(new_n275), .B1(new_n274), .B2(new_n350), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n307), .B(new_n324), .C1(new_n349), .C2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n342), .B1(new_n335), .B2(G68), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n273), .B1(new_n354), .B2(KEYINPUT16), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n352), .B1(new_n355), .B2(new_n347), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n319), .A2(new_n323), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT18), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n352), .ZN(new_n360));
  INV_X1    g0160(.A(G200), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n318), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n322), .A2(new_n297), .A3(new_n267), .A4(new_n308), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n348), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT17), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n348), .A2(new_n364), .A3(KEYINPUT17), .A4(new_n360), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n359), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n249), .A2(G232), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n251), .A2(G238), .A3(G1698), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n330), .A2(G107), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n257), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n262), .A2(G244), .A3(new_n263), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n267), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT71), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n375), .A2(new_n380), .A3(new_n377), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(G200), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n285), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(G20), .B2(G77), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n281), .A2(new_n282), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n350), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n273), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n276), .A2(G77), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n275), .A2(new_n389), .B1(G77), .B2(new_n274), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n382), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n297), .B1(new_n379), .B2(new_n381), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n379), .A2(new_n381), .ZN(new_n395));
  INV_X1    g0195(.A(G179), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n379), .A2(new_n293), .A3(new_n381), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n306), .A2(new_n370), .A3(new_n394), .A4(new_n399), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n274), .A2(G68), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n401), .B(KEYINPUT12), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n276), .A2(G68), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n283), .A2(new_n214), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n285), .A2(new_n253), .B1(new_n207), .B2(G68), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n272), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT11), .ZN(new_n407));
  OAI221_X1 g0207(.A(new_n402), .B1(new_n275), .B2(new_n403), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n406), .A2(new_n407), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n262), .A2(G238), .A3(new_n263), .ZN(new_n411));
  NOR2_X1   g0211(.A1(G226), .A2(G1698), .ZN(new_n412));
  INV_X1    g0212(.A(G232), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(G1698), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n251), .B1(G33), .B2(G97), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n411), .B(new_n267), .C1(new_n415), .C2(new_n256), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT13), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(G1698), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(G226), .B2(G1698), .ZN(new_n419));
  INV_X1    g0219(.A(G97), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n419), .A2(new_n330), .B1(new_n309), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n257), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT13), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(new_n411), .A4(new_n267), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n417), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G200), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n417), .A2(G190), .A3(new_n424), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n410), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n293), .B1(new_n417), .B2(new_n424), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT14), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n430), .A2(new_n431), .B1(new_n425), .B2(new_n396), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(KEYINPUT72), .A3(new_n431), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n425), .A2(new_n431), .A3(G169), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT72), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n410), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n429), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT73), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n441), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n400), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G1698), .ZN(new_n447));
  OAI211_X1 g0247(.A(G257), .B(new_n447), .C1(new_n328), .C2(new_n329), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT81), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n251), .A2(KEYINPUT81), .A3(G257), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n330), .A2(G303), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n251), .A2(G264), .A3(G1698), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n454), .A2(KEYINPUT82), .A3(new_n257), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT82), .B1(new_n454), .B2(new_n257), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n207), .C1(G33), .C2(new_n420), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n459), .B(new_n272), .C1(new_n207), .C2(G116), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT20), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n206), .A2(G33), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n274), .A2(new_n463), .A3(new_n226), .A4(new_n271), .ZN(new_n464));
  MUX2_X1   g0264(.A(new_n274), .B(new_n464), .S(G116), .Z(new_n465));
  AND2_X1   g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT5), .B(G41), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n262), .A2(G274), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n262), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n470), .B(G179), .C1(new_n217), .C2(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n457), .A2(new_n466), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n470), .B1(new_n475), .B2(new_n217), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n454), .A2(new_n257), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT82), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n454), .A2(KEYINPUT82), .A3(new_n257), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n462), .A2(new_n465), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G169), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT21), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n478), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n455), .B2(new_n456), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT21), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n293), .B1(new_n462), .B2(new_n465), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n477), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(KEYINPUT83), .B(new_n466), .C1(new_n483), .C2(new_n361), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n297), .B2(new_n488), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n466), .B1(new_n483), .B2(new_n361), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT83), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n492), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(G250), .B(new_n447), .C1(new_n328), .C2(new_n329), .ZN(new_n499));
  OAI211_X1 g0299(.A(G257), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n500));
  INV_X1    g0300(.A(G294), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n499), .B(new_n500), .C1(new_n309), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n257), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n262), .A2(new_n474), .A3(G264), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(new_n470), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n293), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n503), .A2(new_n504), .A3(new_n396), .A4(new_n470), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n207), .B(G87), .C1(new_n328), .C2(new_n329), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT22), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT22), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n251), .A2(new_n510), .A3(new_n207), .A4(G87), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G116), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G20), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT23), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n207), .B2(G107), .ZN(new_n516));
  INV_X1    g0316(.A(G107), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(KEYINPUT23), .A3(G20), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n514), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT24), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT24), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n512), .A2(new_n522), .A3(new_n519), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n273), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT25), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n274), .B2(G107), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n274), .A2(new_n525), .A3(G107), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n527), .A2(new_n528), .B1(new_n517), .B2(new_n464), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n506), .B(new_n507), .C1(new_n524), .C2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n523), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n522), .B1(new_n512), .B2(new_n519), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n272), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n529), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n505), .A2(G200), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n503), .A2(new_n504), .A3(G190), .A4(new_n470), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n530), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(G250), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n540));
  OAI211_X1 g0340(.A(G244), .B(new_n447), .C1(new_n328), .C2(new_n329), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n458), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT4), .B1(new_n249), .B2(G244), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n257), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n262), .A2(new_n474), .A3(G257), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n470), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G169), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n470), .A2(new_n546), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n541), .A2(new_n542), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n251), .A2(KEYINPUT4), .A3(G244), .A4(new_n447), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(new_n458), .A4(new_n540), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n550), .B1(new_n257), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G179), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n517), .A2(KEYINPUT76), .A3(KEYINPUT6), .A4(G97), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT76), .ZN(new_n558));
  NAND2_X1  g0358(.A1(KEYINPUT6), .A2(G97), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(G107), .ZN(new_n560));
  AND2_X1   g0360(.A1(G97), .A2(G107), .ZN(new_n561));
  NOR2_X1   g0361(.A1(G97), .A2(G107), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n557), .B(new_n560), .C1(new_n563), .C2(KEYINPUT6), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(G20), .B1(new_n386), .B2(G77), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n334), .A2(new_n325), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G107), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n272), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n464), .A2(G97), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n274), .A2(new_n420), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n570), .A2(KEYINPUT77), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT77), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n556), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n361), .B1(new_n545), .B2(new_n547), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n577), .A2(KEYINPUT79), .B1(new_n548), .B2(new_n297), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n569), .A2(KEYINPUT78), .A3(new_n574), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT78), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n273), .B1(new_n565), .B2(new_n567), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n572), .A2(new_n573), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT79), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n554), .A2(new_n584), .A3(G190), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n578), .A2(new_n579), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(G238), .B(new_n447), .C1(new_n328), .C2(new_n329), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n587), .A2(new_n513), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n251), .A2(G244), .A3(G1698), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n256), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(G250), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n468), .B2(KEYINPUT80), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n592), .B(new_n262), .C1(KEYINPUT80), .C2(new_n468), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n262), .A2(G274), .A3(new_n468), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n293), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n589), .A2(new_n513), .A3(new_n587), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n257), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n598), .A2(new_n396), .A3(new_n594), .A4(new_n593), .ZN(new_n599));
  NAND3_X1  g0399(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n207), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n562), .A2(new_n310), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n207), .B(G68), .C1(new_n328), .C2(new_n329), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n285), .B2(new_n420), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n272), .ZN(new_n608));
  INV_X1    g0408(.A(new_n383), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n609), .A2(new_n274), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n608), .B(new_n610), .C1(new_n464), .C2(new_n383), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n596), .A2(new_n599), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n590), .B2(new_n595), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n598), .A2(G190), .A3(new_n594), .A4(new_n593), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n464), .A2(new_n310), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n608), .A2(new_n610), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n539), .A2(new_n576), .A3(new_n586), .A4(new_n618), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n446), .A2(new_n498), .A3(new_n619), .ZN(G372));
  INV_X1    g0420(.A(new_n399), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n621), .A2(new_n428), .B1(new_n438), .B2(new_n439), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n358), .B(new_n353), .C1(new_n622), .C2(new_n369), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n303), .A2(new_n305), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n296), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n586), .A2(new_n576), .A3(new_n618), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n481), .A2(new_n482), .ZN(new_n627));
  INV_X1    g0427(.A(new_n476), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n484), .A3(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n489), .B1(new_n488), .B2(new_n490), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n629), .B(new_n530), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n626), .A2(new_n537), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n612), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n556), .A2(new_n575), .A3(new_n612), .A4(new_n617), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(KEYINPUT26), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n579), .A2(new_n583), .B1(new_n549), .B2(new_n555), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n618), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n625), .B1(new_n446), .B2(new_n642), .ZN(G369));
  NAND3_X1  g0443(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n466), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n492), .B(new_n652), .C1(new_n494), .C2(new_n497), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n651), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n506), .A2(new_n507), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n533), .B2(new_n534), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n649), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n649), .B1(new_n524), .B2(new_n529), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n530), .A2(new_n537), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n656), .A2(G330), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n649), .B(KEYINPUT85), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n530), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT84), .B1(new_n492), .B2(new_n649), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT84), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n654), .A2(new_n668), .A3(new_n650), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n666), .B1(new_n670), .B2(new_n663), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n664), .A2(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n210), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n602), .A2(G116), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G1), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n225), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(new_n675), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  INV_X1    g0480(.A(new_n665), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n641), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT29), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n612), .B(KEYINPUT89), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n635), .A2(KEYINPUT90), .A3(new_n638), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n637), .A2(KEYINPUT26), .A3(new_n618), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT90), .B1(new_n635), .B2(new_n638), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n586), .A2(new_n537), .A3(new_n576), .A4(new_n618), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n492), .B2(new_n530), .ZN(new_n692));
  OAI211_X1 g0492(.A(KEYINPUT29), .B(new_n650), .C1(new_n690), .C2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT31), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n590), .A2(new_n595), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n503), .A2(new_n504), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n697), .A3(new_n554), .A4(new_n628), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n695), .B1(new_n698), .B2(new_n457), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n598), .A2(new_n594), .A3(new_n593), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n503), .A2(new_n504), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n700), .A2(new_n701), .A3(new_n476), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(KEYINPUT30), .A3(new_n627), .A4(new_n554), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n488), .A2(KEYINPUT87), .A3(new_n396), .A4(new_n700), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n548), .A2(KEYINPUT88), .A3(new_n505), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT88), .B1(new_n548), .B2(new_n505), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT87), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n700), .A2(new_n396), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n483), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n704), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n694), .B1(new_n713), .B2(new_n650), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n586), .A2(new_n576), .A3(new_n618), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n538), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n495), .A2(new_n496), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n717), .B(new_n493), .C1(new_n297), .C2(new_n488), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n716), .A2(new_n718), .A3(new_n492), .A4(new_n681), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n699), .A2(new_n703), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n712), .A2(new_n705), .A3(new_n708), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g0522(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n722), .A2(new_n665), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n714), .A2(new_n719), .A3(new_n725), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n684), .A2(new_n693), .B1(G330), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n680), .B1(new_n727), .B2(G1), .ZN(G364));
  NOR2_X1   g0528(.A1(new_n656), .A2(G330), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n656), .A2(G330), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n207), .A2(G13), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n206), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n674), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n730), .A2(new_n731), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n226), .B1(G20), .B2(new_n293), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n207), .A2(G179), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n310), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G190), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G159), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(KEYINPUT32), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n207), .A2(new_n396), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(new_n297), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n742), .B(new_n747), .C1(G68), .C2(new_n750), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n748), .A2(new_n743), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n251), .B1(new_n753), .B2(new_n253), .ZN(new_n754));
  NOR4_X1   g0554(.A1(new_n207), .A2(new_n396), .A3(new_n297), .A4(G200), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n754), .B1(G58), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n740), .A2(new_n297), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n746), .A2(KEYINPUT32), .B1(G107), .B2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n297), .A2(G179), .A3(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n207), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n748), .A2(G190), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G97), .A2(new_n762), .B1(new_n764), .B2(G50), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n751), .A2(new_n756), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G329), .A2(new_n745), .B1(new_n755), .B2(G322), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n251), .B1(new_n752), .B2(G311), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n764), .A2(G326), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT33), .B(G317), .ZN(new_n771));
  INV_X1    g0571(.A(new_n741), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n750), .A2(new_n771), .B1(new_n772), .B2(G303), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n762), .A2(G294), .B1(new_n758), .B2(G283), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n769), .A2(new_n770), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n739), .B1(new_n766), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n738), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT92), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n673), .A2(new_n251), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n225), .A2(new_n467), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n782), .B(new_n783), .C1(new_n245), .C2(new_n467), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n673), .A2(new_n330), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n785), .A2(G355), .B1(new_n216), .B2(new_n673), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n781), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n776), .A2(new_n736), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n779), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n788), .B1(new_n656), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n737), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  INV_X1    g0592(.A(new_n398), .ZN(new_n793));
  AOI21_X1  g0593(.A(G179), .B1(new_n379), .B2(new_n381), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n793), .A2(new_n794), .A3(new_n391), .A4(new_n649), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n649), .B1(new_n388), .B2(new_n390), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n392), .B2(new_n393), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n795), .B1(new_n399), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT94), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n682), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT95), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n636), .A2(new_n639), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n681), .B(new_n798), .C1(new_n692), .C2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n726), .A2(G330), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n800), .A2(new_n801), .A3(new_n805), .A4(new_n803), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n800), .A2(new_n803), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(KEYINPUT95), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n735), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n798), .A2(new_n778), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G116), .A2(new_n752), .B1(new_n755), .B2(G294), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n814), .B(new_n330), .C1(new_n815), .C2(new_n744), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G303), .A2(new_n764), .B1(new_n758), .B2(G87), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n517), .B2(new_n741), .ZN(new_n818));
  INV_X1    g0618(.A(G283), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n761), .A2(new_n420), .B1(new_n749), .B2(new_n819), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n816), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n251), .B1(new_n744), .B2(new_n822), .C1(new_n214), .C2(new_n741), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n761), .A2(new_n337), .B1(new_n757), .B2(new_n338), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G159), .A2(new_n752), .B1(new_n755), .B2(G143), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G137), .A2(new_n764), .B1(new_n750), .B2(G150), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT93), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n826), .A2(KEYINPUT93), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n825), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT34), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n823), .B(new_n824), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n821), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n738), .A2(new_n777), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n835), .A2(new_n739), .B1(G77), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n735), .B1(new_n813), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT96), .B1(new_n812), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT96), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n807), .A2(new_n808), .B1(KEYINPUT95), .B2(new_n810), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n842), .B(new_n839), .C1(new_n843), .C2(new_n735), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n841), .A2(new_n844), .ZN(G384));
  NOR2_X1   g0645(.A1(new_n732), .A2(new_n206), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n344), .A2(new_n272), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n354), .A2(KEYINPUT16), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n360), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n647), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n359), .B2(new_n369), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n349), .A2(new_n352), .B1(new_n324), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n365), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n849), .B1(new_n324), .B2(new_n850), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n356), .B2(new_n364), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n854), .A2(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n852), .A2(new_n858), .A3(KEYINPUT38), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n356), .A2(new_n647), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT99), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n367), .A2(new_n861), .A3(new_n368), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(new_n358), .A3(new_n353), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n861), .B1(new_n367), .B2(new_n368), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n357), .A2(new_n647), .B1(new_n348), .B2(new_n360), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n866), .B2(KEYINPUT98), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n854), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n853), .A2(KEYINPUT98), .A3(KEYINPUT37), .A4(new_n365), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n859), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n797), .A2(new_n399), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n397), .A2(new_n398), .A3(new_n650), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n439), .A2(new_n649), .ZN(new_n877));
  INV_X1    g0677(.A(new_n434), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT72), .B1(new_n430), .B2(new_n431), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n878), .A2(new_n432), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n428), .B(new_n877), .C1(new_n880), .C2(new_n410), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n439), .B(new_n649), .C1(new_n438), .C2(new_n429), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n876), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n650), .B1(new_n720), .B2(new_n721), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n884), .B1(new_n885), .B2(new_n724), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n498), .A2(new_n619), .A3(new_n665), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT40), .B1(new_n873), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n852), .A2(new_n858), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n872), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n852), .A2(new_n858), .A3(KEYINPUT38), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT40), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n719), .B(new_n884), .C1(new_n885), .C2(new_n724), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n894), .A3(new_n883), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n445), .A2(new_n894), .ZN(new_n897));
  OAI21_X1  g0697(.A(G330), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n898), .A2(KEYINPUT100), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n897), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(KEYINPUT100), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n438), .A2(new_n439), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n903), .A2(new_n649), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n904), .B(new_n905), .C1(new_n873), .C2(KEYINPUT39), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n881), .A2(new_n882), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n803), .B2(new_n875), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n891), .A2(new_n892), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n908), .A2(new_n909), .B1(new_n359), .B2(new_n647), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n445), .A2(new_n684), .A3(new_n693), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n625), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n911), .B(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n846), .B1(new_n902), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n914), .B2(new_n902), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n678), .A2(new_n253), .A3(new_n339), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(G68), .B2(new_n201), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n918), .A2(new_n206), .A3(G13), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT97), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT36), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n227), .A2(G20), .A3(G116), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n564), .B2(KEYINPUT35), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(KEYINPUT35), .B2(new_n564), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n920), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n921), .B2(new_n924), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n916), .A2(new_n926), .ZN(G367));
  INV_X1    g0727(.A(KEYINPUT43), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n579), .A2(new_n583), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n586), .B(new_n576), .C1(new_n929), .C2(new_n681), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n637), .A2(new_n665), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n658), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n665), .B1(new_n933), .B2(new_n576), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n492), .A2(KEYINPUT84), .A3(new_n649), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n668), .B1(new_n654), .B2(new_n650), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n663), .B(new_n932), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT42), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n662), .B1(new_n667), .B2(new_n669), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(KEYINPUT42), .A3(new_n932), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n934), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n928), .B1(new_n942), .B2(KEYINPUT102), .ZN(new_n943));
  INV_X1    g0743(.A(new_n934), .ZN(new_n944));
  AND4_X1   g0744(.A1(KEYINPUT42), .A2(new_n670), .A3(new_n663), .A4(new_n932), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT42), .B1(new_n940), .B2(new_n932), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT102), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT43), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n616), .A2(new_n650), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n618), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n951), .A2(KEYINPUT101), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n950), .A2(new_n612), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(KEYINPUT101), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n942), .A2(new_n956), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n943), .A2(new_n949), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n955), .B1(new_n943), .B2(new_n949), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT103), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n932), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n664), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n942), .A2(KEYINPUT102), .A3(new_n928), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT43), .B1(new_n947), .B2(new_n948), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n956), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT103), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n943), .A2(new_n949), .A3(new_n957), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n960), .A2(new_n963), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n963), .B1(new_n960), .B2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n670), .A2(new_n663), .ZN(new_n972));
  INV_X1    g0772(.A(new_n666), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT44), .B1(new_n974), .B2(new_n961), .ZN(new_n975));
  OAI211_X1 g0775(.A(KEYINPUT44), .B(new_n961), .C1(new_n940), .C2(new_n666), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT45), .B1(new_n671), .B2(new_n932), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT45), .ZN(new_n979));
  NOR4_X1   g0779(.A1(new_n940), .A2(new_n961), .A3(new_n979), .A4(new_n666), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n975), .A2(new_n977), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(G330), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n982), .B(new_n662), .C1(new_n653), .C2(new_n655), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n670), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n663), .B1(new_n656), .B2(G330), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n985), .B1(new_n986), .B2(new_n983), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n731), .A2(new_n662), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n988), .A2(new_n664), .A3(new_n670), .ZN(new_n989));
  AND3_X1   g0789(.A1(new_n727), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n979), .B1(new_n974), .B2(new_n961), .ZN(new_n991));
  INV_X1    g0791(.A(new_n980), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT44), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n671), .B2(new_n932), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n976), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n664), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n984), .A2(new_n990), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n727), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n674), .B(KEYINPUT41), .Z(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n734), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n970), .A2(new_n971), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n956), .A2(new_n779), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n781), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n210), .B2(new_n383), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n782), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(new_n238), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n735), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n772), .A2(G116), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT46), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n251), .B1(new_n755), .B2(G303), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G283), .A2(new_n752), .B1(new_n745), .B2(G317), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n761), .A2(new_n517), .B1(new_n749), .B2(new_n501), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n763), .A2(new_n815), .B1(new_n757), .B2(new_n420), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT104), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n758), .A2(G77), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n337), .B2(new_n741), .C1(new_n341), .C2(new_n749), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G68), .A2(new_n762), .B1(new_n764), .B2(G143), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n201), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n330), .B1(new_n1022), .B2(new_n752), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G137), .A2(new_n745), .B1(new_n755), .B2(G150), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1018), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT47), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1009), .B1(new_n1027), .B2(new_n738), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1004), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(KEYINPUT105), .B1(new_n1003), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n960), .A2(new_n969), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n962), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n999), .A2(new_n1001), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n733), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n960), .A2(new_n969), .A3(new_n963), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT105), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n1029), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1031), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(G387));
  INV_X1    g0841(.A(new_n990), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n727), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n989), .A2(new_n987), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1043), .A2(new_n1044), .A3(KEYINPUT109), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n674), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT109), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1044), .A2(new_n733), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G303), .A2(new_n752), .B1(new_n755), .B2(G317), .ZN(new_n1050));
  XOR2_X1   g0850(.A(KEYINPUT107), .B(G322), .Z(new_n1051));
  OAI221_X1 g0851(.A(new_n1050), .B1(new_n815), .B2(new_n749), .C1(new_n763), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT48), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n762), .A2(G283), .B1(new_n772), .B2(G294), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT49), .Z(new_n1058));
  AOI21_X1  g0858(.A(new_n251), .B1(new_n745), .B2(G326), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n216), .B2(new_n757), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n762), .A2(new_n609), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n253), .B2(new_n741), .C1(new_n286), .C2(new_n749), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n755), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n251), .B1(new_n1064), .B2(new_n214), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n753), .A2(new_n338), .B1(new_n744), .B2(new_n284), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n763), .A2(new_n341), .B1(new_n757), .B2(new_n420), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n738), .B1(new_n1061), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n785), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n1070), .A2(new_n676), .B1(G107), .B2(new_n210), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n350), .A2(new_n214), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT50), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n676), .B(new_n467), .C1(new_n338), .C2(new_n253), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n782), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n235), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(KEYINPUT106), .A2(new_n1076), .B1(new_n1077), .B2(G45), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1076), .A2(KEYINPUT106), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1071), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1069), .B(new_n735), .C1(new_n781), .C2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT108), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n662), .B2(new_n779), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1049), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1048), .A2(new_n1086), .ZN(G393));
  INV_X1    g0887(.A(new_n997), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n664), .B1(new_n993), .B2(new_n996), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n961), .A2(new_n779), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1005), .B1(new_n420), .B2(new_n210), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1007), .A2(new_n242), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n735), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1064), .A2(new_n341), .B1(new_n284), .B2(new_n763), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT51), .Z(new_n1096));
  AOI21_X1  g0896(.A(new_n330), .B1(new_n745), .B2(G143), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n286), .B2(new_n753), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n749), .A2(new_n201), .B1(new_n757), .B2(new_n310), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n761), .A2(new_n253), .B1(new_n741), .B2(new_n338), .ZN(new_n1100));
  OR4_X1    g0900(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT110), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n761), .A2(new_n216), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n330), .B1(new_n517), .B2(new_n757), .C1(new_n753), .C2(new_n501), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1104), .B(new_n1105), .C1(G303), .C2(new_n750), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n764), .A2(G317), .B1(new_n755), .B2(G311), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT52), .Z(new_n1108));
  OAI22_X1  g0908(.A1(new_n744), .A2(new_n1051), .B1(new_n741), .B2(new_n819), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1110), .A2(KEYINPUT111), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(KEYINPUT111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1106), .A2(new_n1108), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1103), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1094), .B1(new_n1115), .B2(new_n738), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1090), .A2(new_n734), .B1(new_n1091), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1042), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n674), .A3(new_n998), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(G390));
  OAI21_X1  g0920(.A(new_n905), .B1(new_n873), .B2(KEYINPUT39), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT112), .B1(new_n908), .B2(new_n904), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT112), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n904), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n665), .B1(new_n633), .B2(new_n640), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n795), .B1(new_n1125), .B2(new_n874), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1123), .B(new_n1124), .C1(new_n1126), .C2(new_n907), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1121), .A2(new_n1122), .A3(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n650), .B(new_n874), .C1(new_n690), .C2(new_n692), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n907), .B1(new_n1129), .B2(new_n875), .ZN(new_n1130));
  OR3_X1    g0930(.A1(new_n1130), .A2(new_n873), .A3(new_n904), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(G330), .B(new_n883), .C1(new_n886), .C2(new_n887), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT113), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n894), .A2(KEYINPUT113), .A3(G330), .A4(new_n883), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1132), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n665), .A2(new_n724), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n885), .A2(KEYINPUT31), .B1(new_n713), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(G330), .B(new_n798), .C1(new_n887), .C2(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1141), .A2(new_n907), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1128), .A2(new_n1142), .A3(new_n1131), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1138), .A2(new_n734), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(KEYINPUT115), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT115), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1138), .A2(new_n1146), .A3(new_n734), .A4(new_n1143), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n735), .B1(new_n350), .B2(new_n837), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT116), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n764), .A2(G283), .B1(new_n752), .B2(G97), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n517), .B2(new_n749), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT117), .Z(new_n1153));
  OAI22_X1  g0953(.A1(new_n338), .A2(new_n757), .B1(new_n741), .B2(new_n310), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n330), .B1(new_n744), .B2(new_n501), .C1(new_n1064), .C2(new_n216), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(G77), .C2(new_n762), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n741), .A2(new_n284), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT53), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n330), .B1(new_n745), .B2(G125), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G159), .A2(new_n762), .B1(new_n764), .B2(G128), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G137), .A2(new_n750), .B1(new_n1022), .B2(new_n758), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT54), .B(G143), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n752), .A2(new_n1163), .B1(new_n755), .B2(G132), .ZN(new_n1164));
  AND4_X1   g0964(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1153), .A2(new_n1156), .B1(new_n1158), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1150), .B1(new_n1166), .B2(new_n739), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1121), .B2(new_n777), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1148), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n400), .A2(new_n442), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1171), .A2(G330), .A3(new_n443), .A4(new_n894), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n912), .A2(new_n625), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1141), .A2(new_n907), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1135), .A2(new_n1174), .A3(new_n1136), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1126), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1129), .A2(new_n875), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n876), .B(KEYINPUT94), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n894), .A3(G330), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1178), .B1(new_n1180), .B2(new_n907), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n1142), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1173), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1138), .A2(new_n1183), .A3(new_n1143), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n674), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT114), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1128), .A2(new_n1142), .A3(new_n1131), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1128), .A2(new_n1131), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1186), .B1(new_n1189), .B2(new_n1183), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1177), .A2(new_n1182), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1173), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1193), .B(KEYINPUT114), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1185), .B1(new_n1190), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1170), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(G378));
  INV_X1    g0997(.A(KEYINPUT120), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n911), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(KEYINPUT121), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT121), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n911), .A2(new_n1198), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n624), .A2(new_n295), .ZN(new_n1203));
  XOR2_X1   g1003(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n292), .A2(new_n850), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT119), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1204), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n306), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1205), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1207), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n306), .A2(new_n1208), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n296), .B(new_n1204), .C1(new_n303), .C2(new_n305), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n896), .A2(G330), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(KEYINPUT38), .B1(new_n865), .B2(new_n870), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n894), .B(new_n883), .C1(new_n1218), .C2(new_n859), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n888), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1219), .A2(KEYINPUT40), .B1(new_n1220), .B2(new_n893), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1215), .B1(new_n1221), .B2(new_n982), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1200), .A2(new_n1202), .A3(new_n1217), .A4(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1201), .B1(new_n911), .B2(new_n1198), .ZN(new_n1224));
  AOI211_X1 g1024(.A(KEYINPUT120), .B(KEYINPUT121), .C1(new_n906), .C2(new_n910), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1216), .B1(new_n896), .B2(G330), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n982), .B(new_n1215), .C1(new_n889), .C2(new_n895), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n1224), .A2(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1223), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1216), .A2(new_n777), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n763), .A2(new_n216), .B1(new_n757), .B2(new_n337), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G97), .B2(new_n750), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n251), .A2(G41), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G283), .B2(new_n745), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n609), .A2(new_n752), .B1(new_n755), .B2(G107), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n762), .A2(G68), .B1(new_n772), .B2(G77), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1232), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT58), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1233), .B(new_n214), .C1(G33), .C2(G41), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(G125), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1242), .A2(new_n763), .B1(new_n749), .B2(new_n822), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G137), .A2(new_n752), .B1(new_n755), .B2(G128), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n741), .B2(new_n1162), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1243), .B(new_n1245), .C1(G150), .C2(new_n762), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n758), .A2(G159), .ZN(new_n1249));
  AOI211_X1 g1049(.A(G33), .B(G41), .C1(new_n745), .C2(G124), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1241), .B1(new_n1238), .B2(new_n1237), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n738), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT118), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n736), .B(new_n1255), .C1(new_n201), .C2(new_n836), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1229), .A2(new_n734), .B1(new_n1230), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1173), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n911), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1222), .A2(new_n1217), .A3(new_n906), .A4(new_n910), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1260), .A3(KEYINPUT57), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n674), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1184), .A2(new_n1192), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT57), .B1(new_n1229), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1257), .B1(new_n1262), .B2(new_n1264), .ZN(G375));
  NAND2_X1  g1065(.A1(new_n907), .A2(new_n777), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n517), .A2(new_n753), .B1(new_n1064), .B2(new_n819), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n251), .B(new_n1267), .C1(G303), .C2(new_n745), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n216), .A2(new_n749), .B1(new_n763), .B2(new_n501), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(G97), .B2(new_n772), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1268), .A2(new_n1019), .A3(new_n1062), .A4(new_n1270), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n761), .A2(new_n214), .B1(new_n741), .B2(new_n341), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G132), .B2(new_n764), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n330), .B1(new_n745), .B2(G128), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(G150), .A2(new_n752), .B1(new_n755), .B2(G137), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n750), .A2(new_n1163), .B1(new_n758), .B2(G58), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n739), .B1(new_n1271), .B2(new_n1277), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n736), .B(new_n1278), .C1(new_n338), .C2(new_n836), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1266), .A2(new_n1279), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1175), .A2(new_n1176), .B1(new_n1181), .B2(new_n1142), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1281), .B2(new_n733), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT122), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(KEYINPUT122), .B(new_n1280), .C1(new_n1281), .C2(new_n733), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1281), .A2(new_n1173), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1193), .A2(new_n1001), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(G381));
  INV_X1    g1089(.A(G390), .ZN(new_n1290));
  INV_X1    g1090(.A(G384), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1086), .B(new_n791), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(G378), .A2(G381), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1296));
  OR2_X1    g1096(.A1(G375), .A2(KEYINPUT123), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1295), .A2(new_n1040), .A3(new_n1296), .A4(new_n1297), .ZN(G407));
  NAND2_X1  g1098(.A1(new_n648), .A2(G213), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(G378), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(new_n1297), .A3(new_n1296), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(G407), .A2(G213), .A3(new_n1301), .ZN(G409));
  AOI21_X1  g1102(.A(new_n675), .B1(new_n1189), .B2(new_n1183), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1194), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT114), .B1(new_n1305), .B2(new_n1193), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1303), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1168), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1229), .A2(new_n1001), .A3(new_n1263), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1259), .A2(new_n1260), .A3(new_n734), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1256), .A2(new_n1230), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1307), .B(new_n1308), .C1(new_n1309), .C2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(G375), .B2(new_n1196), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1299), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT124), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(G384), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n841), .A2(KEYINPUT124), .A3(new_n844), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1286), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1281), .A2(KEYINPUT60), .A3(new_n1173), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n674), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1193), .A2(KEYINPUT60), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1321), .B1(new_n1287), .B2(new_n1322), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1317), .B(new_n1318), .C1(new_n1319), .C2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1287), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(new_n674), .A3(new_n1320), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1326), .A2(KEYINPUT124), .A3(new_n1291), .A4(new_n1286), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n648), .A2(G213), .A3(G2897), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1324), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1324), .B2(new_n1327), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT61), .B1(new_n1315), .B2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1314), .A2(new_n1299), .A3(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n791), .B1(new_n1048), .B2(new_n1086), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1336), .A2(new_n1293), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1003), .A2(new_n1030), .A3(new_n1290), .ZN(new_n1338));
  AOI21_X1  g1138(.A(G390), .B1(new_n1037), .B2(new_n1029), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1337), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  XNOR2_X1  g1140(.A(G390), .B(KEYINPUT125), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1031), .A2(new_n1039), .A3(new_n1341), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n971), .A2(new_n1002), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1030), .B1(new_n1343), .B2(new_n1036), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1337), .B1(new_n1344), .B2(G390), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1346));
  AOI22_X1  g1146(.A1(new_n1334), .A2(new_n1335), .B1(new_n1340), .B2(new_n1346), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1314), .A2(KEYINPUT63), .A3(new_n1299), .A4(new_n1333), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT126), .ZN(new_n1349));
  AND2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1351));
  OAI211_X1 g1151(.A(new_n1332), .B(new_n1347), .C1(new_n1350), .C2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1334), .A2(KEYINPUT62), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1315), .A2(new_n1331), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT61), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT62), .ZN(new_n1356));
  NAND4_X1  g1156(.A1(new_n1314), .A2(new_n1356), .A3(new_n1299), .A4(new_n1333), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1353), .A2(new_n1354), .A3(new_n1355), .A4(new_n1357), .ZN(new_n1358));
  AND3_X1   g1158(.A1(new_n1346), .A2(KEYINPUT127), .A3(new_n1340), .ZN(new_n1359));
  AOI21_X1  g1159(.A(KEYINPUT127), .B1(new_n1346), .B2(new_n1340), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1358), .A2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1352), .A2(new_n1362), .ZN(G405));
  NAND2_X1  g1163(.A1(new_n1346), .A2(new_n1340), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1364), .A2(new_n1327), .A3(new_n1324), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1346), .A2(new_n1333), .A3(new_n1340), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  XNOR2_X1  g1167(.A(G378), .B(G375), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1367), .A2(new_n1369), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1365), .A2(new_n1368), .A3(new_n1366), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1370), .A2(new_n1371), .ZN(G402));
endmodule


