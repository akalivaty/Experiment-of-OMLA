//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(G155gat), .B(G162gat), .Z(new_n204));
  XNOR2_X1  g003(.A(G141gat), .B(G148gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT80), .B(KEYINPUT3), .Z(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G141gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT78), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n218), .A2(KEYINPUT79), .A3(KEYINPUT2), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT79), .B1(new_n218), .B2(KEYINPUT2), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n207), .B(new_n208), .C1(new_n217), .C2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT74), .ZN(new_n225));
  AND2_X1   g024(.A1(G211gat), .A2(G218gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G211gat), .A2(G218gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G211gat), .ZN(new_n229));
  INV_X1    g028(.A(G218gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G211gat), .A2(G218gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(KEYINPUT74), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n228), .A2(new_n233), .A3(KEYINPUT73), .ZN(new_n234));
  NAND2_X1  g033(.A1(G197gat), .A2(G204gat), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(G197gat), .A2(G204gat), .ZN(new_n237));
  OAI22_X1  g036(.A1(new_n236), .A2(new_n237), .B1(new_n226), .B2(KEYINPUT22), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n234), .B(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n203), .B1(new_n224), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n239), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT3), .B1(new_n241), .B2(new_n223), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n210), .A2(new_n212), .ZN(new_n243));
  AND2_X1   g042(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n244));
  NOR2_X1   g043(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n215), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n219), .A2(new_n220), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n240), .B1(new_n242), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n208), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n228), .A2(new_n233), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT29), .B1(new_n253), .B2(new_n238), .ZN(new_n254));
  INV_X1    g053(.A(G197gat), .ZN(new_n255));
  INV_X1    g054(.A(G204gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT22), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n257), .A2(new_n235), .B1(new_n258), .B2(new_n232), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(new_n228), .A3(new_n233), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n252), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT85), .B1(new_n261), .B2(new_n250), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n226), .A2(new_n227), .A3(new_n225), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT74), .B1(new_n231), .B2(new_n232), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n238), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(new_n223), .A3(new_n260), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n208), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n207), .B1(new_n217), .B2(new_n221), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n224), .A2(new_n239), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n262), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n272), .A2(new_n273), .A3(new_n203), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(new_n272), .B2(new_n203), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n251), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G22gat), .ZN(new_n277));
  INV_X1    g076(.A(G22gat), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n278), .B(new_n251), .C1(new_n274), .C2(new_n275), .ZN(new_n279));
  XNOR2_X1  g078(.A(G78gat), .B(G106gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT31), .B(G50gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n277), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(new_n277), .B2(new_n279), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G127gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G134gat), .ZN(new_n287));
  INV_X1    g086(.A(G134gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G127gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT70), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT1), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n287), .A2(new_n289), .A3(new_n291), .A4(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n295));
  INV_X1    g094(.A(G120gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G113gat), .ZN(new_n297));
  INV_X1    g096(.A(G113gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G120gat), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n295), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G113gat), .B(G120gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n295), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n286), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n306));
  XNOR2_X1  g105(.A(G127gat), .B(G134gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n297), .A2(new_n299), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n290), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n301), .A2(new_n303), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(KEYINPUT23), .ZN(new_n314));
  INV_X1    g113(.A(G169gat), .ZN(new_n315));
  INV_X1    g114(.A(G176gat), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT23), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT65), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G183gat), .A2(G190gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT24), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G183gat), .ZN(new_n322));
  INV_X1    g121(.A(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n321), .A2(new_n324), .A3(KEYINPUT65), .A4(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n318), .A2(KEYINPUT25), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT25), .B1(new_n318), .B2(new_n326), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n313), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT26), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n331), .A3(new_n312), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n313), .A2(KEYINPUT26), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n319), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n322), .A2(KEYINPUT27), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT27), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G183gat), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT67), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT27), .B(G183gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT67), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT28), .A4(new_n323), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n323), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n334), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n311), .B1(new_n329), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT64), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n318), .A2(new_n326), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n318), .A2(KEYINPUT25), .A3(new_n326), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n334), .ZN(new_n355));
  INV_X1    g154(.A(new_n345), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n335), .A2(new_n337), .A3(KEYINPUT67), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n323), .A2(KEYINPUT28), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n357), .A2(new_n338), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n355), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n307), .B(new_n361), .C1(new_n302), .C2(new_n295), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n309), .A2(KEYINPUT69), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n287), .A2(new_n289), .A3(new_n306), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n304), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n302), .A2(KEYINPUT1), .ZN(new_n366));
  OAI22_X1  g165(.A1(new_n362), .A2(new_n363), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n354), .A2(new_n360), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n347), .A2(new_n349), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT33), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G15gat), .B(G43gat), .Z(new_n373));
  XNOR2_X1  g172(.A(G71gat), .B(G99gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n375), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n369), .B(KEYINPUT32), .C1(new_n371), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT71), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT34), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n347), .A2(new_n368), .ZN(new_n382));
  INV_X1    g181(.A(new_n349), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI211_X1 g183(.A(KEYINPUT34), .B(new_n349), .C1(new_n347), .C2(new_n368), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n386), .A2(new_n376), .A3(new_n378), .ZN(new_n387));
  INV_X1    g186(.A(new_n384), .ZN(new_n388));
  INV_X1    g187(.A(new_n385), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n376), .A2(new_n378), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n380), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n379), .A2(KEYINPUT71), .A3(new_n386), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n202), .B1(new_n285), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT76), .ZN(new_n395));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n329), .A2(new_n346), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n395), .B(new_n396), .C1(new_n397), .C2(KEYINPUT29), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT29), .B1(new_n354), .B2(new_n360), .ZN(new_n399));
  INV_X1    g198(.A(new_n396), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT76), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n396), .B(KEYINPUT75), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n402), .B1(new_n329), .B2(new_n346), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n398), .A2(new_n401), .A3(new_n241), .A4(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n399), .A2(new_n402), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n397), .A2(new_n396), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n239), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G8gat), .B(G36gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n409), .B(new_n410), .Z(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n404), .A2(new_n407), .A3(new_n411), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(KEYINPUT30), .A3(new_n414), .ZN(new_n415));
  OR3_X1    g214(.A1(new_n408), .A2(KEYINPUT30), .A3(new_n412), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT81), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n311), .A2(new_n250), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT81), .B1(new_n367), .B2(new_n269), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n367), .A2(new_n269), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n419), .A2(new_n420), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT3), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n367), .B(new_n222), .C1(new_n250), .C2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n311), .A2(new_n250), .A3(KEYINPUT4), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n429), .A2(new_n423), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n422), .A2(KEYINPUT82), .A3(new_n424), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n427), .A2(KEYINPUT5), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G1gat), .B(G29gat), .Z(new_n436));
  XNOR2_X1  g235(.A(G57gat), .B(G85gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  AOI21_X1  g239(.A(KEYINPUT4), .B1(new_n311), .B2(new_n250), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n419), .A2(new_n420), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(KEYINPUT4), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT5), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n431), .A2(new_n444), .A3(new_n423), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n435), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n446), .ZN(new_n452));
  INV_X1    g251(.A(new_n440), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n447), .A2(KEYINPUT84), .A3(new_n448), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n451), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(KEYINPUT6), .A3(new_n453), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n417), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n379), .A2(KEYINPUT71), .A3(new_n386), .ZN(new_n459));
  INV_X1    g258(.A(new_n386), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n379), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n386), .A2(new_n376), .A3(new_n378), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n459), .B1(new_n463), .B2(new_n380), .ZN(new_n464));
  INV_X1    g263(.A(new_n282), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n272), .A2(new_n203), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT86), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n272), .A2(new_n273), .A3(new_n203), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n278), .B1(new_n469), .B2(new_n251), .ZN(new_n470));
  INV_X1    g269(.A(new_n279), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n277), .A2(new_n279), .A3(new_n282), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n464), .A2(new_n474), .A3(KEYINPUT91), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n394), .A2(new_n458), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT35), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n415), .A2(new_n416), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n422), .A2(KEYINPUT82), .A3(new_n424), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT82), .B1(new_n422), .B2(new_n424), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n431), .A2(new_n423), .A3(new_n432), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n444), .B1(new_n485), .B2(new_n429), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n484), .A2(new_n486), .B1(new_n443), .B2(new_n445), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT6), .B1(new_n487), .B2(new_n440), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n453), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n452), .A2(KEYINPUT87), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n457), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n452), .A2(KEYINPUT89), .A3(KEYINPUT6), .A4(new_n453), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(KEYINPUT88), .B(new_n488), .C1(new_n490), .C2(new_n491), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n494), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n481), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n477), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT40), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n422), .A2(new_n424), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT39), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n443), .A2(new_n431), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n505), .B1(new_n424), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n508), .A3(new_n424), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n440), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n503), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n506), .A2(new_n424), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(KEYINPUT39), .A3(new_n504), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n513), .A2(KEYINPUT40), .A3(new_n440), .A4(new_n509), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n511), .B(new_n514), .C1(new_n490), .C2(new_n491), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n474), .B1(new_n515), .B2(new_n478), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n411), .B1(new_n408), .B2(KEYINPUT37), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT90), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT37), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n404), .A2(new_n521), .A3(new_n407), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n518), .B2(KEYINPUT90), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT38), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n398), .A2(new_n401), .A3(new_n239), .A4(new_n403), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n405), .A2(new_n406), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n525), .B(KEYINPUT37), .C1(new_n239), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n411), .A2(KEYINPUT38), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n522), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(new_n414), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n517), .B1(new_n530), .B2(new_n500), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n456), .A2(new_n457), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n478), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n464), .A2(KEYINPUT36), .ZN(new_n534));
  XOR2_X1   g333(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n535));
  NAND2_X1  g334(.A1(new_n463), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n533), .A2(new_n285), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n502), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT92), .B(G197gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT11), .B(G169gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT12), .Z(new_n545));
  NAND2_X1  g344(.A1(G29gat), .A2(G36gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT93), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR3_X1   g348(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(KEYINPUT15), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(KEYINPUT95), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n546), .B(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n554), .A2(new_n558), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n550), .A2(KEYINPUT94), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n550), .A2(KEYINPUT94), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n549), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n553), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT17), .ZN(new_n566));
  XNOR2_X1  g365(.A(G15gat), .B(G22gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT16), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n568), .B2(G1gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(G1gat), .B2(new_n567), .ZN(new_n570));
  INV_X1    g369(.A(G8gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G229gat), .A2(G233gat), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n572), .A2(KEYINPUT96), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(KEYINPUT96), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n565), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT18), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n574), .B(KEYINPUT13), .Z(new_n581));
  INV_X1    g380(.A(new_n577), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n565), .B1(new_n575), .B2(new_n576), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n578), .A2(new_n579), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n545), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  INV_X1    g387(.A(new_n545), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n588), .A2(new_n580), .A3(new_n584), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT101), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT101), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(G85gat), .A3(G92gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n595), .A3(KEYINPUT7), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT102), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n596), .B(new_n597), .C1(KEYINPUT7), .C2(new_n592), .ZN(new_n599));
  NAND2_X1  g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  INV_X1    g399(.A(G85gat), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(KEYINPUT8), .A2(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  OR3_X1    g404(.A1(new_n604), .A2(KEYINPUT103), .A3(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n605), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(KEYINPUT103), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n566), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n606), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n565), .ZN(new_n612));
  NAND3_X1  g411(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  AND2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G134gat), .B(G162gat), .Z(new_n619));
  AOI21_X1  g418(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT104), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n621), .B(KEYINPUT104), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n616), .B2(new_n617), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  OR2_X1    g428(.A1(G71gat), .A2(G78gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G57gat), .B(G64gat), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT9), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT97), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n630), .A2(new_n629), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n635), .B(new_n636), .C1(new_n632), .C2(new_n631), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n629), .B1(new_n630), .B2(new_n632), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n639));
  INV_X1    g438(.A(G57gat), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n640), .B2(G64gat), .ZN(new_n641));
  INV_X1    g440(.A(G64gat), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n641), .B1(G57gat), .B2(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n639), .A2(new_n640), .A3(G64gat), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n638), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n634), .A2(new_n637), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT99), .B(KEYINPUT21), .Z(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(G127gat), .B(G155gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT20), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(G183gat), .B(G211gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n646), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n575), .A2(new_n576), .B1(KEYINPUT21), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT100), .B(KEYINPUT19), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n655), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n628), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n607), .A2(new_n608), .A3(new_n656), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n609), .A2(new_n646), .A3(new_n606), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n611), .A2(KEYINPUT10), .A3(new_n656), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n663), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT106), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G120gat), .B(G148gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(G176gat), .B(G204gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(KEYINPUT106), .B(new_n676), .C1(new_n671), .C2(new_n672), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n661), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n539), .A2(new_n591), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n539), .A2(KEYINPUT107), .A3(new_n591), .A4(new_n683), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n532), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g490(.A(KEYINPUT16), .B(G8gat), .Z(new_n692));
  NAND3_X1  g491(.A1(new_n688), .A2(new_n417), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n693), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT108), .B1(new_n697), .B2(KEYINPUT42), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n571), .B1(new_n688), .B2(new_n417), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n693), .B1(new_n699), .B2(new_n695), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n696), .B1(new_n698), .B2(new_n700), .ZN(G1325gat));
  INV_X1    g500(.A(G15gat), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n688), .A2(new_n702), .A3(new_n462), .A4(new_n461), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n534), .A2(new_n536), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n686), .B2(new_n687), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n705), .B2(new_n702), .ZN(G1326gat));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n285), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT43), .B(G22gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  NAND2_X1  g508(.A1(new_n627), .A2(KEYINPUT109), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n624), .A2(new_n711), .A3(new_n626), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n499), .A2(new_n498), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n440), .B1(new_n452), .B2(KEYINPUT87), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n487), .A2(new_n489), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT88), .B1(new_n718), .B2(new_n488), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n529), .A2(new_n414), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n518), .A2(KEYINPUT90), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(new_n519), .A3(new_n522), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n721), .B1(new_n723), .B2(KEYINPUT38), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n516), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n704), .B1(new_n474), .B2(new_n458), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n476), .A2(KEYINPUT35), .B1(new_n500), .B2(new_n481), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n714), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n627), .B1(new_n502), .B2(new_n538), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n681), .A2(new_n591), .A3(new_n660), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G29gat), .B1(new_n736), .B2(new_n532), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n730), .A2(new_n591), .A3(new_n660), .A4(new_n681), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n532), .A2(G29gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n739), .A2(new_n738), .A3(new_n740), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n737), .A2(new_n741), .A3(new_n742), .ZN(G1328gat));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR4_X1   g545(.A1(new_n739), .A2(G36gat), .A3(new_n478), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G36gat), .B1(new_n736), .B2(new_n478), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(G1329gat));
  INV_X1    g550(.A(new_n704), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n735), .A2(G43gat), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n739), .A2(new_n463), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(G43gat), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT47), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n753), .B(new_n757), .C1(G43gat), .C2(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1330gat));
  INV_X1    g558(.A(G50gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n739), .B2(new_n474), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n285), .A2(G50gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n736), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g563(.A(new_n591), .ZN(new_n765));
  AND4_X1   g564(.A1(new_n539), .A2(new_n765), .A3(new_n661), .A4(new_n680), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n689), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n417), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT49), .B(G64gat), .Z(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(G1333gat));
  NAND2_X1  g571(.A1(new_n766), .A2(new_n752), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n463), .A2(G71gat), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n773), .A2(G71gat), .B1(new_n766), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n766), .A2(new_n285), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  INV_X1    g577(.A(new_n660), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n591), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n628), .B(new_n780), .C1(new_n727), .C2(new_n728), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n539), .A2(KEYINPUT51), .A3(new_n628), .A4(new_n780), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n681), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(new_n601), .A3(new_n689), .ZN(new_n786));
  INV_X1    g585(.A(new_n780), .ZN(new_n787));
  NOR4_X1   g586(.A1(new_n733), .A2(new_n532), .A3(new_n681), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n788), .B2(new_n601), .ZN(G1336gat));
  NAND2_X1  g588(.A1(new_n783), .A2(new_n784), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n681), .A2(new_n478), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(G92gat), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n733), .A2(new_n787), .A3(new_n792), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(G92gat), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n795), .A2(new_n602), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n783), .A2(new_n784), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n781), .A2(KEYINPUT111), .A3(new_n782), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n802), .A2(new_n793), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n805), .ZN(G1337gat));
  NAND3_X1  g605(.A1(new_n732), .A2(new_n680), .A3(new_n780), .ZN(new_n807));
  OAI21_X1  g606(.A(G99gat), .B1(new_n807), .B2(new_n704), .ZN(new_n808));
  INV_X1    g607(.A(new_n785), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n463), .A2(G99gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(G1338gat));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812));
  XOR2_X1   g611(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n813));
  NOR2_X1   g612(.A1(new_n474), .A2(G106gat), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n785), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n732), .A2(new_n285), .A3(new_n680), .A4(new_n780), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G106gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n680), .A2(new_n814), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n803), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n812), .B(new_n818), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n815), .A2(new_n817), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n822), .B1(new_n817), .B2(new_n820), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT114), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(G1339gat));
  NOR2_X1   g626(.A1(new_n682), .A2(new_n591), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n669), .A2(new_n670), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n662), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n669), .A2(new_n663), .A3(new_n670), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n676), .B1(new_n671), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n585), .A2(new_n586), .A3(new_n545), .ZN(new_n839));
  INV_X1    g638(.A(new_n574), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n566), .A2(new_n572), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n582), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g643(.A(KEYINPUT115), .B(new_n840), .C1(new_n841), .C2(new_n582), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n582), .A2(new_n583), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n581), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n839), .B1(new_n544), .B2(new_n847), .ZN(new_n848));
  OR3_X1    g647(.A1(new_n671), .A2(new_n672), .A3(new_n677), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n835), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n838), .A2(new_n848), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n713), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n848), .A2(new_n679), .A3(new_n678), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n838), .A2(new_n591), .A3(new_n849), .A4(new_n850), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n680), .A2(KEYINPUT116), .A3(new_n848), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n852), .B1(new_n858), .B2(new_n713), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n829), .B1(new_n859), .B2(new_n779), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n860), .A2(new_n474), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n689), .A2(new_n478), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n463), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(new_n298), .A3(new_n765), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n394), .A2(new_n475), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n860), .A2(new_n689), .A3(new_n478), .A4(new_n866), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(new_n765), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n865), .B1(new_n868), .B2(new_n298), .ZN(G1340gat));
  OAI21_X1  g668(.A(new_n296), .B1(new_n867), .B2(new_n681), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n680), .A2(G120gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n864), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT117), .ZN(G1341gat));
  OAI21_X1  g672(.A(G127gat), .B1(new_n864), .B2(new_n660), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n779), .A2(new_n286), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n867), .B2(new_n875), .ZN(G1342gat));
  OAI21_X1  g675(.A(G134gat), .B1(new_n864), .B2(new_n627), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n627), .A2(G134gat), .A3(new_n417), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n860), .A2(new_n689), .A3(new_n866), .A4(new_n878), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n877), .A2(KEYINPUT118), .A3(new_n880), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1343gat));
  NOR2_X1   g685(.A1(new_n752), .A2(new_n862), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n860), .B2(new_n285), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n474), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n847), .A2(new_n544), .ZN(new_n892));
  AND4_X1   g691(.A1(new_n590), .A2(new_n678), .A3(new_n892), .A4(new_n679), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n836), .A2(KEYINPUT119), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n833), .A2(new_n895), .A3(new_n835), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n837), .A3(new_n896), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n850), .A2(new_n591), .A3(new_n849), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n893), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n628), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n660), .B1(new_n900), .B2(new_n852), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n891), .B1(new_n901), .B2(new_n829), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n591), .B(new_n887), .C1(new_n888), .C2(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n903), .A2(G141gat), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n860), .A2(new_n689), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n752), .A2(new_n474), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n478), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n765), .A2(G141gat), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT58), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n903), .A2(G141gat), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n912), .B(new_n913), .C1(new_n907), .C2(new_n909), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n911), .A2(new_n914), .ZN(G1344gat));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n681), .B1(new_n887), .B2(KEYINPUT121), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(KEYINPUT121), .B2(new_n887), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n850), .A2(new_n849), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n919), .A2(new_n628), .A3(new_n848), .A4(new_n838), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n899), .B2(new_n628), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n828), .B1(new_n921), .B2(new_n660), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n889), .B1(new_n922), .B2(new_n474), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n860), .A2(new_n890), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n211), .B1(new_n925), .B2(KEYINPUT122), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n850), .A2(new_n591), .A3(new_n849), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT55), .B1(new_n836), .B2(KEYINPUT119), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n896), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n627), .B1(new_n930), .B2(new_n893), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n779), .B1(new_n931), .B2(new_n920), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n285), .B1(new_n932), .B2(new_n828), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n933), .A2(new_n889), .B1(new_n860), .B2(new_n890), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n927), .B1(new_n934), .B2(new_n918), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n916), .B1(new_n926), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n916), .A2(G148gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n888), .A2(new_n902), .ZN(new_n938));
  INV_X1    g737(.A(new_n887), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n937), .B1(new_n940), .B2(new_n680), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n681), .A2(G148gat), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n907), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(KEYINPUT120), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n907), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  OAI22_X1  g746(.A1(new_n936), .A2(new_n941), .B1(new_n945), .B2(new_n947), .ZN(G1345gat));
  NOR2_X1   g747(.A1(new_n907), .A2(new_n660), .ZN(new_n949));
  AOI21_X1  g748(.A(G155gat), .B1(new_n949), .B2(KEYINPUT123), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n951), .B1(new_n907), .B2(new_n660), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n779), .A2(G155gat), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT124), .ZN(new_n954));
  AOI22_X1  g753(.A1(new_n950), .A2(new_n952), .B1(new_n940), .B2(new_n954), .ZN(G1346gat));
  INV_X1    g754(.A(new_n713), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n956), .B(new_n887), .C1(new_n888), .C2(new_n902), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G162gat), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n627), .A2(G162gat), .A3(new_n417), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n905), .A2(new_n906), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n958), .A2(KEYINPUT125), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1347gat));
  NOR3_X1   g764(.A1(new_n689), .A2(new_n478), .A3(new_n463), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n861), .A2(new_n966), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n967), .A2(new_n315), .A3(new_n765), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n860), .A2(new_n532), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n969), .A2(new_n866), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(new_n417), .A3(new_n591), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n968), .B1(new_n971), .B2(new_n315), .ZN(G1348gat));
  NAND3_X1  g771(.A1(new_n970), .A2(new_n316), .A3(new_n791), .ZN(new_n973));
  OAI21_X1  g772(.A(G176gat), .B1(new_n967), .B2(new_n681), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(G1349gat));
  OAI21_X1  g774(.A(G183gat), .B1(new_n967), .B2(new_n660), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n969), .A2(new_n417), .A3(new_n866), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n779), .A2(new_n339), .A3(new_n341), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(KEYINPUT60), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT60), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n976), .B(new_n982), .C1(new_n978), .C2(new_n979), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n981), .A2(new_n983), .ZN(G1350gat));
  NAND2_X1  g783(.A1(new_n956), .A2(new_n323), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n978), .A2(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n861), .A2(new_n628), .A3(new_n966), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n987), .B1(new_n988), .B2(G190gat), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n988), .A2(G190gat), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(KEYINPUT61), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n991), .B1(new_n994), .B2(new_n995), .ZN(G1351gat));
  NAND2_X1  g795(.A1(new_n923), .A2(new_n924), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n689), .A2(new_n478), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(new_n704), .A3(new_n998), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n999), .A2(new_n255), .A3(new_n765), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n752), .A2(new_n474), .A3(new_n478), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n969), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g801(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g802(.A(G197gat), .B1(new_n1003), .B2(new_n591), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n1000), .A2(new_n1004), .ZN(G1352gat));
  NAND2_X1  g804(.A1(new_n680), .A2(new_n256), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n1007));
  OAI22_X1  g806(.A1(new_n1002), .A2(new_n1006), .B1(new_n1007), .B2(KEYINPUT62), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1008), .B1(KEYINPUT127), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g809(.A(G204gat), .B1(new_n999), .B2(new_n681), .ZN(new_n1011));
  OAI211_X1 g810(.A(new_n1007), .B(KEYINPUT62), .C1(new_n1002), .C2(new_n1006), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(G1353gat));
  NAND3_X1  g812(.A1(new_n1003), .A2(new_n229), .A3(new_n779), .ZN(new_n1014));
  NAND4_X1  g813(.A1(new_n997), .A2(new_n704), .A3(new_n779), .A4(new_n998), .ZN(new_n1015));
  AND3_X1   g814(.A1(new_n1015), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1016));
  AOI21_X1  g815(.A(KEYINPUT63), .B1(new_n1015), .B2(G211gat), .ZN(new_n1017));
  OAI21_X1  g816(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(G1354gat));
  OAI21_X1  g817(.A(G218gat), .B1(new_n999), .B2(new_n627), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1003), .A2(new_n230), .A3(new_n956), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1019), .A2(new_n1020), .ZN(G1355gat));
endmodule


