//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n569, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n624, new_n627, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G567), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(new_n457));
  INV_X1    g032(.A(new_n451), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n457), .B1(G2106), .B2(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G101), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI211_X1 g043(.A(KEYINPUT67), .B(new_n465), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n470), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  OAI221_X1 g052(.A(new_n462), .B1(new_n463), .B2(new_n466), .C1(new_n469), .C2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n479));
  OR2_X1    g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n479), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT69), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n464), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  OAI22_X1  g065(.A1(new_n488), .A2(new_n489), .B1(new_n466), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n487), .A2(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n471), .A2(new_n473), .A3(G138), .A4(new_n465), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n464), .A2(KEYINPUT4), .A3(G138), .A4(new_n465), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n464), .A2(G126), .A3(G2105), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G651), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n510), .B(KEYINPUT5), .C1(new_n511), .C2(KEYINPUT72), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n513), .B1(KEYINPUT71), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  AOI21_X1  g090(.A(KEYINPUT71), .B1(new_n515), .B2(G543), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n512), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT73), .B1(new_n509), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n504), .A2(new_n506), .B1(new_n503), .B2(G651), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT5), .B1(new_n510), .B2(new_n511), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n510), .B1(new_n511), .B2(KEYINPUT72), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n519), .A2(new_n520), .A3(new_n523), .A4(new_n512), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT74), .B(G88), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n518), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n519), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  NAND2_X1  g104(.A1(G75), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G62), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n517), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT75), .ZN(new_n533));
  AND3_X1   g108(.A1(new_n532), .A2(new_n533), .A3(G651), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n533), .B1(new_n532), .B2(G651), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n526), .B(new_n529), .C1(new_n534), .C2(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  AND2_X1   g112(.A1(new_n518), .A2(new_n524), .ZN(new_n538));
  OR2_X1    g113(.A1(KEYINPUT76), .A2(G89), .ZN(new_n539));
  NAND2_X1  g114(.A1(KEYINPUT76), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT7), .ZN(new_n542));
  NAND2_X1  g117(.A1(G76), .A2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n543), .B2(new_n505), .ZN(new_n544));
  INV_X1    g119(.A(G51), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n527), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G63), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n517), .A2(new_n547), .B1(new_n542), .B2(new_n543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n546), .B1(G651), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n541), .A2(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n517), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT77), .ZN(new_n556));
  INV_X1    g131(.A(G52), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n518), .A2(new_n524), .ZN(new_n559));
  OAI221_X1 g134(.A(new_n556), .B1(new_n557), .B2(new_n527), .C1(new_n558), .C2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  NAND2_X1  g136(.A1(new_n538), .A2(G81), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n517), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(G43), .A2(new_n528), .B1(new_n565), .B2(G651), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G188));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT78), .B1(new_n559), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n518), .A2(new_n576), .A3(G91), .A4(new_n524), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT79), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n517), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(KEYINPUT80), .A3(G651), .ZN(new_n586));
  INV_X1    g161(.A(G53), .ZN(new_n587));
  OR3_X1    g162(.A1(new_n527), .A2(KEYINPUT9), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT9), .B1(new_n527), .B2(new_n587), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n585), .A2(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n578), .A2(new_n590), .ZN(G299));
  INV_X1    g166(.A(G74), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n505), .B1(new_n517), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n528), .B2(G49), .ZN(new_n594));
  INV_X1    g169(.A(G87), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n559), .B2(new_n595), .ZN(G288));
  NAND2_X1  g171(.A1(new_n538), .A2(G86), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n517), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(G48), .A2(new_n528), .B1(new_n600), .B2(G651), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n538), .A2(G85), .ZN(new_n603));
  XNOR2_X1  g178(.A(KEYINPUT81), .B(G47), .ZN(new_n604));
  NAND2_X1  g179(.A1(G72), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n517), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n528), .A2(new_n604), .B1(new_n607), .B2(G651), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n603), .A2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT82), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n517), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(G54), .A2(new_n528), .B1(new_n614), .B2(G651), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  AND3_X1   g191(.A1(new_n518), .A2(G92), .A3(new_n524), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n617), .A2(KEYINPUT10), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(KEYINPUT10), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n610), .B1(G868), .B2(new_n620), .ZN(G284));
  OAI21_X1  g196(.A(new_n610), .B1(G868), .B2(new_n620), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  INV_X1    g198(.A(G299), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G297));
  OAI21_X1  g200(.A(new_n623), .B1(new_n624), .B2(G868), .ZN(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n620), .B1(new_n627), .B2(G860), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT83), .Z(G148));
  INV_X1    g204(.A(new_n620), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n630), .A2(G559), .ZN(new_n631));
  MUX2_X1   g206(.A(new_n567), .B(new_n631), .S(G868), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT84), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g209(.A1(new_n474), .A2(G2105), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G2104), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n635), .A2(G135), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n474), .A2(new_n465), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(G123), .ZN(new_n644));
  OR2_X1    g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n645), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n642), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2096), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n640), .A2(new_n641), .A3(new_n648), .ZN(G156));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT86), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2451), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n654), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT87), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2454), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(G14), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n666), .B2(new_n662), .ZN(G401));
  INV_X1    g243(.A(KEYINPUT18), .ZN(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n672), .B2(KEYINPUT18), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n675), .B(new_n677), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT20), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n685), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n685), .B2(new_n691), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT88), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT90), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n698), .B(new_n699), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n696), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT91), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n700), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n696), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n703), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(new_n708), .ZN(G229));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(G5), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G301), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G1961), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n635), .A2(G140), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n643), .A2(G128), .ZN(new_n716));
  OR2_X1    g291(.A1(G104), .A2(G2105), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n717), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G29), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT92), .B(G29), .Z(new_n721));
  INV_X1    g296(.A(G26), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT28), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G2067), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT99), .B(G28), .Z(new_n729));
  AOI21_X1  g304(.A(G29), .B1(new_n729), .B2(KEYINPUT30), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(KEYINPUT30), .B2(new_n729), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT31), .B(G11), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n647), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n721), .ZN(new_n735));
  NAND2_X1  g310(.A1(G162), .A2(new_n721), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n721), .A2(G35), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(KEYINPUT29), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT29), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n736), .A2(new_n740), .A3(new_n737), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n728), .B(new_n735), .C1(new_n742), .C2(G2090), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n721), .A2(G27), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n721), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT102), .B(G2078), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n714), .A2(new_n743), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n739), .A2(G2090), .A3(new_n741), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(KEYINPUT103), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(KEYINPUT103), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n710), .A2(G21), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G286), .B2(G16), .ZN(new_n753));
  INV_X1    g328(.A(G1966), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n750), .A2(new_n751), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT94), .B(G16), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G19), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n567), .B2(new_n759), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G1341), .Z(new_n762));
  NAND3_X1  g337(.A1(new_n748), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G4), .A2(G16), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n620), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT96), .B(G1348), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n758), .A2(G20), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT23), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G299), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1956), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n763), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G29), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G33), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT25), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G139), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n778), .B1(new_n466), .B2(new_n779), .C1(new_n780), .C2(new_n465), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n775), .B1(new_n782), .B2(new_n774), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT97), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2072), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n480), .A2(G29), .A3(new_n481), .ZN(new_n786));
  INV_X1    g361(.A(new_n721), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT24), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(G34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(G34), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n786), .A2(G2084), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n774), .A2(G32), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n635), .A2(G141), .B1(G105), .B2(new_n461), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n643), .A2(G129), .ZN(new_n795));
  NAND3_X1  g370(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT26), .Z(new_n797));
  AND3_X1   g372(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n793), .B1(new_n798), .B2(new_n774), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT27), .B(G1996), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n785), .A2(new_n792), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT98), .ZN(new_n804));
  AOI21_X1  g379(.A(G2084), .B1(new_n786), .B2(new_n791), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n712), .A2(new_n713), .B1(new_n799), .B2(new_n801), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT101), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n806), .A2(new_n807), .A3(KEYINPUT101), .A4(new_n808), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n773), .A2(new_n804), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(KEYINPUT95), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n721), .A2(G25), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n635), .A2(G131), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n643), .A2(G119), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n465), .A2(G107), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT93), .Z(new_n823));
  AOI21_X1  g398(.A(new_n817), .B1(new_n823), .B2(new_n721), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G1991), .Z(new_n825));
  XOR2_X1   g400(.A(new_n824), .B(new_n825), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n758), .A2(G24), .ZN(new_n827));
  INV_X1    g402(.A(G290), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(new_n758), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n829), .A2(G1986), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n829), .A2(G1986), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n826), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(G6), .A2(G16), .ZN(new_n833));
  INV_X1    g408(.A(G305), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(G16), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT32), .B(G1981), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n835), .B(new_n836), .Z(new_n837));
  NOR2_X1   g412(.A1(new_n759), .A2(G22), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G166), .B2(new_n759), .ZN(new_n839));
  INV_X1    g414(.A(G1971), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  MUX2_X1   g416(.A(G23), .B(G288), .S(G16), .Z(new_n842));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G1976), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n842), .B(KEYINPUT33), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(G1976), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n837), .B(new_n841), .C1(new_n846), .C2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n832), .B1(new_n849), .B2(KEYINPUT34), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT34), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n837), .A2(new_n841), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n844), .B(new_n845), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n816), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n853), .A3(new_n851), .ZN(new_n857));
  INV_X1    g432(.A(new_n816), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n832), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n814), .B1(new_n855), .B2(new_n859), .ZN(G311));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n861));
  AOI211_X1 g436(.A(new_n861), .B(new_n814), .C1(new_n855), .C2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n855), .A2(new_n859), .ZN(new_n863));
  INV_X1    g438(.A(new_n814), .ZN(new_n864));
  AOI21_X1  g439(.A(KEYINPUT104), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n862), .A2(new_n865), .ZN(G150));
  NAND2_X1  g441(.A1(new_n538), .A2(G93), .ZN(new_n867));
  NAND2_X1  g442(.A1(G80), .A2(G543), .ZN(new_n868));
  INV_X1    g443(.A(G67), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n517), .B2(new_n869), .ZN(new_n870));
  AOI22_X1  g445(.A1(G55), .A2(new_n528), .B1(new_n870), .B2(G651), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(G860), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  OAI21_X1  g449(.A(KEYINPUT105), .B1(new_n630), .B2(new_n627), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n630), .A2(KEYINPUT105), .A3(new_n627), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT38), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT38), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n880), .A3(new_n875), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n562), .A2(new_n566), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n882), .A2(new_n872), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n872), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n878), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n885), .B1(new_n878), .B2(new_n881), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT39), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n888), .A2(G860), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT39), .B1(new_n886), .B2(new_n887), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n874), .B1(new_n892), .B2(new_n893), .ZN(G145));
  NAND2_X1  g469(.A1(new_n482), .A2(new_n734), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n480), .A2(new_n481), .A3(new_n647), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(G162), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G162), .B1(new_n895), .B2(new_n896), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT110), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n897), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n497), .A2(new_n499), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT107), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT107), .B1(new_n495), .B2(new_n496), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(new_n719), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n909), .A2(new_n798), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n798), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n781), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n643), .A2(G130), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n465), .A2(G118), .ZN(new_n915));
  OAI21_X1  g490(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(G142), .B2(new_n635), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n637), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(new_n823), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n910), .A2(new_n782), .A3(new_n911), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n913), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n900), .A2(new_n903), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT111), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n920), .B1(new_n913), .B2(new_n921), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI211_X1 g503(.A(KEYINPUT108), .B(new_n920), .C1(new_n913), .C2(new_n921), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n924), .B(new_n925), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT111), .B1(new_n931), .B2(new_n923), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g508(.A1(new_n922), .A2(KEYINPUT109), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n922), .A2(KEYINPUT109), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n934), .B(new_n935), .C1(new_n928), .C2(new_n929), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n898), .A2(new_n899), .ZN(new_n937));
  AOI21_X1  g512(.A(G37), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n933), .A2(KEYINPUT40), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT40), .B1(new_n933), .B2(new_n938), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(G395));
  NOR2_X1   g516(.A1(new_n872), .A2(G868), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n631), .B(new_n885), .Z(new_n943));
  NAND2_X1  g518(.A1(new_n630), .A2(G299), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n624), .A2(new_n620), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT41), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT41), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n943), .A2(new_n946), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT113), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n951), .B(new_n955), .C1(new_n943), .C2(new_n946), .ZN(new_n956));
  XOR2_X1   g531(.A(G305), .B(G288), .Z(new_n957));
  XNOR2_X1  g532(.A(G290), .B(G303), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n957), .B(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n961));
  OR3_X1    g536(.A1(new_n960), .A2(KEYINPUT112), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n960), .B2(KEYINPUT112), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n954), .A2(new_n956), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n952), .A2(new_n953), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(new_n966), .A3(new_n955), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n942), .B1(new_n968), .B2(G868), .ZN(G295));
  AOI21_X1  g544(.A(new_n942), .B1(new_n968), .B2(G868), .ZN(G331));
  INV_X1    g545(.A(G37), .ZN(new_n971));
  OAI21_X1  g546(.A(G168), .B1(new_n883), .B2(new_n884), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n567), .A2(new_n867), .A3(new_n871), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n882), .A2(new_n872), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(G286), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G301), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n972), .A2(new_n975), .A3(G171), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n946), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n950), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(new_n982), .B2(new_n979), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n971), .B1(new_n983), .B2(new_n959), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n977), .A2(new_n978), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n947), .A2(new_n986), .A3(new_n949), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n946), .A2(KEYINPUT114), .A3(KEYINPUT41), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n960), .B1(new_n989), .B2(new_n981), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n984), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n946), .B1(new_n977), .B2(new_n978), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n950), .B2(new_n985), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n994), .B2(new_n960), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n983), .A2(new_n959), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT43), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT44), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n984), .A2(new_n990), .A3(KEYINPUT43), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n991), .B1(new_n995), .B2(new_n996), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n1002), .ZN(G397));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n1004));
  INV_X1    g579(.A(G8), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(G166), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n908), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT50), .ZN(new_n1012));
  OAI211_X1 g587(.A(G40), .B(new_n462), .C1(new_n466), .C2(new_n463), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n469), .B2(new_n477), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n500), .A2(new_n1010), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1015), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G2090), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1012), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n477), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n470), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1013), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n1018), .B2(KEYINPUT45), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n495), .A2(new_n496), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT107), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1384), .B1(new_n1032), .B2(new_n905), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT116), .B1(new_n1033), .B2(KEYINPUT45), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n908), .A2(KEYINPUT116), .A3(KEYINPUT45), .A4(new_n1010), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1027), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1021), .B1(new_n1037), .B2(new_n840), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1009), .B1(new_n1038), .B2(new_n1005), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT120), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(new_n1009), .C1(new_n1038), .C2(new_n1005), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1033), .A2(new_n1025), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(new_n1005), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  INV_X1    g622(.A(G1981), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n597), .A2(new_n1048), .A3(new_n601), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n597), .B2(new_n601), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1051), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(KEYINPUT49), .A3(new_n1049), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1046), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n594), .B(G1976), .C1(new_n559), .C2(new_n595), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1044), .A2(new_n1056), .A3(G8), .A4(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1044), .A2(G8), .A3(new_n845), .A4(G288), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1058), .B1(new_n1060), .B2(new_n1059), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n908), .A2(KEYINPUT45), .A3(new_n1010), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1035), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1971), .B1(new_n1067), .B2(new_n1027), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n908), .A2(new_n1016), .A3(new_n1010), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1016), .B1(new_n500), .B2(new_n1010), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1015), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(G2090), .ZN(new_n1073));
  OAI211_X1 g648(.A(G8), .B(new_n1008), .C1(new_n1068), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1026), .B1(new_n1066), .B2(new_n1035), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n1077), .A2(G1971), .B1(G2090), .B2(new_n1072), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1078), .A2(KEYINPUT117), .A3(G8), .A4(new_n1008), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1063), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1033), .A2(KEYINPUT45), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT45), .ZN(new_n1082));
  OAI221_X1 g657(.A(new_n1014), .B1(new_n477), .B2(new_n469), .C1(new_n1017), .C2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n754), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G2084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1069), .A2(new_n1071), .A3(new_n1085), .ZN(new_n1086));
  AOI211_X1 g661(.A(new_n1005), .B(G286), .C1(new_n1084), .C2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1043), .A2(new_n1080), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(KEYINPUT63), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1008), .B1(new_n1078), .B2(G8), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1080), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1080), .A2(new_n1093), .A3(KEYINPUT121), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1090), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1044), .A2(G2067), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1348), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n620), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1956), .B1(new_n1012), .B2(new_n1019), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT56), .B(G2072), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n1077), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n578), .B2(new_n590), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n578), .A2(new_n590), .A3(new_n1105), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1104), .A2(KEYINPUT122), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1077), .A2(new_n1103), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1102), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1109), .A2(new_n1110), .A3(KEYINPUT122), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1101), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1107), .A2(new_n1106), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1109), .A2(new_n1113), .A3(new_n1110), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n882), .A2(KEYINPUT124), .ZN(new_n1117));
  INV_X1    g692(.A(G1996), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1067), .A2(new_n1118), .A3(new_n1027), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT58), .B(G1341), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1044), .A2(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1119), .A2(KEYINPUT123), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT123), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1117), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(KEYINPUT59), .B(new_n1117), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1104), .B2(new_n1113), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1131));
  NOR4_X1   g706(.A1(new_n630), .A2(new_n1099), .A3(KEYINPUT60), .A4(new_n1100), .ZN(new_n1132));
  OR3_X1    g707(.A1(new_n1099), .A2(new_n620), .A3(new_n1100), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1101), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1132), .B1(new_n1134), .B2(KEYINPUT60), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1113), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1129), .B1(new_n1114), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1131), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1116), .B1(new_n1128), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1083), .B1(new_n1082), .B2(new_n1011), .ZN(new_n1140));
  OAI211_X1 g715(.A(G168), .B(new_n1086), .C1(new_n1140), .C2(G1966), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(G8), .ZN(new_n1142));
  AOI21_X1  g717(.A(G168), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT51), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n1145), .A3(G8), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1072), .A2(new_n713), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1081), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT53), .ZN(new_n1150));
  NOR4_X1   g725(.A1(new_n1013), .A2(new_n1023), .A3(new_n1150), .A4(G2078), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1067), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  AOI211_X1 g727(.A(G2078), .B(new_n1026), .C1(new_n1066), .C2(new_n1035), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1148), .B(new_n1152), .C1(new_n1153), .C2(KEYINPUT53), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(G171), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1148), .ZN(new_n1156));
  INV_X1    g731(.A(G2078), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1067), .A2(new_n1157), .A3(new_n1027), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1158), .B2(new_n1150), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1140), .A2(KEYINPUT53), .A3(new_n1157), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(G301), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1155), .A2(new_n1161), .A3(KEYINPUT54), .ZN(new_n1162));
  AND4_X1   g737(.A1(new_n1043), .A2(new_n1080), .A3(new_n1147), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n1164));
  AOI21_X1  g739(.A(G301), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT53), .B1(new_n1077), .B2(new_n1157), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1151), .B1(new_n1033), .B2(KEYINPUT45), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1066), .B2(new_n1035), .ZN(new_n1168));
  NOR4_X1   g743(.A1(new_n1166), .A2(new_n1168), .A3(G171), .A4(new_n1156), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1164), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT125), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1172), .B(new_n1164), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1139), .A2(new_n1163), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1177));
  NOR2_X1   g752(.A1(G288), .A2(G1976), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT119), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1050), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1046), .ZN(new_n1181));
  OAI22_X1  g756(.A1(new_n1176), .A2(new_n1063), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1144), .A2(new_n1183), .A3(new_n1146), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1165), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1043), .A2(new_n1080), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1182), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1098), .A2(new_n1175), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1081), .A2(new_n1025), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n798), .B(G1996), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n719), .B(new_n727), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1195), .B1(new_n825), .B2(new_n823), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(new_n825), .B2(new_n823), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(G1986), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1198), .B1(new_n1199), .B2(new_n828), .ZN(new_n1200));
  NOR2_X1   g775(.A1(G290), .A2(G1986), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT115), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1192), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1190), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1191), .B1(new_n798), .B2(new_n1194), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1205), .B(KEYINPUT126), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1191), .A2(G1996), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n1207), .B(KEYINPUT46), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT47), .Z(new_n1210));
  NAND2_X1  g785(.A1(new_n1202), .A2(new_n1192), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1211), .ZN(new_n1212));
  AOI22_X1  g787(.A1(new_n1212), .A2(KEYINPUT48), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1213), .B1(KEYINPUT48), .B2(new_n1212), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n823), .A2(new_n825), .ZN(new_n1215));
  OAI22_X1  g790(.A1(new_n1195), .A2(new_n1215), .B1(G2067), .B2(new_n719), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n1192), .ZN(new_n1217));
  AND3_X1   g792(.A1(new_n1210), .A2(new_n1214), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1204), .A2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g794(.A1(new_n994), .A2(new_n960), .ZN(new_n1221));
  OAI21_X1  g795(.A(KEYINPUT43), .B1(new_n984), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n989), .A2(new_n981), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n1223), .A2(new_n959), .ZN(new_n1224));
  NAND3_X1  g798(.A1(new_n1224), .A2(new_n995), .A3(new_n991), .ZN(new_n1225));
  NAND2_X1  g799(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g800(.A1(new_n681), .A2(G319), .A3(new_n682), .ZN(new_n1227));
  XNOR2_X1  g801(.A(new_n1227), .B(KEYINPUT127), .ZN(new_n1228));
  NOR2_X1   g802(.A1(G401), .A2(new_n1228), .ZN(new_n1229));
  AND3_X1   g803(.A1(new_n704), .A2(new_n708), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g804(.A1(new_n933), .A2(new_n938), .ZN(new_n1231));
  AND3_X1   g805(.A1(new_n1226), .A2(new_n1230), .A3(new_n1231), .ZN(G308));
  NAND3_X1  g806(.A1(new_n1226), .A2(new_n1230), .A3(new_n1231), .ZN(G225));
endmodule


