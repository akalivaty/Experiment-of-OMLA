//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n457));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(G125), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n457), .B1(new_n462), .B2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AOI211_X1 g039(.A(KEYINPUT66), .B(new_n464), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT67), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n469), .A2(new_n464), .A3(G101), .A4(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n464), .C1(new_n458), .C2(new_n459), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(KEYINPUT68), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  INV_X1    g053(.A(new_n459), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n464), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n464), .B1(new_n477), .B2(new_n481), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND2_X1  g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n479), .B2(new_n480), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n464), .C1(new_n458), .C2(new_n459), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(KEYINPUT71), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(G102), .B2(G2105), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT69), .B(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(new_n464), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n503), .A2(KEYINPUT69), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(KEYINPUT69), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n499), .B(G2105), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n502), .A2(G2104), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n494), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n498), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(G50), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(new_n516), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n515), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n516), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI221_X1 g101(.A(new_n523), .B1(new_n524), .B2(new_n525), .C1(new_n526), .C2(new_n518), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n527), .A2(new_n530), .ZN(G168));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n518), .A2(new_n532), .B1(new_n524), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n514), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G171));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  INV_X1    g113(.A(G43), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n518), .A2(new_n538), .B1(new_n524), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n514), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  AOI22_X1  g123(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT74), .B1(new_n549), .B2(new_n514), .ZN(new_n550));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  AND2_X1   g126(.A1(KEYINPUT5), .A2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(KEYINPUT5), .A2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(new_n557), .A3(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g134(.A1(KEYINPUT73), .A2(G53), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n516), .A2(G543), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n516), .A2(new_n563), .A3(G543), .A4(new_n560), .ZN(new_n564));
  INV_X1    g139(.A(new_n518), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n562), .A2(new_n564), .B1(new_n565), .B2(G91), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT75), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  OR2_X1    g144(.A1(new_n527), .A2(new_n530), .ZN(G286));
  OAI221_X1 g145(.A(new_n517), .B1(new_n518), .B2(new_n519), .C1(new_n513), .C2(new_n514), .ZN(G303));
  OAI21_X1  g146(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n512), .A2(new_n516), .A3(G87), .ZN(new_n573));
  AND2_X1   g148(.A1(KEYINPUT6), .A2(G651), .ZN(new_n574));
  NOR2_X1   g149(.A1(KEYINPUT6), .A2(G651), .ZN(new_n575));
  OAI211_X1 g150(.A(G49), .B(G543), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n572), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G288));
  OAI211_X1 g157(.A(G48), .B(G543), .C1(new_n574), .C2(new_n575), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n586), .B(new_n587), .C1(new_n554), .C2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n584), .B1(new_n589), .B2(G651), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n565), .A2(G86), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G305));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT78), .B(G47), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n518), .A2(new_n593), .B1(new_n524), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n514), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G54), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n601), .A2(new_n514), .B1(new_n602), .B2(new_n524), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n565), .A2(G92), .ZN(new_n606));
  XOR2_X1   g181(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n600), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n600), .B1(new_n610), .B2(G868), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n567), .B(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n615), .B2(G868), .ZN(G280));
  XNOR2_X1  g191(.A(G280), .B(KEYINPUT81), .ZN(G297));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n610), .B1(new_n618), .B2(G860), .ZN(G148));
  INV_X1    g194(.A(new_n543), .ZN(new_n620));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n609), .A2(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n621), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G111), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n626), .A2(new_n627), .B1(new_n629), .B2(G2105), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n483), .A2(G123), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n486), .A2(new_n632), .A3(G135), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n632), .B1(new_n486), .B2(G135), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n631), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(G2100), .Z(new_n642));
  NAND3_X1  g217(.A1(new_n637), .A2(new_n638), .A3(new_n642), .ZN(G156));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(KEYINPUT84), .ZN(new_n651));
  INV_X1    g226(.A(G1341), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(KEYINPUT84), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n651), .B2(new_n653), .ZN(new_n656));
  OAI21_X1  g231(.A(G1348), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n656), .ZN(new_n658));
  INV_X1    g233(.A(G1348), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n654), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n662), .B(new_n663), .Z(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n664), .B1(new_n657), .B2(new_n660), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n644), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n667), .ZN(new_n669));
  NAND4_X1  g244(.A1(new_n669), .A2(KEYINPUT85), .A3(G14), .A4(new_n665), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G401));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT86), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n679), .A2(new_n673), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT87), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n674), .B(KEYINPUT17), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n681), .B1(new_n673), .B2(new_n682), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n678), .B(new_n683), .C1(new_n684), .C2(new_n675), .ZN(new_n685));
  XOR2_X1   g260(.A(G2096), .B(G2100), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n691), .A2(new_n692), .ZN(new_n696));
  OR3_X1    g271(.A1(new_n690), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n690), .A2(new_n696), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1991), .B(G1996), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  INV_X1    g282(.A(new_n705), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n702), .A2(new_n708), .A3(new_n703), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n707), .B1(new_n706), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(G229));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G21), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G168), .B2(new_n713), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(G1966), .ZN(new_n716));
  INV_X1    g291(.A(new_n636), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT89), .B(G29), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n713), .A2(G19), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT95), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n620), .B2(G16), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(G1341), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(G1341), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n724), .A2(new_n725), .B1(new_n715), .B2(G1966), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n713), .A2(G4), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n609), .B2(G16), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n720), .B(new_n726), .C1(new_n659), .C2(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n719), .A2(G35), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT29), .B(G2090), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n730), .B(new_n731), .C1(new_n490), .C2(new_n718), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT31), .B(G11), .ZN(new_n733));
  INV_X1    g308(.A(G28), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n734), .B2(KEYINPUT30), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  OAI22_X1  g311(.A1(new_n736), .A2(KEYINPUT101), .B1(KEYINPUT30), .B2(new_n734), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n736), .A2(KEYINPUT101), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n713), .A2(G5), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G171), .B2(new_n713), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n739), .B1(new_n741), .B2(G1961), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n732), .B(new_n742), .C1(G1961), .C2(new_n741), .ZN(new_n743));
  NAND2_X1  g318(.A1(G162), .A2(new_n719), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n731), .B1(new_n744), .B2(new_n730), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2072), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT25), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n486), .B2(G139), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n750), .A2(KEYINPUT97), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(KEYINPUT97), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  OAI22_X1  g328(.A1(new_n751), .A2(new_n752), .B1(new_n464), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G29), .ZN(new_n755));
  INV_X1    g330(.A(G29), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G33), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n747), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n729), .A2(new_n746), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G141), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n485), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT99), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT26), .Z(new_n764));
  NAND3_X1  g339(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n483), .B2(G129), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n756), .B1(new_n762), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n756), .A2(G32), .ZN(new_n769));
  OR3_X1    g344(.A1(new_n768), .A2(KEYINPUT100), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT27), .B(G1996), .ZN(new_n771));
  OAI21_X1  g346(.A(KEYINPUT100), .B1(new_n768), .B2(new_n769), .ZN(new_n772));
  AND3_X1   g347(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n713), .A2(G20), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT23), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n615), .B2(new_n713), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1956), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n718), .A2(G26), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT28), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n483), .A2(G128), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n486), .A2(G140), .ZN(new_n783));
  OR2_X1    g358(.A1(G104), .A2(G2105), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n784), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT96), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n782), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n781), .B1(new_n788), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2067), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n728), .A2(new_n659), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT24), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(G34), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(G34), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n718), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n474), .B2(new_n756), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2084), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n719), .A2(G27), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G164), .B2(new_n719), .ZN(new_n799));
  INV_X1    g374(.A(G2078), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n790), .A2(new_n791), .A3(new_n797), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n779), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n755), .A2(new_n747), .A3(new_n757), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT98), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n759), .A2(new_n775), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT34), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT93), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n713), .A2(G22), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT91), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G166), .B2(new_n713), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n810), .B1(G303), .B2(G16), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT92), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G1971), .ZN(new_n818));
  INV_X1    g393(.A(G1971), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n814), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n713), .A2(G23), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n552), .A2(new_n553), .A3(G74), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n576), .B1(new_n823), .B2(new_n514), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n512), .A2(new_n516), .A3(G87), .ZN(new_n825));
  OAI21_X1  g400(.A(KEYINPUT90), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT90), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n572), .A2(new_n573), .A3(new_n827), .A4(new_n576), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n822), .B1(new_n829), .B2(G16), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT33), .B(G1976), .Z(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n818), .A2(new_n820), .A3(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n713), .A2(G6), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G305), .B2(G16), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT32), .B(G1981), .Z(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n830), .A2(new_n832), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n808), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n818), .A2(new_n820), .A3(new_n833), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n844), .A2(new_n841), .A3(KEYINPUT93), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n807), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n834), .A2(new_n842), .A3(new_n808), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT93), .B1(new_n844), .B2(new_n841), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(KEYINPUT34), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n718), .A2(G25), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n483), .A2(G119), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n486), .A2(G131), .ZN(new_n852));
  OR2_X1    g427(.A1(G95), .A2(G2105), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n850), .B1(new_n856), .B2(new_n718), .ZN(new_n857));
  XOR2_X1   g432(.A(KEYINPUT35), .B(G1991), .Z(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n713), .A2(G24), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n598), .B2(new_n713), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G1986), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n860), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n846), .A2(new_n849), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT94), .B(KEYINPUT36), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n846), .A2(new_n849), .A3(new_n865), .A4(new_n867), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n806), .B1(new_n869), .B2(new_n870), .ZN(G311));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  INV_X1    g447(.A(new_n806), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT102), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n875));
  AOI211_X1 g450(.A(new_n875), .B(new_n806), .C1(new_n869), .C2(new_n870), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(new_n876), .ZN(G150));
  NOR2_X1   g452(.A1(new_n609), .A2(new_n618), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT38), .ZN(new_n879));
  XNOR2_X1  g454(.A(KEYINPUT103), .B(G93), .ZN(new_n880));
  INV_X1    g455(.A(G55), .ZN(new_n881));
  OAI22_X1  g456(.A1(new_n518), .A2(new_n880), .B1(new_n524), .B2(new_n881), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(new_n514), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n620), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n543), .A2(new_n885), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n879), .B(new_n889), .Z(new_n890));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n891));
  AOI21_X1  g466(.A(G860), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n886), .A2(G860), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT37), .Z(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(G145));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n636), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g473(.A(KEYINPUT104), .B(new_n631), .C1(new_n634), .C2(new_n635), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(G160), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n898), .A2(new_n474), .A3(new_n899), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n901), .A2(G162), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(G162), .B1(new_n901), .B2(new_n902), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT107), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n902), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n490), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(G162), .A3(new_n902), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n753), .A2(new_n464), .ZN(new_n911));
  INV_X1    g486(.A(new_n752), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n750), .A2(KEYINPUT97), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n788), .A2(new_n510), .ZN(new_n915));
  NAND4_X1  g490(.A1(G164), .A2(new_n782), .A3(new_n783), .A4(new_n787), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n754), .A2(new_n915), .A3(new_n916), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n762), .A2(new_n767), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n483), .A2(G130), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n486), .A2(G142), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n925));
  OR3_X1    g500(.A1(new_n925), .A2(new_n464), .A3(G118), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n464), .B2(G118), .ZN(new_n927));
  OR2_X1    g502(.A1(G106), .A2(G2105), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n926), .A2(G2104), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n923), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n640), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n930), .A2(new_n640), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n855), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n933), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(new_n856), .A3(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n921), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n918), .A2(new_n919), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n922), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n905), .B(new_n910), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n918), .A2(new_n919), .A3(new_n939), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n939), .B1(new_n918), .B2(new_n919), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n937), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n941), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n903), .A2(new_n904), .ZN(new_n951));
  AOI21_X1  g526(.A(G37), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT40), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n943), .A2(new_n948), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(new_n951), .ZN(new_n955));
  INV_X1    g530(.A(G37), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT40), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n954), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n953), .A2(new_n959), .ZN(G395));
  INV_X1    g535(.A(KEYINPUT41), .ZN(new_n961));
  NOR2_X1   g536(.A1(G299), .A2(new_n610), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n615), .A2(new_n609), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n615), .A2(new_n609), .ZN(new_n965));
  NAND2_X1  g540(.A1(G299), .A2(new_n610), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT41), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n623), .B(new_n889), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n969), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n962), .A2(new_n963), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(KEYINPUT108), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n969), .B2(new_n972), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(new_n974), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT42), .ZN(new_n978));
  XNOR2_X1  g553(.A(G290), .B(new_n829), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n829), .B(new_n598), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(G305), .B(G303), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n985), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n970), .A2(new_n974), .A3(new_n990), .A4(new_n976), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n978), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n989), .B1(new_n978), .B2(new_n991), .ZN(new_n993));
  OAI21_X1  g568(.A(G868), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n886), .A2(new_n621), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(G295));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n995), .ZN(G331));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n998));
  NAND3_X1  g573(.A1(G286), .A2(new_n998), .A3(G301), .ZN(new_n999));
  NAND2_X1  g574(.A1(G171), .A2(KEYINPUT110), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n998), .B1(new_n534), .B2(new_n536), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(G168), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n889), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n999), .A2(new_n887), .A3(new_n1002), .A4(new_n888), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(KEYINPUT111), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1003), .A2(new_n1007), .A3(new_n889), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n968), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1004), .A2(KEYINPUT112), .A3(new_n1005), .ZN(new_n1011));
  OR3_X1    g586(.A1(new_n1003), .A2(new_n889), .A3(KEYINPUT112), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n973), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(new_n989), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n956), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n968), .A2(new_n1012), .A3(new_n1011), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n973), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n989), .A2(KEYINPUT113), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n986), .A2(new_n1021), .A3(new_n988), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1017), .A2(new_n1019), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1016), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1009), .A2(new_n968), .B1(new_n1013), .B2(new_n973), .ZN(new_n1026));
  AOI21_X1  g601(.A(G37), .B1(new_n1026), .B2(new_n989), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT43), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT44), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1016), .A2(new_n1023), .A3(KEYINPUT43), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1024), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1036), .ZN(G397));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n502), .A2(G2104), .A3(new_n506), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n476), .A2(G138), .A3(new_n464), .A4(new_n497), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n476), .A2(G126), .A3(G2105), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n509), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n476), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT66), .B1(new_n1046), .B2(new_n464), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n471), .A2(G40), .A3(new_n472), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n462), .A2(new_n457), .A3(G2105), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G2067), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n788), .B(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1054), .B2(new_n939), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT46), .B1(new_n1052), .B2(G1996), .ZN(new_n1056));
  OR3_X1    g631(.A1(new_n1052), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT47), .ZN(new_n1059));
  INV_X1    g634(.A(G1996), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n939), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1054), .B1(new_n939), .B2(new_n1060), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1051), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n855), .B(new_n859), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1052), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1986), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1051), .A2(new_n1070), .A3(new_n598), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1071), .B(KEYINPUT127), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT48), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1069), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n788), .A2(G2067), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n855), .A2(new_n859), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n1064), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT126), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1052), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n1059), .B(new_n1076), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G286), .A2(G8), .ZN(new_n1084));
  NOR2_X1   g659(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n471), .A2(G40), .A3(new_n472), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n463), .A2(new_n465), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n510), .B2(new_n1038), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G2084), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1044), .A2(G1384), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n509), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1384), .B1(new_n1096), .B2(new_n507), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1088), .B(new_n1095), .C1(new_n1097), .C2(KEYINPUT45), .ZN(new_n1098));
  INV_X1    g673(.A(G1966), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1092), .A2(new_n1093), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G8), .ZN(new_n1101));
  OAI211_X1 g676(.A(KEYINPUT51), .B(new_n1084), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1043), .A2(KEYINPUT50), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1105), .A2(new_n1093), .A3(new_n1088), .A4(new_n1086), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1103), .B(G8), .C1(new_n1107), .C2(G286), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1084), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT120), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1111), .B(new_n1084), .C1(new_n1104), .C2(new_n1106), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1102), .B(new_n1108), .C1(new_n1110), .C2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT62), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1095), .A2(new_n1088), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT45), .B1(new_n510), .B2(new_n1038), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n819), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G2090), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1105), .A2(new_n1118), .A3(new_n1088), .A4(new_n1086), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G8), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT55), .B(G8), .C1(new_n515), .C2(new_n520), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n826), .A2(G1976), .A3(new_n828), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(G8), .C1(new_n1043), .C2(new_n1050), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT115), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1097), .A2(new_n1088), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1130), .A2(new_n1131), .A3(G8), .A4(new_n1127), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1132), .A3(KEYINPUT52), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT49), .ZN(new_n1134));
  INV_X1    g709(.A(G1981), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n590), .A2(new_n1135), .A3(new_n591), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(KEYINPUT116), .A2(G86), .ZN(new_n1138));
  NAND2_X1  g713(.A1(KEYINPUT116), .A2(G86), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n565), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1135), .B1(new_n590), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1134), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1141), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(KEYINPUT49), .A3(new_n1136), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1043), .A2(new_n1050), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n1101), .ZN(new_n1147));
  INV_X1    g722(.A(G1976), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT52), .B1(G288), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1128), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1145), .A2(new_n1147), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1125), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1120), .A2(G8), .A3(new_n1152), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1126), .A2(new_n1133), .A3(new_n1151), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT53), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1098), .B2(G2078), .ZN(new_n1156));
  INV_X1    g731(.A(G1961), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1050), .B1(new_n510), .B2(new_n1094), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1159), .A2(new_n1160), .A3(new_n800), .A4(new_n1045), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT53), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1160), .B1(new_n1163), .B2(new_n800), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1156), .B(new_n1158), .C1(new_n1162), .C2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(G171), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1154), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1111), .B1(new_n1100), .B2(new_n1084), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1107), .A2(KEYINPUT120), .A3(new_n1109), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1170), .A2(new_n1171), .A3(new_n1102), .A4(new_n1108), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1114), .A2(new_n1167), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1147), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1133), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n1101), .B(new_n1125), .C1(new_n1117), .C2(new_n1119), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1148), .A3(new_n581), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1136), .B(KEYINPUT117), .Z(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1177), .A2(new_n1178), .B1(new_n1181), .B2(new_n1147), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1100), .A2(new_n1101), .A3(G286), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1177), .A2(new_n1153), .A3(new_n1126), .A4(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT63), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1184), .A2(KEYINPUT118), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1185), .B1(new_n1184), .B2(KEYINPUT118), .ZN(new_n1187));
  OAI211_X1 g762(.A(new_n1173), .B(new_n1182), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(KEYINPUT56), .B(G2072), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1159), .A2(new_n1045), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(G1956), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1191), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT57), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n559), .A2(new_n566), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1193), .B1(new_n559), .B2(new_n566), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1190), .A2(new_n1192), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1197), .B1(new_n1192), .B2(new_n1190), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n659), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1146), .A2(new_n1053), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n609), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1198), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT119), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI211_X1 g780(.A(KEYINPUT119), .B(new_n1198), .C1(new_n1199), .C2(new_n1202), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1199), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1208), .A2(KEYINPUT61), .A3(new_n1198), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1198), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1210), .B1(new_n1211), .B2(new_n1199), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT60), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1200), .A2(KEYINPUT60), .A3(new_n1201), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1215), .A2(new_n610), .A3(new_n1216), .ZN(new_n1217));
  AND3_X1   g792(.A1(new_n1209), .A2(new_n1212), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1163), .A2(new_n1060), .ZN(new_n1219));
  XOR2_X1   g794(.A(KEYINPUT58), .B(G1341), .Z(new_n1220));
  NAND2_X1  g795(.A1(new_n1130), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n620), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  OAI22_X1  g797(.A1(new_n1222), .A2(KEYINPUT59), .B1(new_n610), .B2(new_n1216), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1223), .B1(KEYINPUT59), .B2(new_n1222), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1207), .B1(new_n1218), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g800(.A(new_n1152), .B1(new_n1120), .B2(G8), .ZN(new_n1226));
  NOR3_X1   g801(.A1(new_n1176), .A2(new_n1226), .A3(new_n1178), .ZN(new_n1227));
  AND2_X1   g802(.A1(new_n1113), .A2(new_n1227), .ZN(new_n1228));
  AND2_X1   g803(.A1(new_n1156), .A2(G301), .ZN(new_n1229));
  AOI211_X1 g804(.A(new_n1155), .B(G2078), .C1(new_n510), .C2(new_n1094), .ZN(new_n1230));
  OR2_X1    g805(.A1(new_n462), .A2(KEYINPUT122), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n462), .A2(KEYINPUT122), .ZN(new_n1232));
  NAND3_X1  g807(.A1(new_n1231), .A2(new_n1232), .A3(G2105), .ZN(new_n1233));
  AND3_X1   g808(.A1(new_n1233), .A2(KEYINPUT123), .A3(new_n1048), .ZN(new_n1234));
  AOI21_X1  g809(.A(KEYINPUT123), .B1(new_n1233), .B2(new_n1048), .ZN(new_n1235));
  OAI211_X1 g810(.A(new_n1230), .B(new_n1045), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1229), .A2(new_n1158), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1166), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g813(.A(KEYINPUT54), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  OAI211_X1 g815(.A(new_n1229), .B(new_n1158), .C1(new_n1164), .C2(new_n1162), .ZN(new_n1241));
  NAND3_X1  g816(.A1(new_n1156), .A2(new_n1236), .A3(new_n1158), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n1242), .A2(KEYINPUT124), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1243), .A2(G171), .ZN(new_n1244));
  NOR2_X1   g819(.A1(new_n1242), .A2(KEYINPUT124), .ZN(new_n1245));
  OAI211_X1 g820(.A(KEYINPUT54), .B(new_n1241), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g821(.A1(new_n1228), .A2(new_n1240), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g822(.A(new_n1225), .B1(new_n1247), .B2(KEYINPUT125), .ZN(new_n1248));
  INV_X1    g823(.A(KEYINPUT125), .ZN(new_n1249));
  NAND4_X1  g824(.A1(new_n1228), .A2(new_n1240), .A3(new_n1249), .A4(new_n1246), .ZN(new_n1250));
  AOI21_X1  g825(.A(new_n1188), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g826(.A(new_n598), .B(G1986), .ZN(new_n1252));
  OAI21_X1  g827(.A(new_n1069), .B1(new_n1052), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g828(.A(new_n1083), .B1(new_n1251), .B2(new_n1253), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g829(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1256));
  INV_X1    g830(.A(G319), .ZN(new_n1257));
  NOR2_X1   g831(.A1(G227), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g832(.A(new_n1258), .B1(new_n710), .B2(new_n711), .ZN(new_n1259));
  AOI21_X1  g833(.A(new_n1259), .B1(new_n668), .B2(new_n670), .ZN(new_n1260));
  OAI21_X1  g834(.A(new_n1260), .B1(new_n954), .B2(new_n957), .ZN(new_n1261));
  NOR2_X1   g835(.A1(new_n1256), .A2(new_n1261), .ZN(G308));
  OAI221_X1 g836(.A(new_n1260), .B1(new_n954), .B2(new_n957), .C1(new_n1034), .C2(new_n1035), .ZN(G225));
endmodule


