

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798;

  AND2_X1 U379 ( .A1(n636), .A2(n371), .ZN(n659) );
  XNOR2_X1 U380 ( .A(n358), .B(n357), .ZN(n394) );
  NOR2_X1 U381 ( .A1(n796), .A2(KEYINPUT44), .ZN(n358) );
  INV_X1 U382 ( .A(n564), .ZN(n357) );
  NOR2_X1 U383 ( .A1(n773), .A2(n591), .ZN(n592) );
  XNOR2_X1 U384 ( .A(n531), .B(n530), .ZN(n796) );
  NOR2_X1 U385 ( .A1(n529), .A2(n367), .ZN(n531) );
  XNOR2_X1 U386 ( .A(n590), .B(n589), .ZN(n612) );
  NOR2_X1 U387 ( .A1(n601), .A2(n547), .ZN(n476) );
  BUF_X1 U388 ( .A(n537), .Z(n359) );
  BUF_X1 U389 ( .A(n736), .Z(n360) );
  NOR2_X1 U390 ( .A1(n602), .A2(n569), .ZN(n379) );
  XNOR2_X1 U391 ( .A(n588), .B(n474), .ZN(n537) );
  XNOR2_X1 U392 ( .A(n472), .B(G469), .ZN(n588) );
  XNOR2_X1 U393 ( .A(n463), .B(n462), .ZN(n736) );
  NOR2_X1 U394 ( .A1(n678), .A2(G902), .ZN(n463) );
  NOR2_X1 U395 ( .A1(n686), .A2(G902), .ZN(n472) );
  BUF_X1 U396 ( .A(G146), .Z(n361) );
  XNOR2_X1 U397 ( .A(KEYINPUT8), .B(KEYINPUT75), .ZN(n454) );
  XNOR2_X1 U398 ( .A(KEYINPUT76), .B(KEYINPUT90), .ZN(n455) );
  XNOR2_X2 U399 ( .A(n453), .B(G953), .ZN(n479) );
  NOR2_X1 U400 ( .A1(n658), .A2(n798), .ZN(n374) );
  XNOR2_X2 U401 ( .A(n362), .B(n420), .ZN(n637) );
  NAND2_X2 U402 ( .A1(n396), .A2(n393), .ZN(n362) );
  XOR2_X2 U403 ( .A(n483), .B(n482), .Z(n366) );
  XNOR2_X1 U404 ( .A(KEYINPUT5), .B(G116), .ZN(n381) );
  XNOR2_X1 U405 ( .A(KEYINPUT80), .B(G110), .ZN(n422) );
  INV_X2 U406 ( .A(G131), .ZN(n428) );
  INV_X1 U407 ( .A(G116), .ZN(n488) );
  INV_X1 U408 ( .A(n361), .ZN(n432) );
  INV_X1 U409 ( .A(G953), .ZN(n786) );
  INV_X1 U410 ( .A(KEYINPUT64), .ZN(n453) );
  AND2_X2 U411 ( .A1(n387), .A2(n386), .ZN(n369) );
  AND2_X1 U412 ( .A1(n404), .A2(n622), .ZN(n403) );
  INV_X1 U413 ( .A(KEYINPUT45), .ZN(n420) );
  INV_X1 U414 ( .A(KEYINPUT48), .ZN(n401) );
  NAND2_X1 U415 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U416 ( .A(n402), .B(n401), .ZN(n636) );
  NAND2_X1 U417 ( .A1(n405), .A2(n403), .ZN(n402) );
  OR2_X1 U418 ( .A1(n562), .A2(n563), .ZN(n391) );
  XNOR2_X1 U419 ( .A(n374), .B(n373), .ZN(n405) );
  XNOR2_X1 U420 ( .A(n407), .B(n406), .ZN(n624) );
  XNOR2_X1 U421 ( .A(n533), .B(n532), .ZN(n759) );
  XNOR2_X1 U422 ( .A(n376), .B(KEYINPUT21), .ZN(n735) );
  XNOR2_X1 U423 ( .A(n661), .B(n432), .ZN(n471) );
  XNOR2_X1 U424 ( .A(n489), .B(n398), .ZN(n397) );
  XNOR2_X1 U425 ( .A(n464), .B(n422), .ZN(n478) );
  XNOR2_X1 U426 ( .A(n477), .B(n425), .ZN(n661) );
  XNOR2_X1 U427 ( .A(n506), .B(n426), .ZN(n425) );
  NAND2_X1 U428 ( .A1(n424), .A2(n423), .ZN(n464) );
  XNOR2_X1 U429 ( .A(n522), .B(KEYINPUT4), .ZN(n477) );
  XNOR2_X1 U430 ( .A(n377), .B(n442), .ZN(n639) );
  AND2_X1 U431 ( .A1(n563), .A2(KEYINPUT44), .ZN(n392) );
  XNOR2_X1 U432 ( .A(n488), .B(G107), .ZN(n520) );
  XNOR2_X1 U433 ( .A(n427), .B(G134), .ZN(n426) );
  INV_X1 U434 ( .A(KEYINPUT73), .ZN(n434) );
  NOR2_X1 U435 ( .A1(n637), .A2(n634), .ZN(n729) );
  BUF_X1 U436 ( .A(n567), .Z(n630) );
  NAND2_X1 U437 ( .A1(n587), .A2(n736), .ZN(n602) );
  NOR2_X1 U438 ( .A1(n735), .A2(n585), .ZN(n586) );
  INV_X1 U439 ( .A(G137), .ZN(n427) );
  INV_X1 U440 ( .A(n567), .ZN(n414) );
  OR2_X1 U441 ( .A1(n601), .A2(n382), .ZN(n626) );
  NOR2_X1 U442 ( .A1(n561), .A2(n560), .ZN(n562) );
  INV_X1 U443 ( .A(KEYINPUT15), .ZN(n442) );
  XNOR2_X1 U444 ( .A(G902), .B(KEYINPUT95), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n435), .B(n381), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U447 ( .A(G104), .B(G107), .ZN(n466) );
  NAND2_X1 U448 ( .A1(n434), .A2(G101), .ZN(n423) );
  NOR2_X1 U449 ( .A1(n617), .A2(n616), .ZN(n404) );
  NAND2_X1 U450 ( .A1(n460), .A2(G221), .ZN(n376) );
  NAND2_X1 U451 ( .A1(n414), .A2(n413), .ZN(n412) );
  NOR2_X1 U452 ( .A1(n756), .A2(KEYINPUT19), .ZN(n413) );
  XNOR2_X1 U453 ( .A(n487), .B(n486), .ZN(n505) );
  INV_X1 U454 ( .A(G104), .ZN(n486) );
  XNOR2_X1 U455 ( .A(G122), .B(G113), .ZN(n487) );
  NAND2_X1 U456 ( .A1(G234), .A2(G237), .ZN(n494) );
  XNOR2_X1 U457 ( .A(n626), .B(n603), .ZN(n604) );
  NAND2_X1 U458 ( .A1(KEYINPUT92), .A2(n390), .ZN(n389) );
  INV_X1 U459 ( .A(KEYINPUT44), .ZN(n390) );
  OR2_X1 U460 ( .A1(G237), .A2(G902), .ZN(n492) );
  INV_X1 U461 ( .A(KEYINPUT19), .ZN(n416) );
  INV_X1 U462 ( .A(G902), .ZN(n571) );
  NOR2_X1 U463 ( .A1(G953), .A2(G237), .ZN(n507) );
  NAND2_X1 U464 ( .A1(n385), .A2(n364), .ZN(n384) );
  NAND2_X1 U465 ( .A1(n411), .A2(n410), .ZN(n409) );
  INV_X1 U466 ( .A(n585), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n443), .B(n444), .ZN(n460) );
  XNOR2_X1 U468 ( .A(n380), .B(n464), .ZN(n436) );
  XNOR2_X1 U469 ( .A(G128), .B(G137), .ZN(n447) );
  XNOR2_X1 U470 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n449) );
  XNOR2_X1 U471 ( .A(G134), .B(G122), .ZN(n518) );
  XOR2_X1 U472 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n503) );
  XNOR2_X1 U473 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U474 ( .A(KEYINPUT96), .B(KEYINPUT18), .ZN(n483) );
  XOR2_X1 U475 ( .A(KEYINPUT17), .B(KEYINPUT85), .Z(n480) );
  INV_X1 U476 ( .A(n491), .ZN(n398) );
  XNOR2_X1 U477 ( .A(n379), .B(n372), .ZN(n378) );
  INV_X1 U478 ( .A(KEYINPUT39), .ZN(n406) );
  NOR2_X1 U479 ( .A1(n599), .A2(n757), .ZN(n407) );
  NOR2_X1 U480 ( .A1(n736), .A2(n735), .ZN(n732) );
  NAND2_X1 U481 ( .A1(n611), .A2(n498), .ZN(n500) );
  BUF_X1 U482 ( .A(n479), .Z(n662) );
  NOR2_X1 U483 ( .A1(n662), .A2(G952), .ZN(n698) );
  XNOR2_X1 U484 ( .A(n605), .B(KEYINPUT113), .ZN(n606) );
  AND2_X1 U485 ( .A1(n538), .A2(n608), .ZN(n539) );
  NAND2_X1 U486 ( .A1(n545), .A2(n360), .ZN(n669) );
  AND2_X1 U487 ( .A1(n414), .A2(n418), .ZN(n363) );
  AND2_X1 U488 ( .A1(n562), .A2(KEYINPUT92), .ZN(n364) );
  OR2_X1 U489 ( .A1(n418), .A2(n416), .ZN(n365) );
  NAND2_X1 U490 ( .A1(n594), .A2(n596), .ZN(n367) );
  AND2_X1 U491 ( .A1(n732), .A2(n550), .ZN(n368) );
  NAND2_X1 U492 ( .A1(G210), .A2(n492), .ZN(n370) );
  AND2_X1 U493 ( .A1(n723), .A2(n725), .ZN(n371) );
  INV_X1 U494 ( .A(n756), .ZN(n418) );
  XOR2_X1 U495 ( .A(KEYINPUT109), .B(KEYINPUT28), .Z(n372) );
  XNOR2_X1 U496 ( .A(n581), .B(n580), .ZN(n798) );
  XOR2_X1 U497 ( .A(n593), .B(KEYINPUT65), .Z(n373) );
  XOR2_X2 U498 ( .A(G146), .B(G125), .Z(n482) );
  NAND2_X1 U499 ( .A1(n391), .A2(n388), .ZN(n386) );
  OR2_X2 U500 ( .A1(n796), .A2(n565), .ZN(n431) );
  XNOR2_X1 U501 ( .A(n375), .B(n456), .ZN(n517) );
  XNOR2_X1 U502 ( .A(n455), .B(n454), .ZN(n375) );
  NAND2_X1 U503 ( .A1(n394), .A2(n566), .ZN(n393) );
  NAND2_X1 U504 ( .A1(n378), .A2(n550), .ZN(n590) );
  NAND2_X1 U505 ( .A1(n716), .A2(n383), .ZN(n382) );
  INV_X1 U506 ( .A(n602), .ZN(n383) );
  NAND2_X1 U507 ( .A1(n369), .A2(n384), .ZN(n396) );
  INV_X1 U508 ( .A(n431), .ZN(n385) );
  NAND2_X1 U509 ( .A1(n431), .A2(n392), .ZN(n387) );
  NAND2_X1 U510 ( .A1(n562), .A2(n389), .ZN(n388) );
  NAND2_X1 U511 ( .A1(n695), .A2(n639), .ZN(n419) );
  XNOR2_X2 U512 ( .A(n399), .B(n781), .ZN(n695) );
  XNOR2_X2 U513 ( .A(n397), .B(n490), .ZN(n781) );
  XNOR2_X2 U514 ( .A(n400), .B(n485), .ZN(n399) );
  XNOR2_X2 U515 ( .A(n366), .B(n484), .ZN(n400) );
  XNOR2_X2 U516 ( .A(n481), .B(n480), .ZN(n484) );
  XNOR2_X1 U517 ( .A(n471), .B(n437), .ZN(n651) );
  NAND2_X1 U518 ( .A1(n433), .A2(KEYINPUT73), .ZN(n424) );
  NAND2_X1 U519 ( .A1(n624), .A2(n716), .ZN(n581) );
  NAND2_X1 U520 ( .A1(n579), .A2(n430), .ZN(n599) );
  AND2_X1 U521 ( .A1(n550), .A2(n408), .ZN(n578) );
  NOR2_X1 U522 ( .A1(n736), .A2(n409), .ZN(n408) );
  INV_X1 U523 ( .A(n735), .ZN(n411) );
  NAND2_X2 U524 ( .A1(n415), .A2(n412), .ZN(n611) );
  AND2_X2 U525 ( .A1(n417), .A2(n365), .ZN(n415) );
  NAND2_X1 U526 ( .A1(n567), .A2(KEYINPUT19), .ZN(n417) );
  XNOR2_X2 U527 ( .A(n419), .B(n370), .ZN(n567) );
  XNOR2_X2 U528 ( .A(n428), .B(KEYINPUT78), .ZN(n506) );
  XNOR2_X2 U529 ( .A(G143), .B(G128), .ZN(n522) );
  XNOR2_X1 U530 ( .A(n478), .B(n467), .ZN(n469) );
  XOR2_X1 U531 ( .A(n491), .B(G113), .Z(n429) );
  XNOR2_X1 U532 ( .A(KEYINPUT30), .B(n570), .ZN(n430) );
  XNOR2_X1 U533 ( .A(n471), .B(n470), .ZN(n686) );
  INV_X1 U534 ( .A(G140), .ZN(n465) );
  XNOR2_X1 U535 ( .A(n436), .B(n429), .ZN(n437) );
  XNOR2_X1 U536 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U537 ( .A(n511), .B(n510), .ZN(n512) );
  INV_X1 U538 ( .A(KEYINPUT112), .ZN(n603) );
  INV_X1 U539 ( .A(n698), .ZN(n655) );
  INV_X1 U540 ( .A(G101), .ZN(n433) );
  NAND2_X1 U541 ( .A1(n507), .A2(G210), .ZN(n435) );
  XOR2_X1 U542 ( .A(KEYINPUT3), .B(G119), .Z(n491) );
  NAND2_X1 U543 ( .A1(n651), .A2(n571), .ZN(n440) );
  INV_X1 U544 ( .A(KEYINPUT100), .ZN(n438) );
  XNOR2_X1 U545 ( .A(n438), .B(G472), .ZN(n439) );
  XNOR2_X2 U546 ( .A(n440), .B(n439), .ZN(n569) );
  INV_X1 U547 ( .A(KEYINPUT6), .ZN(n441) );
  XNOR2_X1 U548 ( .A(n569), .B(n441), .ZN(n601) );
  XOR2_X1 U549 ( .A(KEYINPUT20), .B(KEYINPUT99), .Z(n444) );
  NAND2_X1 U550 ( .A1(G234), .A2(n639), .ZN(n443) );
  XOR2_X1 U551 ( .A(KEYINPUT77), .B(KEYINPUT10), .Z(n446) );
  XNOR2_X1 U552 ( .A(n482), .B(G140), .ZN(n445) );
  XNOR2_X1 U553 ( .A(n446), .B(n445), .ZN(n660) );
  XOR2_X1 U554 ( .A(G110), .B(G119), .Z(n448) );
  XNOR2_X1 U555 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U556 ( .A(KEYINPUT98), .B(KEYINPUT84), .Z(n450) );
  XNOR2_X1 U557 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U558 ( .A(n452), .B(n451), .Z(n458) );
  NAND2_X1 U559 ( .A1(n479), .A2(G234), .ZN(n456) );
  NAND2_X1 U560 ( .A1(n517), .A2(G221), .ZN(n457) );
  XNOR2_X1 U561 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U562 ( .A(n459), .B(n660), .ZN(n678) );
  AND2_X1 U563 ( .A1(n460), .A2(G217), .ZN(n461) );
  XNOR2_X1 U564 ( .A(KEYINPUT25), .B(n461), .ZN(n462) );
  AND2_X1 U565 ( .A1(n662), .A2(G227), .ZN(n468) );
  INV_X1 U566 ( .A(KEYINPUT70), .ZN(n473) );
  XNOR2_X1 U567 ( .A(n473), .B(KEYINPUT1), .ZN(n474) );
  NAND2_X1 U568 ( .A1(n732), .A2(n537), .ZN(n547) );
  XNOR2_X1 U569 ( .A(KEYINPUT33), .B(KEYINPUT81), .ZN(n475) );
  XNOR2_X1 U570 ( .A(n476), .B(n475), .ZN(n747) );
  XNOR2_X1 U571 ( .A(n478), .B(n477), .ZN(n485) );
  NAND2_X1 U572 ( .A1(n479), .A2(G224), .ZN(n481) );
  INV_X1 U573 ( .A(n505), .ZN(n490) );
  XNOR2_X1 U574 ( .A(KEYINPUT16), .B(n520), .ZN(n489) );
  NAND2_X1 U575 ( .A1(n492), .A2(G214), .ZN(n493) );
  XNOR2_X1 U576 ( .A(n493), .B(KEYINPUT97), .ZN(n756) );
  XNOR2_X1 U577 ( .A(KEYINPUT14), .B(n494), .ZN(n731) );
  INV_X1 U578 ( .A(G898), .ZN(n783) );
  AND2_X1 U579 ( .A1(n783), .A2(G902), .ZN(n495) );
  NAND2_X1 U580 ( .A1(n495), .A2(G953), .ZN(n496) );
  NAND2_X1 U581 ( .A1(n786), .A2(G952), .ZN(n574) );
  NAND2_X1 U582 ( .A1(n496), .A2(n574), .ZN(n497) );
  AND2_X1 U583 ( .A1(n731), .A2(n497), .ZN(n498) );
  INV_X1 U584 ( .A(KEYINPUT0), .ZN(n499) );
  XNOR2_X2 U585 ( .A(n500), .B(n499), .ZN(n551) );
  NAND2_X1 U586 ( .A1(n747), .A2(n551), .ZN(n501) );
  XNOR2_X1 U587 ( .A(n501), .B(KEYINPUT34), .ZN(n529) );
  XNOR2_X1 U588 ( .A(G143), .B(KEYINPUT12), .ZN(n502) );
  XNOR2_X1 U589 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U590 ( .A(n505), .B(n504), .ZN(n511) );
  XNOR2_X1 U591 ( .A(n506), .B(KEYINPUT102), .ZN(n509) );
  NAND2_X1 U592 ( .A1(G214), .A2(n507), .ZN(n508) );
  XNOR2_X1 U593 ( .A(n660), .B(n512), .ZN(n673) );
  NOR2_X1 U594 ( .A1(n673), .A2(G902), .ZN(n516) );
  XOR2_X1 U595 ( .A(KEYINPUT13), .B(KEYINPUT103), .Z(n514) );
  XNOR2_X1 U596 ( .A(KEYINPUT104), .B(G475), .ZN(n513) );
  XNOR2_X1 U597 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U598 ( .A(n516), .B(n515), .ZN(n594) );
  NAND2_X1 U599 ( .A1(n517), .A2(G217), .ZN(n526) );
  XNOR2_X1 U600 ( .A(n518), .B(KEYINPUT105), .ZN(n519) );
  XNOR2_X1 U601 ( .A(n520), .B(n519), .ZN(n524) );
  XNOR2_X1 U602 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n521) );
  XNOR2_X1 U603 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U604 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U605 ( .A(n526), .B(n525), .ZN(n682) );
  OR2_X1 U606 ( .A1(n682), .A2(G902), .ZN(n528) );
  XNOR2_X1 U607 ( .A(KEYINPUT106), .B(G478), .ZN(n527) );
  XNOR2_X1 U608 ( .A(n528), .B(n527), .ZN(n596) );
  INV_X1 U609 ( .A(KEYINPUT35), .ZN(n530) );
  OR2_X1 U610 ( .A1(n594), .A2(n596), .ZN(n533) );
  INV_X1 U611 ( .A(KEYINPUT108), .ZN(n532) );
  AND2_X1 U612 ( .A1(n759), .A2(n411), .ZN(n534) );
  NAND2_X1 U613 ( .A1(n551), .A2(n534), .ZN(n536) );
  XNOR2_X1 U614 ( .A(KEYINPUT69), .B(KEYINPUT22), .ZN(n535) );
  XNOR2_X2 U615 ( .A(n536), .B(n535), .ZN(n556) );
  AND2_X1 U616 ( .A1(n601), .A2(n360), .ZN(n538) );
  XNOR2_X1 U617 ( .A(n359), .B(KEYINPUT94), .ZN(n608) );
  NAND2_X1 U618 ( .A1(n556), .A2(n539), .ZN(n541) );
  XNOR2_X1 U619 ( .A(KEYINPUT67), .B(KEYINPUT32), .ZN(n540) );
  XNOR2_X1 U620 ( .A(n541), .B(n540), .ZN(n797) );
  INV_X1 U621 ( .A(n797), .ZN(n546) );
  INV_X1 U622 ( .A(n569), .ZN(n552) );
  NOR2_X1 U623 ( .A1(n359), .A2(n552), .ZN(n542) );
  NAND2_X1 U624 ( .A1(n556), .A2(n542), .ZN(n544) );
  INV_X1 U625 ( .A(KEYINPUT68), .ZN(n543) );
  XNOR2_X1 U626 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U627 ( .A1(n546), .A2(n669), .ZN(n565) );
  INV_X1 U628 ( .A(KEYINPUT31), .ZN(n549) );
  NOR2_X1 U629 ( .A1(n569), .A2(n547), .ZN(n743) );
  AND2_X1 U630 ( .A1(n551), .A2(n743), .ZN(n548) );
  XNOR2_X1 U631 ( .A(n549), .B(n548), .ZN(n719) );
  INV_X1 U632 ( .A(n588), .ZN(n550) );
  NAND2_X1 U633 ( .A1(n368), .A2(n551), .ZN(n553) );
  NOR2_X1 U634 ( .A1(n553), .A2(n552), .ZN(n704) );
  NOR2_X1 U635 ( .A1(n719), .A2(n704), .ZN(n555) );
  INV_X1 U636 ( .A(n596), .ZN(n554) );
  OR2_X1 U637 ( .A1(n594), .A2(n554), .ZN(n703) );
  XNOR2_X1 U638 ( .A(n703), .B(KEYINPUT107), .ZN(n623) );
  AND2_X1 U639 ( .A1(n594), .A2(n554), .ZN(n716) );
  NOR2_X1 U640 ( .A1(n623), .A2(n716), .ZN(n619) );
  NOR2_X1 U641 ( .A1(n555), .A2(n619), .ZN(n561) );
  INV_X1 U642 ( .A(n360), .ZN(n557) );
  NAND2_X1 U643 ( .A1(n601), .A2(n557), .ZN(n558) );
  NOR2_X1 U644 ( .A1(n359), .A2(n558), .ZN(n559) );
  NAND2_X1 U645 ( .A1(n556), .A2(n559), .ZN(n701) );
  INV_X1 U646 ( .A(n701), .ZN(n560) );
  INV_X1 U647 ( .A(KEYINPUT92), .ZN(n563) );
  INV_X1 U648 ( .A(KEYINPUT74), .ZN(n564) );
  INV_X1 U649 ( .A(n565), .ZN(n566) );
  INV_X1 U650 ( .A(KEYINPUT38), .ZN(n568) );
  XNOR2_X1 U651 ( .A(n630), .B(n568), .ZN(n757) );
  NOR2_X1 U652 ( .A1(n569), .A2(n756), .ZN(n570) );
  INV_X1 U653 ( .A(n662), .ZN(n573) );
  NOR2_X1 U654 ( .A1(n571), .A2(G900), .ZN(n572) );
  NAND2_X1 U655 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U656 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U657 ( .A1(n731), .A2(n576), .ZN(n585) );
  INV_X1 U658 ( .A(KEYINPUT83), .ZN(n577) );
  XNOR2_X1 U659 ( .A(n578), .B(n577), .ZN(n579) );
  INV_X1 U660 ( .A(KEYINPUT40), .ZN(n580) );
  NOR2_X1 U661 ( .A1(n757), .A2(n756), .ZN(n582) );
  NAND2_X1 U662 ( .A1(n582), .A2(n759), .ZN(n584) );
  XNOR2_X1 U663 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n583) );
  XNOR2_X1 U664 ( .A(n584), .B(n583), .ZN(n773) );
  XOR2_X1 U665 ( .A(KEYINPUT79), .B(n586), .Z(n587) );
  INV_X1 U666 ( .A(KEYINPUT110), .ZN(n589) );
  INV_X1 U667 ( .A(n612), .ZN(n591) );
  XNOR2_X1 U668 ( .A(n592), .B(KEYINPUT42), .ZN(n658) );
  XOR2_X1 U669 ( .A(KEYINPUT91), .B(KEYINPUT46), .Z(n593) );
  INV_X1 U670 ( .A(n594), .ZN(n595) );
  NOR2_X1 U671 ( .A1(n595), .A2(n630), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n713) );
  INV_X1 U674 ( .A(KEYINPUT89), .ZN(n618) );
  NOR2_X1 U675 ( .A1(KEYINPUT47), .A2(n618), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n713), .A2(n600), .ZN(n610) );
  NAND2_X1 U677 ( .A1(n604), .A2(n363), .ZN(n607) );
  XOR2_X1 U678 ( .A(KEYINPUT36), .B(KEYINPUT93), .Z(n605) );
  XNOR2_X1 U679 ( .A(n607), .B(n606), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n722) );
  NAND2_X1 U681 ( .A1(n610), .A2(n722), .ZN(n617) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT86), .ZN(n709) );
  NOR2_X1 U684 ( .A1(n619), .A2(KEYINPUT47), .ZN(n614) );
  NOR2_X1 U685 ( .A1(n614), .A2(KEYINPUT89), .ZN(n615) );
  NOR2_X1 U686 ( .A1(n709), .A2(n615), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n709), .A2(n618), .ZN(n620) );
  INV_X1 U688 ( .A(n619), .ZN(n748) );
  NAND2_X1 U689 ( .A1(n620), .A2(n748), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n621), .A2(KEYINPUT47), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n624), .A2(n623), .ZN(n723) );
  NAND2_X1 U692 ( .A1(n723), .A2(KEYINPUT2), .ZN(n625) );
  XOR2_X1 U693 ( .A(KEYINPUT87), .B(n625), .Z(n632) );
  NOR2_X1 U694 ( .A1(n359), .A2(n626), .ZN(n627) );
  NAND2_X1 U695 ( .A1(n418), .A2(n627), .ZN(n628) );
  XNOR2_X1 U696 ( .A(n628), .B(KEYINPUT43), .ZN(n629) );
  NAND2_X1 U697 ( .A1(n630), .A2(n629), .ZN(n725) );
  INV_X1 U698 ( .A(n725), .ZN(n631) );
  NOR2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U700 ( .A1(n636), .A2(n633), .ZN(n634) );
  AND2_X1 U701 ( .A1(n639), .A2(KEYINPUT72), .ZN(n635) );
  NOR2_X1 U702 ( .A1(n729), .A2(n635), .ZN(n648) );
  XNOR2_X1 U703 ( .A(n659), .B(KEYINPUT82), .ZN(n638) );
  INV_X1 U704 ( .A(n637), .ZN(n726) );
  NAND2_X1 U705 ( .A1(n638), .A2(n726), .ZN(n646) );
  INV_X1 U706 ( .A(n639), .ZN(n641) );
  INV_X1 U707 ( .A(KEYINPUT2), .ZN(n642) );
  NOR2_X1 U708 ( .A1(n642), .A2(KEYINPUT72), .ZN(n640) );
  NAND2_X1 U709 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U710 ( .A1(n642), .A2(KEYINPUT72), .ZN(n643) );
  NAND2_X1 U711 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n647) );
  INV_X1 U713 ( .A(KEYINPUT66), .ZN(n649) );
  XNOR2_X2 U714 ( .A(n650), .B(n649), .ZN(n692) );
  NAND2_X1 U715 ( .A1(n692), .A2(G472), .ZN(n653) );
  XOR2_X1 U716 ( .A(n651), .B(KEYINPUT62), .Z(n652) );
  XNOR2_X1 U717 ( .A(n653), .B(n652), .ZN(n654) );
  INV_X1 U718 ( .A(n654), .ZN(n656) );
  NAND2_X1 U719 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U720 ( .A(n657), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U721 ( .A(G137), .B(n658), .Z(G39) );
  XOR2_X1 U722 ( .A(n661), .B(n660), .Z(n664) );
  XNOR2_X1 U723 ( .A(n659), .B(n664), .ZN(n663) );
  NAND2_X1 U724 ( .A1(n663), .A2(n662), .ZN(n668) );
  XOR2_X1 U725 ( .A(G227), .B(n664), .Z(n665) );
  NAND2_X1 U726 ( .A1(n665), .A2(G900), .ZN(n666) );
  NAND2_X1 U727 ( .A1(G953), .A2(n666), .ZN(n667) );
  NAND2_X1 U728 ( .A1(n668), .A2(n667), .ZN(G72) );
  INV_X1 U729 ( .A(n669), .ZN(n670) );
  XOR2_X1 U730 ( .A(G110), .B(n670), .Z(G12) );
  NAND2_X1 U731 ( .A1(n692), .A2(G475), .ZN(n675) );
  XNOR2_X1 U732 ( .A(KEYINPUT71), .B(KEYINPUT123), .ZN(n671) );
  XOR2_X1 U733 ( .A(n671), .B(KEYINPUT59), .Z(n672) );
  XNOR2_X1 U734 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U735 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X2 U736 ( .A1(n676), .A2(n698), .ZN(n677) );
  XNOR2_X1 U737 ( .A(n677), .B(KEYINPUT60), .ZN(G60) );
  BUF_X1 U738 ( .A(n692), .Z(n685) );
  NAND2_X1 U739 ( .A1(n685), .A2(G217), .ZN(n680) );
  XNOR2_X1 U740 ( .A(n678), .B(KEYINPUT124), .ZN(n679) );
  XNOR2_X1 U741 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n681), .A2(n698), .ZN(G66) );
  NAND2_X1 U743 ( .A1(n685), .A2(G478), .ZN(n683) );
  XNOR2_X1 U744 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U745 ( .A1(n684), .A2(n698), .ZN(G63) );
  NAND2_X1 U746 ( .A1(n685), .A2(G469), .ZN(n690) );
  XOR2_X1 U747 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n688) );
  XNOR2_X1 U748 ( .A(n686), .B(KEYINPUT122), .ZN(n687) );
  XNOR2_X1 U749 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U750 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U751 ( .A1(n691), .A2(n698), .ZN(G54) );
  NAND2_X1 U752 ( .A1(n692), .A2(G210), .ZN(n697) );
  XNOR2_X1 U753 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n693) );
  XOR2_X1 U754 ( .A(n693), .B(KEYINPUT55), .Z(n694) );
  XNOR2_X1 U755 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U756 ( .A(n697), .B(n696), .ZN(n699) );
  NOR2_X2 U757 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U758 ( .A(n700), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U759 ( .A(n701), .B(G101), .ZN(G3) );
  NAND2_X1 U760 ( .A1(n704), .A2(n716), .ZN(n702) );
  XNOR2_X1 U761 ( .A(n702), .B(G104), .ZN(G6) );
  XNOR2_X1 U762 ( .A(G107), .B(KEYINPUT27), .ZN(n708) );
  XOR2_X1 U763 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n706) );
  INV_X1 U764 ( .A(n703), .ZN(n718) );
  NAND2_X1 U765 ( .A1(n704), .A2(n718), .ZN(n705) );
  XNOR2_X1 U766 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U767 ( .A(n708), .B(n707), .ZN(G9) );
  XOR2_X1 U768 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n711) );
  INV_X1 U769 ( .A(n709), .ZN(n714) );
  NAND2_X1 U770 ( .A1(n714), .A2(n718), .ZN(n710) );
  XNOR2_X1 U771 ( .A(n711), .B(n710), .ZN(n712) );
  XOR2_X1 U772 ( .A(G128), .B(n712), .Z(G30) );
  XOR2_X1 U773 ( .A(G143), .B(n713), .Z(G45) );
  NAND2_X1 U774 ( .A1(n714), .A2(n716), .ZN(n715) );
  XNOR2_X1 U775 ( .A(n715), .B(n361), .ZN(G48) );
  NAND2_X1 U776 ( .A1(n719), .A2(n716), .ZN(n717) );
  XNOR2_X1 U777 ( .A(n717), .B(G113), .ZN(G15) );
  NAND2_X1 U778 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U779 ( .A(n720), .B(G116), .ZN(G18) );
  XOR2_X1 U780 ( .A(G125), .B(KEYINPUT37), .Z(n721) );
  XNOR2_X1 U781 ( .A(n722), .B(n721), .ZN(G27) );
  INV_X1 U782 ( .A(n723), .ZN(n724) );
  XOR2_X1 U783 ( .A(G134), .B(n724), .Z(G36) );
  XNOR2_X1 U784 ( .A(G140), .B(n725), .ZN(G42) );
  NAND2_X1 U785 ( .A1(n726), .A2(n659), .ZN(n728) );
  XOR2_X1 U786 ( .A(KEYINPUT2), .B(KEYINPUT88), .Z(n727) );
  AND2_X1 U787 ( .A1(n728), .A2(n727), .ZN(n730) );
  NOR2_X1 U788 ( .A1(n730), .A2(n729), .ZN(n779) );
  INV_X1 U789 ( .A(n731), .ZN(n770) );
  OR2_X1 U790 ( .A1(n732), .A2(n359), .ZN(n733) );
  XNOR2_X1 U791 ( .A(KEYINPUT50), .B(n733), .ZN(n734) );
  NAND2_X1 U792 ( .A1(n734), .A2(n569), .ZN(n741) );
  XOR2_X1 U793 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n738) );
  NAND2_X1 U794 ( .A1(n360), .A2(n735), .ZN(n737) );
  XNOR2_X1 U795 ( .A(n738), .B(n737), .ZN(n739) );
  XNOR2_X1 U796 ( .A(n739), .B(KEYINPUT116), .ZN(n740) );
  NOR2_X1 U797 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U798 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U799 ( .A(KEYINPUT51), .B(n744), .Z(n745) );
  XNOR2_X1 U800 ( .A(n745), .B(KEYINPUT118), .ZN(n746) );
  NOR2_X1 U801 ( .A1(n746), .A2(n773), .ZN(n767) );
  BUF_X1 U802 ( .A(n747), .Z(n772) );
  NAND2_X1 U803 ( .A1(n748), .A2(n418), .ZN(n755) );
  INV_X1 U804 ( .A(n755), .ZN(n749) );
  NAND2_X1 U805 ( .A1(n749), .A2(KEYINPUT119), .ZN(n753) );
  INV_X1 U806 ( .A(n759), .ZN(n751) );
  INV_X1 U807 ( .A(n757), .ZN(n750) );
  NAND2_X1 U808 ( .A1(n751), .A2(n750), .ZN(n752) );
  OR2_X1 U809 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U810 ( .A1(n772), .A2(n754), .ZN(n764) );
  OR2_X1 U811 ( .A1(n755), .A2(n757), .ZN(n761) );
  NAND2_X1 U812 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U813 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U814 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U815 ( .A1(KEYINPUT119), .A2(n762), .ZN(n763) );
  NOR2_X1 U816 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U817 ( .A(n765), .B(KEYINPUT120), .ZN(n766) );
  NOR2_X1 U818 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U819 ( .A(n768), .B(KEYINPUT52), .ZN(n769) );
  NOR2_X1 U820 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U821 ( .A1(n771), .A2(G952), .ZN(n777) );
  INV_X1 U822 ( .A(n772), .ZN(n774) );
  NOR2_X1 U823 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U824 ( .A1(n775), .A2(G953), .ZN(n776) );
  NAND2_X1 U825 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U826 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U827 ( .A(n780), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U828 ( .A(G101), .B(n781), .Z(n782) );
  XNOR2_X1 U829 ( .A(G110), .B(n782), .ZN(n785) );
  AND2_X1 U830 ( .A1(n783), .A2(G953), .ZN(n784) );
  NOR2_X1 U831 ( .A1(n785), .A2(n784), .ZN(n795) );
  NAND2_X1 U832 ( .A1(n726), .A2(n786), .ZN(n792) );
  XOR2_X1 U833 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n788) );
  NAND2_X1 U834 ( .A1(G224), .A2(G953), .ZN(n787) );
  XNOR2_X1 U835 ( .A(n788), .B(n787), .ZN(n789) );
  NAND2_X1 U836 ( .A1(G898), .A2(n789), .ZN(n790) );
  XNOR2_X1 U837 ( .A(n790), .B(KEYINPUT126), .ZN(n791) );
  NAND2_X1 U838 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U839 ( .A(n793), .B(KEYINPUT127), .Z(n794) );
  XNOR2_X1 U840 ( .A(n795), .B(n794), .ZN(G69) );
  XOR2_X1 U841 ( .A(n796), .B(G122), .Z(G24) );
  XOR2_X1 U842 ( .A(G119), .B(n797), .Z(G21) );
  XOR2_X1 U843 ( .A(G131), .B(n798), .Z(G33) );
endmodule

