//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1239, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND3_X1  g0014(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(G58), .A2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G50), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n204), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n214), .B1(new_n215), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n227), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G13), .ZN(new_n248));
  NOR3_X1   g0048(.A1(new_n248), .A2(new_n209), .A3(G1), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n220), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT12), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n208), .A2(G20), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(G68), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT66), .B1(new_n258), .B2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT66), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(new_n209), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G50), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n267), .A2(new_n268), .B1(new_n209), .B2(G68), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n254), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT11), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n251), .B(new_n257), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G1), .A3(G13), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n280), .A3(G274), .ZN(new_n281));
  INV_X1    g0081(.A(new_n278), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n280), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n281), .B1(new_n283), .B2(new_n221), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT70), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT65), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT65), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G1698), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n286), .A2(new_n288), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G226), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n285), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n286), .A2(new_n288), .A3(G232), .A4(G1698), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G97), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT3), .B(G33), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT65), .B(G1698), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n299), .A2(new_n300), .A3(KEYINPUT70), .A4(G226), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n295), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n280), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n284), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g0104(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT72), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n305), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n296), .A2(new_n297), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n299), .A2(new_n300), .A3(G226), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n308), .B1(new_n285), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n280), .B1(new_n310), .B2(new_n301), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n307), .B1(new_n311), .B2(new_n284), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n302), .A2(new_n303), .ZN(new_n314));
  INV_X1    g0114(.A(new_n284), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(KEYINPUT72), .A3(new_n307), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n313), .A2(G169), .A3(new_n317), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n318), .A2(KEYINPUT14), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT14), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n313), .A2(new_n320), .A3(G169), .A4(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n304), .A2(new_n305), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT13), .B1(new_n316), .B2(KEYINPUT73), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT73), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n304), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g0125(.A(G179), .B(new_n322), .C1(new_n323), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n275), .B1(new_n319), .B2(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(G190), .B(new_n322), .C1(new_n323), .C2(new_n325), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n313), .A2(G200), .A3(new_n317), .ZN(new_n330));
  AND3_X1   g0130(.A1(new_n329), .A2(new_n330), .A3(new_n274), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n255), .A2(G77), .A3(new_n256), .ZN(new_n334));
  INV_X1    g0134(.A(new_n254), .ZN(new_n335));
  XOR2_X1   g0135(.A(KEYINPUT8), .B(G58), .Z(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(new_n266), .B1(G20), .B2(G77), .ZN(new_n337));
  XOR2_X1   g0137(.A(KEYINPUT15), .B(G87), .Z(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n262), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n335), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  AOI211_X1 g0140(.A(new_n334), .B(new_n340), .C1(new_n264), .C2(new_n249), .ZN(new_n341));
  INV_X1    g0141(.A(G244), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n281), .B1(new_n342), .B2(new_n283), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n343), .A2(KEYINPUT69), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n299), .A2(G238), .A3(G1698), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n205), .B2(new_n299), .ZN(new_n346));
  INV_X1    g0146(.A(new_n299), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n290), .A2(new_n292), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n347), .A2(new_n348), .A3(new_n227), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n303), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n343), .A2(KEYINPUT69), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n344), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G169), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n341), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n352), .ZN(new_n355));
  INV_X1    g0155(.A(G179), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n352), .A2(G200), .ZN(new_n360));
  INV_X1    g0160(.A(G190), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n360), .B(new_n341), .C1(new_n361), .C2(new_n352), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n299), .A2(G223), .A3(G1698), .ZN(new_n365));
  INV_X1    g0165(.A(G222), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n365), .B1(new_n264), .B2(new_n299), .C1(new_n366), .C2(new_n293), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n367), .A2(new_n303), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n281), .B1(new_n283), .B2(new_n294), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n256), .A2(G50), .ZN(new_n371));
  XOR2_X1   g0171(.A(new_n371), .B(KEYINPUT67), .Z(new_n372));
  INV_X1    g0172(.A(new_n255), .ZN(new_n373));
  INV_X1    g0173(.A(new_n249), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n372), .A2(new_n373), .B1(G50), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n202), .A2(G20), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n336), .A2(new_n262), .B1(G150), .B2(new_n266), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n335), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n370), .A2(G190), .B1(new_n379), .B2(KEYINPUT9), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G200), .ZN(new_n382));
  OAI22_X1  g0182(.A1(new_n370), .A2(new_n382), .B1(new_n379), .B2(KEYINPUT9), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT10), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n383), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT10), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n386), .A3(new_n380), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n364), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n370), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(G179), .ZN(new_n391));
  INV_X1    g0191(.A(new_n379), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n370), .B2(G169), .ZN(new_n393));
  OR3_X1    g0193(.A1(new_n391), .A2(new_n393), .A3(KEYINPUT68), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT68), .B1(new_n391), .B2(new_n393), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n226), .A2(new_n220), .ZN(new_n399));
  OAI21_X1  g0199(.A(G20), .B1(new_n399), .B2(new_n216), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n266), .A2(G159), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n287), .A2(KEYINPUT74), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT74), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT3), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n405), .A3(G33), .ZN(new_n406));
  AOI21_X1  g0206(.A(G20), .B1(new_n406), .B2(new_n286), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT7), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n220), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n286), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n411), .B2(G33), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT7), .B1(new_n412), .B2(G20), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n402), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT16), .ZN(new_n415));
  XOR2_X1   g0215(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n416));
  NOR2_X1   g0216(.A1(new_n408), .A2(G20), .ZN(new_n417));
  AOI21_X1  g0217(.A(G33), .B1(new_n403), .B2(new_n405), .ZN(new_n418));
  INV_X1    g0218(.A(new_n288), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n408), .B1(new_n299), .B2(G20), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n220), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n416), .B1(new_n422), .B2(new_n402), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n415), .A2(new_n254), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n336), .A2(new_n256), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n373), .A2(new_n425), .B1(new_n374), .B2(new_n336), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n290), .A2(new_n292), .A3(G223), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G226), .A2(G1698), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n412), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G87), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n280), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n281), .B1(new_n283), .B2(new_n227), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n428), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n435), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n412), .A2(new_n431), .B1(G33), .B2(G87), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n437), .B(KEYINPUT76), .C1(new_n280), .C2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(G200), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n434), .A2(G190), .A3(new_n435), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n424), .B(new_n427), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT77), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n398), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n436), .A2(new_n439), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n353), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n437), .B(new_n356), .C1(new_n280), .C2(new_n438), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n335), .B1(new_n414), .B2(KEYINPUT16), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n426), .B1(new_n449), .B2(new_n423), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT18), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n445), .A2(new_n382), .ZN(new_n452));
  INV_X1    g0252(.A(new_n441), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n454), .A2(KEYINPUT77), .A3(KEYINPUT17), .A4(new_n450), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n424), .A2(new_n427), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n456), .A2(new_n457), .A3(new_n446), .A4(new_n447), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n444), .A2(new_n451), .A3(new_n455), .A4(new_n458), .ZN(new_n459));
  NOR4_X1   g0259(.A1(new_n333), .A2(new_n389), .A3(new_n397), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT4), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(new_n342), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n299), .A2(new_n300), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n299), .A2(G250), .A3(G1698), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n406), .A2(G244), .A3(new_n286), .A4(new_n300), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n461), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n280), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT78), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT5), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(G41), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n276), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n277), .A2(G1), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(G41), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n280), .A2(G274), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n208), .B(G45), .C1(new_n276), .C2(KEYINPUT5), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n471), .A2(G41), .ZN(new_n480));
  OAI211_X1 g0280(.A(G257), .B(new_n280), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n353), .B1(new_n469), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n482), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n485), .B1(new_n461), .B2(new_n467), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n484), .B(new_n356), .C1(new_n486), .C2(new_n280), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n205), .B1(new_n420), .B2(new_n421), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT6), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n489), .A2(new_n204), .A3(G107), .ZN(new_n490));
  XNOR2_X1  g0290(.A(G97), .B(G107), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n492), .A2(new_n209), .B1(new_n264), .B2(new_n267), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n254), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n208), .A2(G33), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n255), .A2(new_n495), .ZN(new_n496));
  MUX2_X1   g0296(.A(new_n374), .B(new_n496), .S(G97), .Z(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n483), .A2(new_n487), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT79), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT79), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n483), .A2(new_n487), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n466), .A2(new_n468), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n482), .B1(new_n503), .B2(new_n303), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G190), .ZN(new_n505));
  OAI21_X1  g0305(.A(G200), .B1(new_n469), .B2(new_n482), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n494), .A3(new_n497), .A4(new_n506), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n500), .A2(new_n502), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n406), .A2(new_n286), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n300), .A2(G238), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT80), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G116), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n258), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n406), .A2(G244), .A3(G1698), .A4(new_n286), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n290), .A2(new_n292), .A3(G238), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT80), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n286), .A4(new_n406), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n511), .A2(new_n514), .A3(new_n515), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n303), .ZN(new_n520));
  OR3_X1    g0320(.A1(new_n277), .A2(G1), .A3(G274), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n223), .B1(new_n277), .B2(G1), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n521), .A2(new_n280), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT81), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n523), .B1(new_n519), .B2(new_n303), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT81), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n356), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n374), .A2(new_n338), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n263), .B2(new_n204), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n412), .A2(new_n209), .A3(G68), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n209), .B1(new_n297), .B2(new_n532), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT82), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(KEYINPUT82), .B(new_n209), .C1(new_n297), .C2(new_n532), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n538), .C1(G87), .C2(new_n206), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n533), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT83), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n335), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT83), .A4(new_n539), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n531), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n338), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(new_n496), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n528), .B1(new_n520), .B2(new_n524), .ZN(new_n547));
  AOI211_X1 g0347(.A(KEYINPUT81), .B(new_n523), .C1(new_n519), .C2(new_n303), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n353), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n530), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n526), .A2(G190), .A3(new_n529), .ZN(new_n551));
  OAI21_X1  g0351(.A(G200), .B1(new_n547), .B2(new_n548), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n496), .A2(new_n222), .ZN(new_n553));
  AOI211_X1 g0353(.A(new_n531), .B(new_n553), .C1(new_n542), .C2(new_n543), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n508), .A2(new_n550), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n255), .A2(G116), .A3(new_n495), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n249), .A2(new_n512), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n252), .A2(new_n253), .B1(G20), .B2(new_n512), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n465), .B(new_n209), .C1(G33), .C2(new_n204), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n559), .A2(KEYINPUT20), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT20), .B1(new_n559), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n557), .B(new_n558), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G264), .A2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n348), .B2(new_n228), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n412), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n347), .A2(G303), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n280), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n280), .B1(new_n479), .B2(new_n480), .ZN(new_n569));
  INV_X1    g0369(.A(G270), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n569), .A2(new_n570), .B1(new_n476), .B2(new_n477), .ZN(new_n571));
  OAI211_X1 g0371(.A(G169), .B(new_n563), .C1(new_n568), .C2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n571), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n565), .A2(new_n412), .B1(G303), .B2(new_n347), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n575), .B1(new_n576), .B2(new_n280), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n577), .A2(KEYINPUT21), .A3(G169), .A4(new_n563), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n568), .A2(new_n571), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(G179), .A3(new_n563), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n574), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n563), .B1(new_n577), .B2(G200), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n582), .A2(KEYINPUT84), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n582), .A2(KEYINPUT84), .B1(G190), .B2(new_n579), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT86), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n290), .A2(new_n292), .A3(G250), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G257), .A2(G1698), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n412), .A2(new_n589), .B1(G33), .B2(G294), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n586), .B1(new_n590), .B2(new_n280), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G294), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n300), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n593), .B2(new_n509), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(KEYINPUT86), .A3(new_n303), .ZN(new_n595));
  OAI211_X1 g0395(.A(G264), .B(new_n280), .C1(new_n479), .C2(new_n480), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n477), .B2(new_n476), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n591), .A2(new_n595), .A3(new_n361), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT88), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n412), .A2(new_n589), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n280), .B1(new_n601), .B2(new_n592), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n597), .B1(new_n602), .B2(KEYINPUT86), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT88), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n361), .A4(new_n591), .ZN(new_n605));
  INV_X1    g0405(.A(new_n478), .ZN(new_n606));
  INV_X1    g0406(.A(new_n596), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT87), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n594), .A2(new_n303), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT87), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n596), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n606), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n600), .B(new_n605), .C1(new_n612), .C2(G200), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n249), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT25), .B1(new_n249), .B2(new_n205), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n496), .A2(new_n205), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT22), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n209), .A2(G87), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n618), .B1(new_n347), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT23), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n209), .B2(G107), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n622), .A2(new_n623), .B1(new_n513), .B2(new_n209), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n412), .A2(new_n209), .ZN(new_n625));
  NAND2_X1  g0425(.A1(KEYINPUT22), .A2(G87), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n620), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g0427(.A(KEYINPUT85), .B(KEYINPUT24), .Z(new_n628));
  XNOR2_X1  g0428(.A(new_n627), .B(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n617), .B1(new_n629), .B2(new_n254), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n613), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n617), .ZN(new_n632));
  INV_X1    g0432(.A(new_n628), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n627), .B(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n634), .B2(new_n335), .ZN(new_n635));
  AOI211_X1 g0435(.A(new_n356), .B(new_n606), .C1(new_n608), .C2(new_n611), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n353), .B1(new_n603), .B2(new_n591), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n585), .A2(new_n631), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n556), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n460), .A2(new_n640), .ZN(G372));
  NAND2_X1  g0441(.A1(new_n500), .A2(new_n502), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n550), .A2(new_n555), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT26), .ZN(new_n644));
  INV_X1    g0444(.A(new_n581), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n637), .B1(G179), .B2(new_n612), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(new_n630), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n525), .A2(KEYINPUT89), .A3(G200), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n527), .B2(new_n382), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n551), .A2(new_n651), .A3(new_n554), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n508), .A2(new_n647), .A3(new_n631), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n525), .A2(new_n353), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n530), .A2(new_n546), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  INV_X1    g0456(.A(new_n499), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n652), .A2(new_n655), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n644), .A2(new_n653), .A3(new_n655), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n460), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n451), .A2(new_n458), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n318), .A2(KEYINPUT14), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n326), .A3(new_n321), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n332), .A2(new_n359), .B1(new_n663), .B2(new_n275), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n444), .A2(new_n455), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n397), .B1(new_n666), .B2(new_n388), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n660), .A2(new_n667), .ZN(G369));
  NAND3_X1  g0468(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n563), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n585), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n645), .B2(new_n675), .ZN(new_n677));
  XOR2_X1   g0477(.A(KEYINPUT90), .B(G330), .Z(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n631), .A2(new_n638), .ZN(new_n681));
  INV_X1    g0481(.A(new_n674), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n681), .B1(new_n630), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n638), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n674), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n645), .A2(new_n674), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n681), .A2(new_n688), .B1(new_n684), .B2(new_n682), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT91), .ZN(G399));
  NAND2_X1  g0491(.A1(new_n212), .A2(new_n276), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT92), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n218), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT31), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n575), .B(G179), .C1(new_n280), .C2(new_n576), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n608), .B2(new_n611), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n526), .A2(new_n701), .A3(new_n504), .A4(new_n529), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n547), .A2(new_n548), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(KEYINPUT30), .A3(new_n504), .A4(new_n701), .ZN(new_n706));
  NOR4_X1   g0506(.A1(new_n527), .A2(new_n504), .A3(new_n579), .A4(G179), .ZN(new_n707));
  INV_X1    g0507(.A(new_n612), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n704), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n674), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n640), .A2(new_n682), .B1(new_n699), .B2(new_n711), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n702), .A2(new_n703), .B1(new_n707), .B2(new_n708), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT93), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n706), .B1(new_n713), .B2(new_n714), .ZN(new_n716));
  OAI211_X1 g0516(.A(KEYINPUT31), .B(new_n674), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n678), .B1(new_n712), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n659), .A2(new_n682), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n652), .A2(new_n655), .A3(new_n657), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT26), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n550), .A2(new_n555), .A3(new_n656), .A4(new_n642), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n653), .A3(new_n655), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n721), .B1(new_n725), .B2(new_n682), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n718), .A2(new_n720), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n698), .B1(new_n727), .B2(G1), .ZN(G364));
  NOR2_X1   g0528(.A1(new_n248), .A2(G20), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n208), .B1(new_n729), .B2(G45), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n694), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n680), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n679), .B2(new_n677), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n212), .A2(new_n299), .ZN(new_n735));
  INV_X1    g0535(.A(G355), .ZN(new_n736));
  OAI22_X1  g0536(.A1(new_n735), .A2(new_n736), .B1(G116), .B2(new_n212), .ZN(new_n737));
  INV_X1    g0537(.A(new_n212), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n412), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n218), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n740), .B1(new_n277), .B2(new_n741), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n246), .A2(new_n277), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n737), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n248), .A2(new_n258), .A3(KEYINPUT94), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT94), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G13), .B2(G33), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n253), .B1(G20), .B2(new_n353), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n732), .B1(new_n744), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n361), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n356), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G190), .A2(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n209), .A2(new_n356), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n760), .A2(KEYINPUT95), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(KEYINPUT95), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n299), .B1(new_n758), .B2(new_n204), .C1(new_n763), .C2(new_n264), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n755), .B1(new_n761), .B2(new_n762), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n764), .B1(G58), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n209), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n759), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT96), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(KEYINPUT32), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n772), .A2(KEYINPUT32), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n760), .A2(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n361), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n768), .A2(new_n361), .A3(G200), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n777), .A2(new_n268), .B1(new_n778), .B2(new_n205), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n775), .A2(G190), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n220), .B1(new_n782), .B2(new_n222), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n767), .A2(new_n773), .A3(new_n774), .A4(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n776), .A2(G326), .B1(new_n757), .B2(G294), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n787), .B2(new_n763), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT97), .Z(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n781), .A2(new_n790), .B1(new_n778), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n769), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n299), .B1(new_n793), .B2(G329), .ZN(new_n794));
  INV_X1    g0594(.A(G303), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n795), .B2(new_n782), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G322), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n798), .B2(new_n765), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n785), .B1(new_n789), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n754), .B1(new_n800), .B2(new_n751), .ZN(new_n801));
  INV_X1    g0601(.A(new_n750), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n677), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n734), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NAND2_X1  g0605(.A1(new_n359), .A2(new_n682), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n341), .A2(new_n682), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n358), .B1(new_n363), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n719), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n809), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n659), .A2(new_n682), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n718), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n732), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n718), .A2(new_n810), .A3(new_n812), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n748), .A2(new_n751), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n731), .B1(new_n264), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n751), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n347), .B1(new_n769), .B2(new_n787), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(G97), .B2(new_n757), .ZN(new_n821));
  INV_X1    g0621(.A(G294), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n512), .B2(new_n763), .C1(new_n822), .C2(new_n765), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n222), .A2(new_n778), .B1(new_n782), .B2(new_n205), .ZN(new_n824));
  XNOR2_X1  g0624(.A(KEYINPUT98), .B(G283), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n795), .A2(new_n777), .B1(new_n781), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n823), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n780), .A2(G150), .B1(new_n776), .B2(G137), .ZN(new_n828));
  INV_X1    g0628(.A(G143), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n829), .B2(new_n765), .C1(new_n770), .C2(new_n763), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT34), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n412), .B1(new_n833), .B2(new_n769), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n778), .A2(new_n220), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G58), .B2(new_n757), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n268), .B2(new_n782), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n832), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n830), .A2(new_n831), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n827), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n818), .B1(new_n819), .B2(new_n840), .C1(new_n811), .C2(new_n749), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n816), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G384));
  INV_X1    g0643(.A(new_n492), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n512), .B(new_n215), .C1(new_n844), .C2(KEYINPUT35), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(KEYINPUT35), .B2(new_n844), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT36), .ZN(new_n847));
  OAI21_X1  g0647(.A(G77), .B1(new_n226), .B2(new_n220), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n218), .A2(new_n848), .B1(G50), .B2(new_n220), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n849), .A2(G1), .A3(new_n248), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT99), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n274), .A2(new_n682), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n328), .A2(new_n332), .A3(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n275), .B(new_n674), .C1(new_n663), .C2(new_n331), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n809), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n585), .A2(new_n631), .A3(new_n638), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n550), .A2(new_n555), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(new_n508), .A4(new_n682), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n711), .A2(new_n699), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT103), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT100), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n416), .B1(new_n414), .B2(new_n869), .ZN(new_n870));
  AOI211_X1 g0670(.A(KEYINPUT100), .B(new_n402), .C1(new_n409), .C2(new_n413), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n449), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n427), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT101), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n872), .A2(KEYINPUT101), .A3(new_n427), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n448), .A2(new_n672), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n868), .B1(new_n878), .B2(new_n442), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n456), .A2(new_n446), .A3(new_n447), .ZN(new_n880));
  INV_X1    g0680(.A(new_n672), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n456), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n880), .A2(new_n882), .A3(new_n868), .A4(new_n442), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n872), .A2(KEYINPUT101), .A3(new_n427), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT101), .B1(new_n872), .B2(new_n427), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n886), .A2(new_n887), .A3(new_n672), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n459), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n867), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n889), .B(KEYINPUT38), .C1(new_n879), .C2(new_n884), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n857), .A2(new_n863), .A3(KEYINPUT103), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n866), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n864), .ZN(new_n898));
  INV_X1    g0698(.A(new_n882), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n459), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n880), .A2(new_n442), .A3(new_n882), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n883), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n867), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n896), .B1(new_n905), .B2(new_n892), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n898), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n897), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n460), .A2(new_n863), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n679), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n905), .A2(new_n913), .A3(new_n892), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT102), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n881), .B1(new_n446), .B2(new_n447), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n886), .A2(new_n887), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n442), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT37), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n883), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n920), .B2(new_n889), .ZN(new_n921));
  INV_X1    g0721(.A(new_n892), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT39), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT102), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n905), .A2(new_n924), .A3(new_n892), .A4(new_n913), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n915), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n328), .A2(new_n674), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n855), .A2(new_n856), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n812), .A2(new_n806), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n893), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n661), .A2(new_n881), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n460), .B1(new_n720), .B2(new_n726), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n667), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n933), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n912), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n208), .B2(new_n729), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n912), .A2(new_n936), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n852), .B1(new_n938), .B2(new_n939), .ZN(G367));
  OR3_X1    g0740(.A1(new_n655), .A2(new_n554), .A3(new_n682), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n652), .B(new_n655), .C1(new_n554), .C2(new_n682), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n498), .A2(new_n674), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n508), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n657), .A2(new_n674), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n681), .A2(new_n688), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT42), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n500), .B(new_n502), .C1(new_n949), .C2(new_n638), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n682), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n953), .A2(KEYINPUT104), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(KEYINPUT42), .B2(new_n952), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT104), .B1(new_n955), .B2(new_n953), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n944), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n960), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n962), .B(new_n944), .C1(new_n957), .C2(new_n958), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n687), .A2(new_n949), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n961), .A2(new_n965), .A3(new_n963), .ZN(new_n968));
  INV_X1    g0768(.A(new_n730), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n694), .B(KEYINPUT41), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n689), .A2(new_n948), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(KEYINPUT105), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT105), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n689), .A2(new_n973), .A3(new_n948), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n689), .A2(new_n948), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT44), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n972), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n680), .A3(new_n686), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n977), .A2(new_n979), .A3(new_n687), .A4(new_n980), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n950), .B1(new_n686), .B2(new_n688), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n680), .A2(KEYINPUT106), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n984), .B(new_n985), .Z(new_n986));
  NAND4_X1  g0786(.A1(new_n982), .A2(new_n727), .A3(new_n983), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n970), .B1(new_n987), .B2(new_n727), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n967), .B(new_n968), .C1(new_n969), .C2(new_n988), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n752), .B1(new_n212), .B2(new_n545), .C1(new_n740), .C2(new_n239), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n732), .A2(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n781), .A2(new_n822), .B1(new_n758), .B2(new_n205), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT46), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n782), .B2(new_n512), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n763), .B2(new_n825), .C1(new_n795), .C2(new_n765), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n992), .B(new_n995), .C1(G311), .C2(new_n776), .ZN(new_n996));
  INV_X1    g0796(.A(new_n782), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(KEYINPUT46), .A3(G116), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT107), .ZN(new_n999));
  INV_X1    g0799(.A(G317), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n509), .B1(new_n204), .B2(new_n778), .C1(new_n1000), .C2(new_n769), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT108), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n996), .A2(new_n999), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT109), .Z(new_n1006));
  NOR2_X1   g0806(.A1(new_n758), .A2(new_n220), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n781), .A2(new_n770), .B1(new_n777), .B2(new_n829), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n778), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1007), .B(new_n1008), .C1(G77), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(G137), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n299), .B1(new_n769), .B2(new_n1011), .C1(new_n226), .C2(new_n782), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n763), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1012), .B1(new_n1013), .B2(G50), .ZN(new_n1014));
  INV_X1    g0814(.A(G150), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1010), .B(new_n1014), .C1(new_n1015), .C2(new_n765), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1006), .A2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT47), .Z(new_n1018));
  OAI221_X1 g0818(.A(new_n991), .B1(new_n802), .B2(new_n943), .C1(new_n1018), .C2(new_n819), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n989), .A2(new_n1019), .ZN(G387));
  XOR2_X1   g0820(.A(new_n694), .B(KEYINPUT111), .Z(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n986), .B2(new_n727), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n727), .B2(new_n986), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n683), .A2(new_n685), .A3(new_n750), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n735), .A2(new_n695), .B1(G107), .B2(new_n212), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n236), .A2(new_n277), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n336), .A2(new_n268), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT50), .Z(new_n1029));
  INV_X1    g0829(.A(new_n695), .ZN(new_n1030));
  AOI211_X1 g0830(.A(G45), .B(new_n1030), .C1(G68), .C2(G77), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n740), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1026), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n732), .B1(new_n1033), .B2(new_n753), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n782), .A2(new_n264), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n412), .B1(new_n1015), .B2(new_n769), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(G97), .C2(new_n1009), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G50), .A2(new_n766), .B1(new_n1013), .B2(G68), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n780), .A2(new_n336), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n758), .A2(new_n545), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G159), .B2(new_n776), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n412), .B1(G326), .B2(new_n793), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n758), .A2(new_n825), .B1(new_n782), .B2(new_n822), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n780), .A2(G311), .B1(new_n776), .B2(G322), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n795), .B2(new_n763), .C1(new_n1000), .C2(new_n765), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n1047), .B2(new_n1046), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1043), .B1(new_n512), .B2(new_n778), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1042), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1034), .B1(new_n1053), .B2(new_n751), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT110), .Z(new_n1055));
  AOI22_X1  g0855(.A1(new_n986), .A2(new_n969), .B1(new_n1025), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1024), .A2(new_n1056), .ZN(G393));
  NAND2_X1  g0857(.A1(new_n739), .A2(new_n243), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n752), .C1(new_n204), .C2(new_n212), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n765), .A2(new_n770), .B1(new_n777), .B2(new_n1015), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n780), .A2(G50), .B1(new_n1009), .B2(G87), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G68), .A2(new_n997), .B1(new_n757), .B2(G77), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n412), .B1(new_n829), .B2(new_n769), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n1013), .B2(new_n336), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n780), .A2(G303), .B1(new_n757), .B2(G116), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n822), .B2(new_n763), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT112), .Z(new_n1069));
  OAI21_X1  g0869(.A(new_n347), .B1(new_n769), .B2(new_n798), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G107), .B2(new_n1009), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(new_n782), .C2(new_n825), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n766), .A2(G311), .B1(G317), .B2(new_n776), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1066), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1075), .B(KEYINPUT113), .Z(new_n1076));
  OAI211_X1 g0876(.A(new_n732), .B(new_n1059), .C1(new_n1076), .C2(new_n819), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT114), .Z(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n802), .B2(new_n948), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n982), .A2(new_n983), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n730), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n986), .A2(new_n727), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT115), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT115), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1080), .A2(new_n1085), .A3(new_n1082), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n987), .A2(new_n1021), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1081), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(G390));
  AOI21_X1  g0890(.A(new_n927), .B1(new_n905), .B2(new_n892), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n725), .A2(new_n682), .A3(new_n808), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1092), .A2(new_n806), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n929), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n927), .B1(new_n930), .B2(new_n929), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1095), .B1(new_n926), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n863), .A2(G330), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n1098), .A2(new_n809), .A3(new_n1094), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n718), .A2(new_n857), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1095), .B(new_n1101), .C1(new_n926), .C2(new_n1096), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n969), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n817), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n732), .B1(new_n336), .B2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n766), .A2(G132), .B1(G128), .B2(new_n776), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT117), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n299), .B1(new_n769), .B2(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n781), .A2(new_n1011), .B1(new_n778), .B2(new_n268), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(G159), .C2(new_n757), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n997), .A2(G150), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT53), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT54), .B(G143), .Z(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n1013), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1107), .A2(new_n1111), .A3(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n780), .A2(G107), .B1(new_n776), .B2(G283), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n204), .B2(new_n763), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT118), .Z(new_n1119));
  OAI221_X1 g0919(.A(new_n347), .B1(new_n769), .B2(new_n822), .C1(new_n222), .C2(new_n782), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n835), .B(new_n1120), .C1(G77), .C2(new_n757), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n512), .B2(new_n765), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1116), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT119), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n819), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1105), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n926), .B2(new_n749), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1103), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1098), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n460), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n934), .A2(new_n1131), .A3(new_n667), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n929), .B1(new_n718), .B2(new_n811), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n930), .B1(new_n1133), .B2(new_n1099), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1094), .B1(new_n1098), .B2(new_n809), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1101), .A2(new_n1135), .A3(new_n1093), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1132), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT116), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1100), .A2(new_n1102), .A3(new_n1137), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1140), .A2(new_n1021), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1129), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(G378));
  AOI21_X1  g0943(.A(new_n731), .B1(new_n268), .B2(new_n817), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G128), .A2(new_n766), .B1(new_n1013), .B2(G137), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n776), .A2(G125), .B1(new_n757), .B2(G150), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n780), .A2(G132), .B1(new_n997), .B2(new_n1114), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1149), .A2(KEYINPUT59), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(KEYINPUT59), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1009), .A2(G159), .ZN(new_n1152));
  AOI211_X1 g0952(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n781), .A2(new_n204), .B1(new_n777), .B2(new_n512), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n778), .A2(new_n226), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G107), .A2(new_n766), .B1(new_n1013), .B2(new_n338), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n276), .B1(new_n769), .B2(new_n791), .ZN(new_n1159));
  NOR4_X1   g0959(.A1(new_n1007), .A2(new_n1159), .A3(new_n1035), .A4(new_n412), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT58), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n276), .B1(new_n411), .B2(new_n258), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n268), .ZN(new_n1166));
  AND4_X1   g0966(.A1(new_n1154), .A2(new_n1163), .A3(new_n1164), .A4(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n388), .B1(new_n391), .B2(new_n393), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n379), .A2(new_n672), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  OR3_X1    g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1144), .B1(new_n819), .B2(new_n1167), .C1(new_n1176), .C2(new_n749), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT120), .Z(new_n1178));
  AOI22_X1  g0978(.A1(new_n864), .A2(new_n865), .B1(new_n891), .B2(new_n892), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT40), .B1(new_n1179), .B2(new_n894), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n907), .A2(G330), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n1176), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1176), .ZN(new_n1183));
  INV_X1    g0983(.A(G330), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n898), .B2(new_n906), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1183), .B1(new_n897), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n931), .A2(new_n932), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n927), .B2(new_n926), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT121), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n1182), .A2(new_n1186), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1176), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n897), .A2(new_n1185), .A3(new_n1183), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n933), .A2(new_n1191), .A3(new_n1192), .A4(KEYINPUT121), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1178), .B1(new_n1194), .B2(new_n969), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1132), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1140), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n933), .B1(new_n1182), .B2(new_n1186), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1191), .A2(new_n1188), .A3(new_n1192), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(KEYINPUT57), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1021), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1140), .A2(new_n1196), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT57), .B1(new_n1194), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1195), .B1(new_n1201), .B2(new_n1203), .ZN(G375));
  NAND2_X1  g1004(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1094), .A2(new_n748), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n732), .B1(G68), .B2(new_n1104), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n781), .A2(new_n512), .B1(new_n777), .B2(new_n822), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1040), .B(new_n1208), .C1(G97), .C2(new_n997), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n347), .B1(new_n769), .B2(new_n795), .C1(new_n264), .C2(new_n778), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1013), .B2(G107), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(new_n791), .C2(new_n765), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT122), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n763), .A2(new_n1015), .B1(new_n758), .B2(new_n268), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT123), .Z(new_n1215));
  OAI22_X1  g1015(.A1(new_n777), .A2(new_n833), .B1(new_n782), .B2(new_n770), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1156), .B(new_n1216), .C1(new_n780), .C2(new_n1114), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n766), .A2(G137), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n509), .B1(G128), .B2(new_n793), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1215), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1212), .A2(KEYINPUT122), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1213), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1207), .B1(new_n1222), .B2(new_n751), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1205), .A2(new_n969), .B1(new_n1206), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1137), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n970), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1205), .A2(new_n1196), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1224), .B1(new_n1227), .B2(new_n1228), .ZN(G381));
  NOR3_X1   g1029(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1230));
  INV_X1    g1030(.A(G375), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1024), .A2(new_n804), .A3(new_n1056), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n842), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT124), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1230), .A2(new_n1142), .A3(new_n1231), .A4(new_n1235), .ZN(G407));
  NAND2_X1  g1036(.A1(new_n673), .A2(G213), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1231), .A2(new_n1142), .A3(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(G407), .A2(new_n1239), .A3(G213), .ZN(G409));
  INV_X1    g1040(.A(KEYINPUT116), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1241), .B(new_n1137), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT116), .B1(new_n1243), .B2(new_n1225), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1141), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1129), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1194), .A2(new_n1226), .A3(new_n1202), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1198), .A2(new_n969), .A3(new_n1199), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1177), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1245), .B(new_n1246), .C1(new_n1247), .C2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(G375), .B2(new_n1142), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT125), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1228), .A2(KEYINPUT60), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1205), .B2(new_n1196), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1253), .A2(new_n1021), .A3(new_n1225), .A4(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(G384), .A3(new_n1224), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G384), .B1(new_n1256), .B2(new_n1224), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT125), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1250), .B(new_n1261), .C1(G375), .C2(new_n1142), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1252), .A2(new_n1237), .A3(new_n1260), .A4(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT63), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1252), .A2(new_n1237), .A3(new_n1262), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1238), .A2(G2897), .ZN(new_n1267));
  OR3_X1    g1067(.A1(new_n1258), .A2(new_n1259), .A3(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1267), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1266), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(G390), .A2(new_n989), .A3(new_n1019), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G387), .A2(new_n1089), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(G393), .A2(G396), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(KEYINPUT126), .B1(new_n1276), .B2(new_n1233), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1275), .A2(new_n1278), .A3(new_n1232), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1273), .A2(new_n1274), .A3(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1277), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(KEYINPUT61), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1251), .A2(new_n1237), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(KEYINPUT63), .A3(new_n1260), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1265), .A2(new_n1272), .A3(new_n1285), .A4(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1289), .B1(new_n1286), .B2(new_n1270), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1263), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1286), .A2(KEYINPUT62), .A3(new_n1260), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1290), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1284), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1288), .B1(new_n1294), .B2(new_n1295), .ZN(G405));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1260), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1231), .A2(G378), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G375), .A2(new_n1142), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1298), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1260), .A2(new_n1297), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1299), .A2(new_n1297), .A3(new_n1260), .A4(new_n1300), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1305), .B(new_n1295), .ZN(G402));
endmodule


