

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784;

  BUF_X1 U370 ( .A(n723), .Z(n348) );
  XNOR2_X1 U371 ( .A(n635), .B(n634), .ZN(n690) );
  NAND2_X1 U372 ( .A1(n350), .A2(n349), .ZN(n552) );
  INV_X2 U373 ( .A(n562), .ZN(n350) );
  INV_X1 U374 ( .A(n551), .ZN(n349) );
  XNOR2_X1 U375 ( .A(n670), .B(KEYINPUT38), .ZN(n620) );
  NAND2_X1 U376 ( .A1(n423), .A2(n420), .ZN(n670) );
  AND2_X1 U377 ( .A1(n425), .A2(n424), .ZN(n423) );
  XNOR2_X1 U378 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n506) );
  XNOR2_X1 U379 ( .A(n621), .B(KEYINPUT39), .ZN(n411) );
  XOR2_X2 U380 ( .A(n700), .B(KEYINPUT59), .Z(n360) );
  XOR2_X2 U381 ( .A(KEYINPUT67), .B(n696), .Z(n697) );
  XNOR2_X2 U382 ( .A(n497), .B(G472), .ZN(n627) );
  XNOR2_X2 U383 ( .A(n591), .B(KEYINPUT35), .ZN(n782) );
  INV_X1 U384 ( .A(n692), .ZN(n397) );
  INV_X2 U385 ( .A(G953), .ZN(n763) );
  AND2_X1 U386 ( .A1(n412), .A2(KEYINPUT85), .ZN(n409) );
  NAND2_X1 U387 ( .A1(n374), .A2(n373), .ZN(n585) );
  XNOR2_X1 U388 ( .A(n558), .B(n557), .ZN(n586) );
  AND2_X1 U389 ( .A1(n385), .A2(n384), .ZN(n383) );
  XNOR2_X1 U390 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U391 ( .A(n370), .B(n369), .ZN(n723) );
  NOR2_X2 U392 ( .A1(n714), .A2(G902), .ZN(n388) );
  NOR2_X1 U393 ( .A1(n387), .A2(n604), .ZN(n605) );
  XNOR2_X1 U394 ( .A(n495), .B(n494), .ZN(n508) );
  XNOR2_X1 U395 ( .A(G119), .B(G113), .ZN(n495) );
  XNOR2_X1 U396 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n494) );
  XNOR2_X1 U397 ( .A(G122), .B(G116), .ZN(n522) );
  XNOR2_X1 U398 ( .A(n427), .B(n443), .ZN(n372) );
  INV_X1 U399 ( .A(KEYINPUT22), .ZN(n443) );
  XNOR2_X1 U400 ( .A(n598), .B(n362), .ZN(n647) );
  INV_X1 U401 ( .A(KEYINPUT6), .ZN(n362) );
  INV_X1 U402 ( .A(n687), .ZN(n417) );
  INV_X1 U403 ( .A(KEYINPUT0), .ZN(n379) );
  XNOR2_X1 U404 ( .A(KEYINPUT10), .B(n464), .ZN(n771) );
  XNOR2_X1 U405 ( .A(G140), .B(G125), .ZN(n464) );
  XNOR2_X1 U406 ( .A(KEYINPUT18), .B(G125), .ZN(n511) );
  INV_X1 U407 ( .A(KEYINPUT108), .ZN(n429) );
  NAND2_X1 U408 ( .A1(n397), .A2(n676), .ZN(n698) );
  NOR2_X1 U409 ( .A1(n675), .A2(n674), .ZN(n676) );
  OR2_X1 U410 ( .A1(n723), .A2(n421), .ZN(n420) );
  NAND2_X1 U411 ( .A1(n422), .A2(n694), .ZN(n421) );
  INV_X1 U412 ( .A(n519), .ZN(n422) );
  NAND2_X1 U413 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U414 ( .A(n383), .ZN(n380) );
  NAND2_X1 U415 ( .A1(n376), .A2(n379), .ZN(n375) );
  NAND2_X1 U416 ( .A1(n381), .A2(n377), .ZN(n376) );
  INV_X1 U417 ( .A(n581), .ZN(n377) );
  AND2_X1 U418 ( .A1(n576), .A2(n430), .ZN(n555) );
  INV_X1 U419 ( .A(n599), .ZN(n430) );
  XNOR2_X1 U420 ( .A(n458), .B(n689), .ZN(n491) );
  XNOR2_X1 U421 ( .A(G134), .B(G131), .ZN(n458) );
  XNOR2_X1 U422 ( .A(n508), .B(n492), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n509), .B(n508), .ZN(n762) );
  XNOR2_X1 U424 ( .A(G110), .B(G107), .ZN(n455) );
  INV_X1 U425 ( .A(n401), .ZN(n667) );
  AND2_X1 U426 ( .A1(n595), .A2(n594), .ZN(n387) );
  AND2_X1 U427 ( .A1(n372), .A2(n647), .ZN(n592) );
  XNOR2_X1 U428 ( .A(n753), .B(KEYINPUT88), .ZN(n654) );
  AND2_X1 U429 ( .A1(G953), .A2(G902), .ZN(n611) );
  NOR2_X1 U430 ( .A1(n499), .A2(n363), .ZN(n500) );
  AND2_X1 U431 ( .A1(n784), .A2(n416), .ZN(n415) );
  NAND2_X1 U432 ( .A1(n417), .A2(KEYINPUT86), .ZN(n416) );
  INV_X1 U433 ( .A(G237), .ZN(n516) );
  XNOR2_X1 U434 ( .A(G143), .B(G113), .ZN(n536) );
  XOR2_X1 U435 ( .A(G104), .B(G131), .Z(n537) );
  XNOR2_X1 U436 ( .A(G122), .B(KEYINPUT12), .ZN(n538) );
  XOR2_X1 U437 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n539) );
  NOR2_X1 U438 ( .A1(G953), .A2(G237), .ZN(n542) );
  XNOR2_X1 U439 ( .A(KEYINPUT96), .B(G140), .ZN(n460) );
  NOR2_X1 U440 ( .A1(n434), .A2(n435), .ZN(n606) );
  NAND2_X1 U441 ( .A1(n438), .A2(n605), .ZN(n434) );
  NAND2_X1 U442 ( .A1(n437), .A2(n436), .ZN(n435) );
  INV_X1 U443 ( .A(n598), .ZN(n363) );
  NAND2_X1 U444 ( .A1(n420), .A2(n639), .ZN(n405) );
  INV_X1 U445 ( .A(G902), .ZN(n547) );
  OR2_X1 U446 ( .A1(n644), .A2(n642), .ZN(n599) );
  XNOR2_X1 U447 ( .A(G134), .B(G107), .ZN(n528) );
  XNOR2_X1 U448 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U449 ( .A(n371), .B(n762), .ZN(n370) );
  XNOR2_X1 U450 ( .A(n514), .B(n454), .ZN(n371) );
  NAND2_X1 U451 ( .A1(G234), .A2(G237), .ZN(n570) );
  NOR2_X1 U452 ( .A1(n647), .A2(n556), .ZN(n558) );
  XNOR2_X1 U453 ( .A(n555), .B(n429), .ZN(n556) );
  NAND2_X1 U454 ( .A1(n352), .A2(n383), .ZN(n373) );
  AND2_X1 U455 ( .A1(n378), .A2(n375), .ZN(n374) );
  AND2_X1 U456 ( .A1(n555), .A2(n363), .ZN(n596) );
  NOR2_X1 U457 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U458 ( .A1(n423), .A2(n382), .ZN(n381) );
  NOR2_X1 U459 ( .A1(n405), .A2(n354), .ZN(n382) );
  XNOR2_X1 U460 ( .A(n535), .B(n534), .ZN(n589) );
  XNOR2_X1 U461 ( .A(G478), .B(KEYINPUT106), .ZN(n534) );
  XNOR2_X1 U462 ( .A(n600), .B(KEYINPUT99), .ZN(n618) );
  NOR2_X1 U463 ( .A1(n630), .A2(n599), .ZN(n600) );
  XNOR2_X1 U464 ( .A(n390), .B(n364), .ZN(n703) );
  XNOR2_X1 U465 ( .A(n493), .B(n365), .ZN(n364) );
  NAND2_X1 U466 ( .A1(n451), .A2(G221), .ZN(n450) );
  INV_X1 U467 ( .A(KEYINPUT83), .ZN(n681) );
  NAND2_X1 U468 ( .A1(n366), .A2(n353), .ZN(n753) );
  XNOR2_X1 U469 ( .A(n368), .B(n367), .ZN(n366) );
  INV_X1 U470 ( .A(KEYINPUT36), .ZN(n367) );
  NAND2_X1 U471 ( .A1(n668), .A2(n651), .ZN(n368) );
  AND2_X1 U472 ( .A1(n583), .A2(n353), .ZN(n442) );
  NAND2_X1 U473 ( .A1(n402), .A2(n351), .ZN(n691) );
  XNOR2_X1 U474 ( .A(n403), .B(KEYINPUT107), .ZN(n402) );
  INV_X1 U475 ( .A(KEYINPUT60), .ZN(n445) );
  XNOR2_X1 U476 ( .A(n387), .B(n386), .ZN(n730) );
  INV_X1 U477 ( .A(G101), .ZN(n386) );
  AND2_X1 U478 ( .A1(n598), .A2(n593), .ZN(n351) );
  AND2_X1 U479 ( .A1(n381), .A2(n355), .ZN(n352) );
  XOR2_X1 U480 ( .A(n401), .B(KEYINPUT91), .Z(n353) );
  INV_X1 U481 ( .A(n423), .ZN(n404) );
  XNOR2_X1 U482 ( .A(n771), .B(n465), .ZN(n545) );
  XOR2_X1 U483 ( .A(KEYINPUT19), .B(KEYINPUT68), .Z(n354) );
  NOR2_X1 U484 ( .A1(n581), .A2(n379), .ZN(n355) );
  AND2_X1 U485 ( .A1(n687), .A2(n672), .ZN(n356) );
  AND2_X1 U486 ( .A1(n442), .A2(n372), .ZN(n357) );
  INV_X1 U487 ( .A(G221), .ZN(n480) );
  XNOR2_X1 U488 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n358) );
  XOR2_X1 U489 ( .A(n622), .B(KEYINPUT40), .Z(n359) );
  INV_X1 U490 ( .A(n749), .ZN(n444) );
  XOR2_X1 U491 ( .A(G131), .B(KEYINPUT127), .Z(n361) );
  XNOR2_X1 U492 ( .A(n457), .B(n769), .ZN(n369) );
  NAND2_X1 U493 ( .A1(n372), .A2(n667), .ZN(n403) );
  NAND2_X1 U494 ( .A1(n383), .A2(n381), .ZN(n656) );
  NAND2_X1 U495 ( .A1(n405), .A2(n354), .ZN(n384) );
  NAND2_X1 U496 ( .A1(n404), .A2(n354), .ZN(n385) );
  XNOR2_X2 U497 ( .A(n388), .B(G469), .ZN(n630) );
  XNOR2_X1 U498 ( .A(n527), .B(n431), .ZN(n389) );
  XNOR2_X1 U499 ( .A(n389), .B(n454), .ZN(n390) );
  XNOR2_X1 U500 ( .A(n769), .B(n454), .ZN(n496) );
  XNOR2_X1 U501 ( .A(n396), .B(n699), .ZN(n391) );
  NAND2_X2 U502 ( .A1(n398), .A2(n698), .ZN(n396) );
  XNOR2_X1 U503 ( .A(n496), .B(n457), .ZN(n515) );
  XNOR2_X1 U504 ( .A(n606), .B(KEYINPUT45), .ZN(n692) );
  NAND2_X1 U505 ( .A1(n413), .A2(KEYINPUT86), .ZN(n392) );
  NAND2_X1 U506 ( .A1(n413), .A2(KEYINPUT86), .ZN(n412) );
  BUF_X1 U507 ( .A(n411), .Z(n393) );
  NAND2_X1 U508 ( .A1(n411), .A2(n747), .ZN(n623) );
  NOR2_X1 U509 ( .A1(n692), .A2(n694), .ZN(n400) );
  BUF_X1 U510 ( .A(n406), .Z(n394) );
  XNOR2_X1 U511 ( .A(n623), .B(n359), .ZN(n406) );
  NAND2_X1 U512 ( .A1(n447), .A2(n726), .ZN(n446) );
  XNOR2_X1 U513 ( .A(n448), .B(n360), .ZN(n447) );
  XNOR2_X1 U514 ( .A(n630), .B(n463), .ZN(n576) );
  BUF_X1 U515 ( .A(n576), .Z(n401) );
  INV_X1 U516 ( .A(n395), .ZN(n693) );
  AND2_X2 U517 ( .A1(n410), .A2(n408), .ZN(n395) );
  NAND2_X1 U518 ( .A1(n721), .A2(G475), .ZN(n448) );
  XNOR2_X2 U519 ( .A(n396), .B(n699), .ZN(n721) );
  NAND2_X1 U520 ( .A1(n399), .A2(n697), .ZN(n398) );
  NAND2_X1 U521 ( .A1(n395), .A2(n400), .ZN(n399) );
  NAND2_X1 U522 ( .A1(n406), .A2(n636), .ZN(n638) );
  XNOR2_X1 U523 ( .A(n394), .B(n361), .ZN(G33) );
  NAND2_X1 U524 ( .A1(n407), .A2(n678), .ZN(n410) );
  NAND2_X1 U525 ( .A1(n414), .A2(n392), .ZN(n407) );
  NAND2_X1 U526 ( .A1(n414), .A2(n392), .ZN(n675) );
  NAND2_X1 U527 ( .A1(n409), .A2(n414), .ZN(n408) );
  NAND2_X1 U528 ( .A1(n393), .A2(n444), .ZN(n673) );
  INV_X1 U529 ( .A(n419), .ZN(n413) );
  AND2_X2 U530 ( .A1(n418), .A2(n415), .ZN(n414) );
  NAND2_X1 U531 ( .A1(n419), .A2(n356), .ZN(n418) );
  XNOR2_X1 U532 ( .A(n666), .B(n665), .ZN(n419) );
  NAND2_X1 U533 ( .A1(n519), .A2(n426), .ZN(n424) );
  NAND2_X1 U534 ( .A1(n723), .A2(n519), .ZN(n425) );
  INV_X1 U535 ( .A(n694), .ZN(n426) );
  NAND2_X1 U536 ( .A1(n585), .A2(n453), .ZN(n427) );
  NAND2_X1 U537 ( .A1(n703), .A2(n547), .ZN(n497) );
  XNOR2_X2 U538 ( .A(n428), .B(G143), .ZN(n527) );
  XNOR2_X2 U539 ( .A(G128), .B(KEYINPUT65), .ZN(n428) );
  XNOR2_X1 U540 ( .A(n587), .B(n358), .ZN(n590) );
  XNOR2_X2 U541 ( .A(n527), .B(n431), .ZN(n769) );
  XNOR2_X2 U542 ( .A(n433), .B(n432), .ZN(n431) );
  XNOR2_X2 U543 ( .A(KEYINPUT64), .B(KEYINPUT70), .ZN(n432) );
  XNOR2_X2 U544 ( .A(KEYINPUT4), .B(G146), .ZN(n433) );
  NAND2_X1 U545 ( .A1(n441), .A2(KEYINPUT44), .ZN(n436) );
  NAND2_X1 U546 ( .A1(n782), .A2(KEYINPUT44), .ZN(n437) );
  NAND2_X1 U547 ( .A1(n440), .A2(n439), .ZN(n438) );
  INV_X1 U548 ( .A(n441), .ZN(n439) );
  NOR2_X1 U549 ( .A1(n782), .A2(KEYINPUT44), .ZN(n440) );
  NAND2_X1 U550 ( .A1(n691), .A2(n783), .ZN(n441) );
  XNOR2_X1 U551 ( .A(n446), .B(n445), .ZN(G60) );
  NAND2_X1 U552 ( .A1(n709), .A2(n547), .ZN(n479) );
  XNOR2_X1 U553 ( .A(n449), .B(n545), .ZN(n709) );
  XNOR2_X1 U554 ( .A(n452), .B(n450), .ZN(n449) );
  INV_X1 U555 ( .A(n521), .ZN(n451) );
  XNOR2_X1 U556 ( .A(n472), .B(n468), .ZN(n452) );
  NOR2_X1 U557 ( .A1(n582), .A2(n642), .ZN(n453) );
  INV_X1 U558 ( .A(KEYINPUT85), .ZN(n678) );
  INV_X1 U559 ( .A(KEYINPUT2), .ZN(n674) );
  INV_X1 U560 ( .A(KEYINPUT1), .ZN(n463) );
  XNOR2_X1 U561 ( .A(n619), .B(KEYINPUT78), .ZN(n648) );
  XNOR2_X1 U562 ( .A(n526), .B(n525), .ZN(n533) );
  XNOR2_X1 U563 ( .A(n682), .B(n681), .ZN(n683) );
  INV_X1 U564 ( .A(KEYINPUT32), .ZN(n584) );
  XOR2_X1 U565 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n505) );
  XNOR2_X1 U566 ( .A(KEYINPUT69), .B(G101), .ZN(n454) );
  XNOR2_X1 U567 ( .A(n455), .B(G104), .ZN(n760) );
  XNOR2_X1 U568 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n456) );
  XNOR2_X1 U569 ( .A(n760), .B(n456), .ZN(n457) );
  INV_X1 U570 ( .A(G137), .ZN(n689) );
  XNOR2_X1 U571 ( .A(n491), .B(KEYINPUT95), .ZN(n770) );
  NAND2_X1 U572 ( .A1(n763), .A2(G227), .ZN(n459) );
  XNOR2_X1 U573 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U574 ( .A(n770), .B(n461), .ZN(n462) );
  XNOR2_X1 U575 ( .A(n515), .B(n462), .ZN(n714) );
  INV_X1 U576 ( .A(G146), .ZN(n465) );
  XNOR2_X2 U577 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n467) );
  XNOR2_X2 U578 ( .A(KEYINPUT79), .B(KEYINPUT97), .ZN(n466) );
  XNOR2_X1 U579 ( .A(n467), .B(n466), .ZN(n468) );
  NAND2_X1 U580 ( .A1(n763), .A2(G234), .ZN(n469) );
  XNOR2_X1 U581 ( .A(n469), .B(KEYINPUT8), .ZN(n521) );
  XNOR2_X2 U582 ( .A(G128), .B(G110), .ZN(n471) );
  XNOR2_X2 U583 ( .A(G119), .B(G137), .ZN(n470) );
  XNOR2_X1 U584 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X2 U585 ( .A(G902), .B(KEYINPUT15), .ZN(n694) );
  NAND2_X1 U586 ( .A1(n694), .A2(G234), .ZN(n474) );
  INV_X1 U587 ( .A(KEYINPUT20), .ZN(n473) );
  XNOR2_X1 U588 ( .A(n474), .B(n473), .ZN(n481) );
  INV_X1 U589 ( .A(n481), .ZN(n475) );
  NAND2_X1 U590 ( .A1(n475), .A2(G217), .ZN(n477) );
  XNOR2_X1 U591 ( .A(KEYINPUT98), .B(KEYINPUT25), .ZN(n476) );
  XNOR2_X1 U592 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U593 ( .A(n479), .B(n478), .ZN(n644) );
  OR2_X1 U594 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U595 ( .A(n482), .B(KEYINPUT21), .ZN(n642) );
  NAND2_X1 U596 ( .A1(n667), .A2(n599), .ZN(n483) );
  XOR2_X1 U597 ( .A(KEYINPUT50), .B(n483), .Z(n502) );
  INV_X1 U598 ( .A(KEYINPUT101), .ZN(n484) );
  NAND2_X1 U599 ( .A1(G116), .A2(n484), .ZN(n487) );
  INV_X1 U600 ( .A(G116), .ZN(n485) );
  NAND2_X1 U601 ( .A1(n485), .A2(KEYINPUT101), .ZN(n486) );
  NAND2_X1 U602 ( .A1(n487), .A2(n486), .ZN(n489) );
  XNOR2_X1 U603 ( .A(KEYINPUT100), .B(KEYINPUT5), .ZN(n488) );
  XNOR2_X1 U604 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U605 ( .A(n491), .B(n490), .ZN(n493) );
  NAND2_X1 U606 ( .A1(n542), .A2(G210), .ZN(n492) );
  INV_X1 U607 ( .A(n627), .ZN(n598) );
  BUF_X1 U608 ( .A(n644), .Z(n593) );
  NAND2_X1 U609 ( .A1(n593), .A2(n642), .ZN(n498) );
  XNOR2_X1 U610 ( .A(n498), .B(KEYINPUT49), .ZN(n499) );
  XNOR2_X1 U611 ( .A(KEYINPUT119), .B(n500), .ZN(n501) );
  NOR2_X1 U612 ( .A1(n502), .A2(n501), .ZN(n503) );
  NOR2_X1 U613 ( .A1(n503), .A2(n596), .ZN(n504) );
  XOR2_X1 U614 ( .A(n505), .B(n504), .Z(n553) );
  XNOR2_X1 U615 ( .A(n506), .B(KEYINPUT16), .ZN(n507) );
  XNOR2_X1 U616 ( .A(n507), .B(n522), .ZN(n509) );
  NAND2_X1 U617 ( .A1(n763), .A2(G224), .ZN(n510) );
  XNOR2_X1 U618 ( .A(n511), .B(n510), .ZN(n513) );
  XNOR2_X1 U619 ( .A(KEYINPUT92), .B(KEYINPUT17), .ZN(n512) );
  XNOR2_X1 U620 ( .A(n513), .B(n512), .ZN(n514) );
  NAND2_X1 U621 ( .A1(n547), .A2(n516), .ZN(n550) );
  NAND2_X1 U622 ( .A1(n550), .A2(G210), .ZN(n518) );
  XNOR2_X1 U623 ( .A(KEYINPUT81), .B(KEYINPUT93), .ZN(n517) );
  XNOR2_X1 U624 ( .A(n518), .B(n517), .ZN(n519) );
  INV_X1 U625 ( .A(n620), .ZN(n562) );
  INV_X1 U626 ( .A(G217), .ZN(n520) );
  OR2_X1 U627 ( .A1(n521), .A2(n520), .ZN(n526) );
  XNOR2_X1 U628 ( .A(n522), .B(KEYINPUT104), .ZN(n524) );
  XOR2_X1 U629 ( .A(KEYINPUT9), .B(KEYINPUT105), .Z(n523) );
  INV_X1 U630 ( .A(n527), .ZN(n531) );
  XOR2_X1 U631 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n529) );
  XNOR2_X1 U632 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U633 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U634 ( .A(n533), .B(n532), .ZN(n711) );
  NOR2_X1 U635 ( .A1(n711), .A2(G902), .ZN(n535) );
  XNOR2_X1 U636 ( .A(n537), .B(n536), .ZN(n541) );
  XNOR2_X1 U637 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U638 ( .A(n541), .B(n540), .Z(n544) );
  NAND2_X1 U639 ( .A1(G214), .A2(n542), .ZN(n543) );
  XNOR2_X1 U640 ( .A(n544), .B(n543), .ZN(n546) );
  XNOR2_X1 U641 ( .A(n546), .B(n545), .ZN(n700) );
  NAND2_X1 U642 ( .A1(n700), .A2(n547), .ZN(n549) );
  XOR2_X1 U643 ( .A(KEYINPUT13), .B(G475), .Z(n548) );
  XNOR2_X1 U644 ( .A(n549), .B(n548), .ZN(n560) );
  INV_X1 U645 ( .A(n560), .ZN(n588) );
  NAND2_X1 U646 ( .A1(n589), .A2(n588), .ZN(n582) );
  AND2_X1 U647 ( .A1(n550), .A2(G214), .ZN(n577) );
  OR2_X1 U648 ( .A1(n582), .A2(n577), .ZN(n551) );
  XNOR2_X2 U649 ( .A(n552), .B(KEYINPUT41), .ZN(n633) );
  NAND2_X1 U650 ( .A1(n553), .A2(n633), .ZN(n554) );
  XNOR2_X1 U651 ( .A(n554), .B(KEYINPUT121), .ZN(n568) );
  XOR2_X1 U652 ( .A(KEYINPUT33), .B(KEYINPUT90), .Z(n557) );
  INV_X1 U653 ( .A(n586), .ZN(n566) );
  INV_X1 U654 ( .A(n577), .ZN(n639) );
  NOR2_X1 U655 ( .A1(n620), .A2(n639), .ZN(n559) );
  NOR2_X1 U656 ( .A1(n559), .A2(n582), .ZN(n564) );
  AND2_X1 U657 ( .A1(n589), .A2(n560), .ZN(n747) );
  INV_X1 U658 ( .A(n747), .ZN(n744) );
  OR2_X1 U659 ( .A1(n589), .A2(n560), .ZN(n749) );
  NAND2_X1 U660 ( .A1(n744), .A2(n749), .ZN(n658) );
  NAND2_X1 U661 ( .A1(n658), .A2(n639), .ZN(n561) );
  NOR2_X1 U662 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U663 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U664 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U665 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U666 ( .A(KEYINPUT52), .B(n569), .ZN(n572) );
  XNOR2_X1 U667 ( .A(KEYINPUT14), .B(n570), .ZN(n615) );
  NAND2_X1 U668 ( .A1(G952), .A2(n615), .ZN(n571) );
  NOR2_X1 U669 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U670 ( .A1(G953), .A2(n573), .ZN(n575) );
  NAND2_X1 U671 ( .A1(n586), .A2(n633), .ZN(n574) );
  NAND2_X1 U672 ( .A1(n575), .A2(n574), .ZN(n684) );
  XNOR2_X1 U673 ( .A(G898), .B(KEYINPUT94), .ZN(n764) );
  INV_X1 U674 ( .A(n764), .ZN(n578) );
  NAND2_X1 U675 ( .A1(n578), .A2(n611), .ZN(n579) );
  NAND2_X1 U676 ( .A1(n763), .A2(G952), .ZN(n612) );
  NAND2_X1 U677 ( .A1(n579), .A2(n612), .ZN(n580) );
  NAND2_X1 U678 ( .A1(n580), .A2(n615), .ZN(n581) );
  AND2_X1 U679 ( .A1(n647), .A2(n593), .ZN(n583) );
  XNOR2_X1 U680 ( .A(n357), .B(n584), .ZN(n783) );
  NAND2_X1 U681 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U682 ( .A1(n589), .A2(n588), .ZN(n650) );
  NAND2_X1 U683 ( .A1(n590), .A2(n650), .ZN(n591) );
  XOR2_X1 U684 ( .A(KEYINPUT89), .B(n592), .Z(n595) );
  NOR2_X1 U685 ( .A1(n401), .A2(n593), .ZN(n594) );
  NAND2_X1 U686 ( .A1(n585), .A2(n596), .ZN(n597) );
  XNOR2_X1 U687 ( .A(n597), .B(KEYINPUT31), .ZN(n750) );
  NAND2_X1 U688 ( .A1(n598), .A2(n585), .ZN(n731) );
  BUF_X1 U689 ( .A(n618), .Z(n601) );
  NOR2_X1 U690 ( .A1(n731), .A2(n601), .ZN(n602) );
  OR2_X1 U691 ( .A1(n750), .A2(n602), .ZN(n603) );
  AND2_X1 U692 ( .A1(n603), .A2(n658), .ZN(n604) );
  NAND2_X1 U693 ( .A1(n692), .A2(n674), .ZN(n607) );
  XNOR2_X1 U694 ( .A(n607), .B(KEYINPUT82), .ZN(n677) );
  NAND2_X1 U695 ( .A1(n627), .A2(n639), .ZN(n609) );
  INV_X1 U696 ( .A(KEYINPUT30), .ZN(n608) );
  XNOR2_X1 U697 ( .A(n609), .B(n608), .ZN(n616) );
  INV_X1 U698 ( .A(G900), .ZN(n610) );
  NAND2_X1 U699 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U700 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U701 ( .A1(n615), .A2(n614), .ZN(n624) );
  INV_X1 U702 ( .A(n624), .ZN(n640) );
  NAND2_X1 U703 ( .A1(n616), .A2(n640), .ZN(n617) );
  NAND2_X1 U704 ( .A1(n648), .A2(n620), .ZN(n621) );
  INV_X1 U705 ( .A(KEYINPUT110), .ZN(n622) );
  NOR2_X1 U706 ( .A1(n642), .A2(n624), .ZN(n625) );
  AND2_X1 U707 ( .A1(n644), .A2(n625), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n629) );
  XOR2_X1 U709 ( .A(KEYINPUT28), .B(KEYINPUT109), .Z(n628) );
  XNOR2_X1 U710 ( .A(n629), .B(n628), .ZN(n631) );
  OR2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n655) );
  INV_X1 U712 ( .A(n655), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n635) );
  XNOR2_X1 U714 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n634) );
  INV_X1 U715 ( .A(n690), .ZN(n636) );
  INV_X1 U716 ( .A(KEYINPUT46), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n638), .B(n637), .ZN(n664) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U720 ( .A1(n593), .A2(n643), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n747), .A2(n645), .ZN(n646) );
  NOR2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n668) );
  INV_X1 U723 ( .A(n670), .ZN(n651) );
  BUF_X1 U724 ( .A(n648), .Z(n649) );
  INV_X1 U725 ( .A(n649), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n652) );
  OR2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n688) );
  NAND2_X1 U728 ( .A1(n654), .A2(n688), .ZN(n662) );
  OR2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n657), .B(KEYINPUT80), .ZN(n745) );
  INV_X1 U731 ( .A(n658), .ZN(n659) );
  OR2_X1 U732 ( .A1(n745), .A2(n659), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(KEYINPUT47), .ZN(n661) );
  NOR2_X1 U734 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n666) );
  XNOR2_X1 U736 ( .A(KEYINPUT71), .B(KEYINPUT48), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n669), .B(KEYINPUT43), .ZN(n671) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n687) );
  INV_X1 U740 ( .A(KEYINPUT86), .ZN(n672) );
  XNOR2_X1 U741 ( .A(n673), .B(KEYINPUT112), .ZN(n784) );
  NAND2_X1 U742 ( .A1(n677), .A2(n698), .ZN(n680) );
  AND2_X1 U743 ( .A1(n693), .A2(n674), .ZN(n679) );
  NOR2_X1 U744 ( .A1(n680), .A2(n679), .ZN(n682) );
  NOR2_X1 U745 ( .A1(n684), .A2(n683), .ZN(n686) );
  XNOR2_X1 U746 ( .A(KEYINPUT53), .B(KEYINPUT122), .ZN(n685) );
  XNOR2_X1 U747 ( .A(n686), .B(n685), .ZN(G75) );
  XNOR2_X1 U748 ( .A(n687), .B(G140), .ZN(G42) );
  XNOR2_X1 U749 ( .A(n688), .B(G143), .ZN(G45) );
  XNOR2_X1 U750 ( .A(n690), .B(n689), .ZN(G39) );
  XNOR2_X1 U751 ( .A(n691), .B(G110), .ZN(G12) );
  XOR2_X1 U752 ( .A(KEYINPUT84), .B(n694), .Z(n695) );
  NAND2_X1 U753 ( .A1(n695), .A2(KEYINPUT2), .ZN(n696) );
  INV_X1 U754 ( .A(KEYINPUT66), .ZN(n699) );
  INV_X1 U755 ( .A(G952), .ZN(n701) );
  NAND2_X1 U756 ( .A1(n701), .A2(G953), .ZN(n726) );
  INV_X1 U757 ( .A(n726), .ZN(n719) );
  NAND2_X1 U758 ( .A1(n721), .A2(G472), .ZN(n705) );
  XOR2_X1 U759 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n702) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(n706) );
  NAND2_X1 U761 ( .A1(n706), .A2(n726), .ZN(n707) );
  XNOR2_X1 U762 ( .A(n707), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U763 ( .A1(n391), .A2(G217), .ZN(n708) );
  XOR2_X1 U764 ( .A(n709), .B(n708), .Z(n710) );
  NOR2_X1 U765 ( .A1(n710), .A2(n719), .ZN(G66) );
  NAND2_X1 U766 ( .A1(n391), .A2(G478), .ZN(n712) );
  XNOR2_X1 U767 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U768 ( .A1(n713), .A2(n719), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n391), .A2(G469), .ZN(n718) );
  BUF_X1 U770 ( .A(n714), .Z(n716) );
  XOR2_X1 U771 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n715) );
  XNOR2_X1 U772 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U773 ( .A(n718), .B(n717), .ZN(n720) );
  NOR2_X1 U774 ( .A1(n720), .A2(n719), .ZN(G54) );
  NAND2_X1 U775 ( .A1(n721), .A2(G210), .ZN(n725) );
  XNOR2_X1 U776 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n722) );
  XNOR2_X1 U777 ( .A(n348), .B(n722), .ZN(n724) );
  XNOR2_X1 U778 ( .A(n725), .B(n724), .ZN(n727) );
  NAND2_X1 U779 ( .A1(n727), .A2(n726), .ZN(n729) );
  XNOR2_X1 U780 ( .A(KEYINPUT87), .B(KEYINPUT56), .ZN(n728) );
  XNOR2_X1 U781 ( .A(n729), .B(n728), .ZN(G51) );
  XNOR2_X1 U782 ( .A(KEYINPUT114), .B(n730), .ZN(G3) );
  INV_X1 U783 ( .A(n731), .ZN(n738) );
  NOR2_X1 U784 ( .A1(n601), .A2(n744), .ZN(n732) );
  NAND2_X1 U785 ( .A1(n738), .A2(n732), .ZN(n733) );
  XNOR2_X1 U786 ( .A(n733), .B(G104), .ZN(G6) );
  XOR2_X1 U787 ( .A(KEYINPUT27), .B(KEYINPUT116), .Z(n735) );
  XNOR2_X1 U788 ( .A(G107), .B(KEYINPUT115), .ZN(n734) );
  XNOR2_X1 U789 ( .A(n735), .B(n734), .ZN(n736) );
  XOR2_X1 U790 ( .A(KEYINPUT26), .B(n736), .Z(n740) );
  NOR2_X1 U791 ( .A1(n601), .A2(n749), .ZN(n737) );
  NAND2_X1 U792 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U793 ( .A(n740), .B(n739), .ZN(G9) );
  NOR2_X1 U794 ( .A1(n745), .A2(n749), .ZN(n742) );
  XNOR2_X1 U795 ( .A(KEYINPUT117), .B(KEYINPUT29), .ZN(n741) );
  XNOR2_X1 U796 ( .A(n742), .B(n741), .ZN(n743) );
  XOR2_X1 U797 ( .A(G128), .B(n743), .Z(G30) );
  NOR2_X1 U798 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U799 ( .A(G146), .B(n746), .Z(G48) );
  NAND2_X1 U800 ( .A1(n750), .A2(n747), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n748), .B(G113), .ZN(G15) );
  NAND2_X1 U802 ( .A1(n750), .A2(n444), .ZN(n751) );
  XNOR2_X1 U803 ( .A(n751), .B(G116), .ZN(G18) );
  XOR2_X1 U804 ( .A(KEYINPUT118), .B(KEYINPUT37), .Z(n752) );
  XNOR2_X1 U805 ( .A(n753), .B(n752), .ZN(n754) );
  XNOR2_X1 U806 ( .A(G125), .B(n754), .ZN(G27) );
  NAND2_X1 U807 ( .A1(n397), .A2(n763), .ZN(n758) );
  NAND2_X1 U808 ( .A1(G953), .A2(G224), .ZN(n755) );
  XNOR2_X1 U809 ( .A(n755), .B(KEYINPUT61), .ZN(n756) );
  NAND2_X1 U810 ( .A1(n756), .A2(n764), .ZN(n757) );
  NAND2_X1 U811 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U812 ( .A(n759), .B(KEYINPUT123), .ZN(n768) );
  XOR2_X1 U813 ( .A(G101), .B(n760), .Z(n761) );
  XNOR2_X1 U814 ( .A(n762), .B(n761), .ZN(n766) );
  NOR2_X1 U815 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U816 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U817 ( .A(n768), .B(n767), .Z(G69) );
  XOR2_X1 U818 ( .A(n771), .B(n770), .Z(n772) );
  XNOR2_X1 U819 ( .A(KEYINPUT124), .B(n772), .ZN(n773) );
  XNOR2_X1 U820 ( .A(n389), .B(n773), .ZN(n776) );
  XNOR2_X1 U821 ( .A(n693), .B(n776), .ZN(n774) );
  NOR2_X1 U822 ( .A1(n774), .A2(G953), .ZN(n775) );
  XNOR2_X1 U823 ( .A(KEYINPUT125), .B(n775), .ZN(n781) );
  XOR2_X1 U824 ( .A(G227), .B(n776), .Z(n777) );
  NAND2_X1 U825 ( .A1(n777), .A2(G900), .ZN(n778) );
  NAND2_X1 U826 ( .A1(G953), .A2(n778), .ZN(n779) );
  XNOR2_X1 U827 ( .A(KEYINPUT126), .B(n779), .ZN(n780) );
  NAND2_X1 U828 ( .A1(n781), .A2(n780), .ZN(G72) );
  XOR2_X1 U829 ( .A(n782), .B(G122), .Z(G24) );
  XNOR2_X1 U830 ( .A(G119), .B(n783), .ZN(G21) );
  XNOR2_X1 U831 ( .A(G134), .B(n784), .ZN(G36) );
endmodule

