//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT67), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT2), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G116), .B(G119), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n195), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  OAI22_X1  g016(.A1(new_n194), .A2(new_n202), .B1(new_n201), .B2(new_n200), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(G146), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G143), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G128), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT66), .B(G128), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(G143), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n207), .B2(G143), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n210), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G134), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G137), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT11), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n220), .B2(G137), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(G137), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n222), .A2(new_n223), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n226), .ZN(new_n228));
  OAI21_X1  g042(.A(G131), .B1(new_n228), .B2(new_n221), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n217), .A2(new_n233), .B1(new_n208), .B2(new_n231), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n222), .A2(new_n225), .A3(new_n226), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n227), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n219), .A2(new_n230), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n204), .B(KEYINPUT30), .C1(new_n238), .C2(KEYINPUT64), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n219), .A2(new_n230), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT68), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT30), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n242), .B2(KEYINPUT68), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n203), .B(new_n239), .C1(new_n244), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n203), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT67), .B1(new_n192), .B2(new_n193), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n200), .A2(new_n201), .A3(new_n195), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n250), .A2(new_n251), .B1(new_n192), .B2(new_n193), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT69), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n240), .A2(new_n249), .A3(new_n241), .A4(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n256));
  NOR2_X1   g070(.A1(G237), .A2(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G210), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n256), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  XOR2_X1   g074(.A(new_n259), .B(new_n260), .Z(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n254), .A2(KEYINPUT28), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n254), .A2(KEYINPUT28), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n238), .A2(new_n252), .ZN(new_n267));
  OR3_X1    g081(.A1(new_n266), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT29), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n263), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n249), .A2(new_n253), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n242), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(new_n264), .B2(new_n265), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n273), .A2(new_n269), .A3(new_n262), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G902), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n187), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n254), .A2(KEYINPUT71), .A3(new_n261), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT71), .B1(new_n254), .B2(new_n261), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT31), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n247), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n280), .B2(new_n247), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n282), .B(new_n283), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  AOI211_X1 g100(.A(KEYINPUT72), .B(new_n281), .C1(new_n280), .C2(new_n247), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n187), .B(new_n277), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT32), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n280), .A2(new_n247), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT31), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT72), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n284), .A2(new_n285), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n282), .A4(new_n283), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n187), .A4(new_n277), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n276), .B1(new_n289), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n211), .A2(G119), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(new_n188), .B2(G128), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT24), .B(G110), .Z(new_n301));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n302), .B1(new_n188), .B2(G128), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI22_X1  g120(.A1(new_n303), .A2(new_n304), .B1(new_n188), .B2(G128), .ZN(new_n307));
  OAI22_X1  g121(.A1(new_n306), .A2(new_n307), .B1(new_n302), .B2(new_n298), .ZN(new_n308));
  OAI22_X1  g122(.A1(new_n300), .A2(new_n301), .B1(new_n308), .B2(G110), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(KEYINPUT74), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(G125), .A3(G140), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(KEYINPUT16), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT16), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n311), .B2(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G146), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n207), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT76), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n207), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n309), .A2(new_n319), .A3(new_n325), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n300), .A2(new_n301), .B1(new_n308), .B2(G110), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT75), .B1(new_n318), .B2(G146), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n315), .A2(new_n329), .A3(new_n205), .A4(new_n317), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n330), .A3(new_n319), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT77), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT22), .B(G137), .ZN(new_n336));
  INV_X1    g150(.A(G953), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n337), .A2(G221), .A3(G234), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n336), .B(new_n338), .Z(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n326), .A2(new_n332), .A3(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n334), .A2(new_n335), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n326), .A2(new_n332), .A3(new_n339), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n334), .A2(new_n340), .A3(new_n342), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT78), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G217), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(G234), .B2(new_n277), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(G902), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n347), .A2(new_n277), .A3(new_n344), .A4(new_n343), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n345), .A2(KEYINPUT25), .A3(new_n277), .A4(new_n347), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n353), .B1(new_n358), .B2(new_n350), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n297), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n362));
  XNOR2_X1  g176(.A(G113), .B(G122), .ZN(new_n363));
  INV_X1    g177(.A(G104), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G237), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n337), .A3(G214), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n214), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n257), .A2(G143), .A3(G214), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT18), .A2(G131), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(KEYINPUT91), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n312), .A2(new_n314), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G146), .ZN(new_n374));
  INV_X1    g188(.A(new_n324), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n323), .B1(new_n207), .B2(new_n320), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n368), .A2(new_n369), .ZN(new_n378));
  INV_X1    g192(.A(new_n370), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n372), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n325), .A2(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT92), .A3(new_n372), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n378), .A2(G131), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n368), .A2(new_n223), .A3(new_n369), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  MUX2_X1   g203(.A(new_n320), .B(new_n373), .S(KEYINPUT19), .Z(new_n390));
  INV_X1    g204(.A(new_n207), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n389), .B(new_n319), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n365), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n378), .A2(KEYINPUT17), .A3(G131), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n389), .B2(KEYINPUT17), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n396), .A2(new_n331), .ZN(new_n397));
  AND4_X1   g211(.A1(KEYINPUT92), .A2(new_n372), .A3(new_n377), .A4(new_n380), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT92), .B1(new_n384), .B2(new_n372), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n397), .B(new_n365), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT93), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n396), .A2(new_n331), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n383), .B2(new_n385), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT93), .B1(new_n404), .B2(new_n365), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n394), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(G475), .A2(G902), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n362), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n400), .A2(new_n401), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n386), .A2(KEYINPUT93), .A3(new_n365), .A4(new_n397), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n393), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n407), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n411), .A2(KEYINPUT20), .A3(new_n412), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n404), .A2(new_n365), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n409), .B2(new_n410), .ZN(new_n416));
  OAI21_X1  g230(.A(G475), .B1(new_n416), .B2(G902), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT95), .B(G952), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(G953), .ZN(new_n419));
  NAND2_X1  g233(.A1(G234), .A2(G237), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(G898), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(G902), .A3(G953), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n422), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n414), .A2(new_n417), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n214), .A2(G128), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n429), .B(KEYINPUT13), .Z(new_n430));
  NAND2_X1  g244(.A1(new_n211), .A2(G143), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G134), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G116), .B(G122), .ZN(new_n434));
  INV_X1    g248(.A(G107), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n429), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n433), .B(new_n436), .C1(G134), .C2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT14), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n190), .A2(KEYINPUT14), .A3(G122), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(G107), .A3(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n442), .A2(KEYINPUT94), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(KEYINPUT94), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n434), .A2(new_n435), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n437), .A2(G134), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n220), .B1(new_n431), .B2(new_n429), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n438), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT9), .B(G234), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n451), .A2(new_n349), .A3(G953), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n438), .B(new_n452), .C1(new_n445), .C2(new_n449), .ZN(new_n455));
  AOI21_X1  g269(.A(G902), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G478), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(KEYINPUT15), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n428), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G214), .B1(G237), .B2(G902), .ZN(new_n462));
  OAI21_X1  g276(.A(G210), .B1(G237), .B2(G902), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n435), .A2(G104), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n364), .A2(G107), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT80), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT3), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n468), .A2(new_n435), .A3(KEYINPUT3), .A4(G104), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n466), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT4), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n472), .A2(KEYINPUT82), .A3(new_n473), .A4(G101), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT82), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n468), .A2(new_n435), .A3(G104), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n465), .B1(new_n478), .B2(new_n470), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n473), .A2(G101), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n252), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n465), .A2(G101), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n469), .B2(new_n471), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g299(.A(G101), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n478), .A2(new_n470), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(new_n466), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n485), .A2(new_n488), .A3(KEYINPUT81), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT81), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n472), .A2(G101), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n473), .B1(new_n487), .B2(new_n483), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n482), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n467), .A2(new_n465), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n484), .B1(new_n486), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n194), .A2(new_n202), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n201), .A2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G113), .B1(new_n189), .B2(KEYINPUT5), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n496), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G110), .B(G122), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n464), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n494), .A2(new_n505), .A3(new_n503), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(KEYINPUT87), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT87), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT81), .B1(new_n485), .B2(new_n488), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n491), .A2(new_n490), .A3(new_n492), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n502), .B1(new_n513), .B2(new_n482), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n510), .B1(new_n514), .B2(new_n505), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n507), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n210), .B(new_n311), .C1(new_n213), .C2(new_n218), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n234), .A2(new_n311), .ZN(new_n519));
  OAI211_X1 g333(.A(G224), .B(new_n337), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G224), .ZN(new_n521));
  OAI221_X1 g335(.A(new_n517), .B1(new_n311), .B2(new_n234), .C1(new_n521), .C2(G953), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n514), .A2(KEYINPUT6), .A3(new_n505), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n516), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT88), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n508), .A2(KEYINPUT87), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n514), .A2(new_n510), .A3(new_n505), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n524), .B1(new_n530), .B2(new_n507), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n523), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n505), .B(KEYINPUT8), .Z(new_n535));
  NOR2_X1   g349(.A1(new_n497), .A2(new_n501), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(new_n496), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n498), .A2(KEYINPUT89), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n500), .B1(new_n498), .B2(KEYINPUT89), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n538), .A2(new_n539), .B1(new_n251), .B2(new_n250), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT90), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n496), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n537), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT7), .B1(new_n337), .B2(G224), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n518), .B2(new_n519), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n520), .B2(new_n522), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(G902), .B1(new_n550), .B2(new_n530), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n463), .B1(new_n534), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n463), .ZN(new_n553));
  INV_X1    g367(.A(new_n551), .ZN(new_n554));
  AOI211_X1 g368(.A(new_n553), .B(new_n554), .C1(new_n527), .C2(new_n533), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n462), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G221), .B1(new_n451), .B2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n210), .A2(KEYINPUT83), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT83), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n208), .A2(new_n561), .A3(new_n209), .A4(G128), .ZN(new_n562));
  INV_X1    g376(.A(new_n208), .ZN(new_n563));
  OAI21_X1  g377(.A(G128), .B1(new_n215), .B2(new_n209), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n560), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n543), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n496), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n567), .A2(new_n568), .B1(new_n219), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n474), .A2(new_n481), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n513), .A2(new_n234), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n237), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(G110), .B(G140), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n337), .A2(G227), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n573), .B1(new_n570), .B2(new_n572), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n577), .B(KEYINPUT79), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n210), .A2(KEYINPUT83), .B1(new_n563), .B2(new_n564), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n496), .B1(new_n584), .B2(new_n562), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n543), .A2(new_n219), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n237), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT84), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT12), .B1(new_n237), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  OAI221_X1 g404(.A(new_n237), .B1(new_n588), .B2(KEYINPUT12), .C1(new_n585), .C2(new_n586), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n583), .B1(new_n592), .B2(new_n574), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n277), .B1(new_n581), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G469), .ZN(new_n595));
  INV_X1    g409(.A(new_n574), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n577), .B1(new_n596), .B2(new_n580), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n592), .A2(new_n574), .A3(new_n578), .ZN(new_n598));
  AOI21_X1  g412(.A(G902), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT86), .B(G469), .Z(new_n600));
  AOI22_X1  g414(.A1(new_n595), .A2(KEYINPUT85), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT85), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n594), .A2(new_n602), .A3(G469), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n559), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n361), .A2(new_n461), .A3(new_n557), .A4(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  NAND2_X1  g420(.A1(new_n556), .A2(KEYINPUT96), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n532), .B1(new_n531), .B2(new_n523), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT6), .B1(new_n514), .B2(new_n505), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n529), .B2(new_n528), .ZN(new_n610));
  INV_X1    g424(.A(new_n523), .ZN(new_n611));
  NOR4_X1   g425(.A1(new_n610), .A2(KEYINPUT88), .A3(new_n611), .A4(new_n524), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n551), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n553), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n534), .A2(new_n463), .A3(new_n551), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n462), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n607), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n417), .B1(new_n408), .B2(new_n413), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n454), .A2(new_n455), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT33), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n454), .A2(new_n623), .A3(new_n455), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(G478), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n457), .A2(new_n277), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n456), .B2(new_n457), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT97), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n625), .A2(new_n627), .A3(KEYINPUT97), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n620), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n633), .A2(new_n427), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n619), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n277), .B1(new_n286), .B2(new_n287), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n604), .A2(new_n288), .A3(new_n359), .A4(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  XNOR2_X1  g456(.A(new_n417), .B(KEYINPUT98), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n643), .A2(new_n414), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n460), .A3(new_n427), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n607), .B2(new_n618), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n639), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NAND2_X1  g463(.A1(new_n358), .A2(new_n350), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n334), .A2(new_n342), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n340), .A2(KEYINPUT36), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n651), .B(new_n652), .Z(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n351), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n637), .A2(new_n288), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n658), .A2(new_n557), .A3(new_n461), .A4(new_n604), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT99), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  NAND2_X1  g476(.A1(new_n289), .A2(new_n296), .ZN(new_n663));
  INV_X1    g477(.A(new_n276), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n604), .A3(new_n655), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n425), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n421), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n644), .A2(new_n460), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n607), .B2(new_n618), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n666), .B1(new_n671), .B2(KEYINPUT100), .ZN(new_n672));
  INV_X1    g486(.A(new_n670), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n619), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XNOR2_X1  g492(.A(new_n669), .B(KEYINPUT39), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n604), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT40), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n290), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n261), .B1(new_n272), .B2(new_n254), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n277), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G472), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n663), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n462), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n620), .A2(new_n460), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n655), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(new_n680), .B2(new_n681), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT38), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n616), .B(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n688), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n214), .ZN(G45));
  NAND2_X1  g510(.A1(new_n595), .A2(KEYINPUT85), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n599), .A2(new_n600), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n603), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n558), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n297), .A2(new_n700), .A3(new_n656), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n620), .A2(new_n632), .A3(new_n669), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n701), .A2(new_n619), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  NAND2_X1  g519(.A1(new_n665), .A2(new_n359), .ZN(new_n706));
  INV_X1    g520(.A(G469), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n698), .B1(new_n707), .B2(new_n599), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n558), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n635), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n646), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  NOR4_X1   g530(.A1(new_n297), .A2(new_n656), .A3(new_n460), .A4(new_n428), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n710), .B1(new_n607), .B2(new_n618), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  NAND2_X1  g534(.A1(new_n273), .A2(new_n262), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n291), .A2(new_n282), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(G472), .A2(G902), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n636), .A2(G472), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n359), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT101), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT101), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n724), .A2(new_n727), .A3(new_n359), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n710), .A2(new_n426), .ZN(new_n730));
  INV_X1    g544(.A(new_n690), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT102), .B1(new_n619), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  AOI211_X1 g547(.A(new_n733), .B(new_n690), .C1(new_n607), .C2(new_n618), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n729), .B(new_n730), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT103), .B(G122), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G24));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n702), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n620), .A2(new_n632), .A3(KEYINPUT104), .A4(new_n669), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n724), .A2(new_n655), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n718), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  AOI21_X1  g559(.A(new_n559), .B1(new_n698), .B2(new_n595), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n614), .A2(new_n746), .A3(new_n615), .A4(new_n462), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n747), .A2(KEYINPUT105), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(KEYINPUT105), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n741), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n706), .A2(KEYINPUT106), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n361), .A2(new_n752), .ZN(new_n753));
  AND4_X1   g567(.A1(KEYINPUT42), .A2(new_n750), .A3(new_n751), .A4(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n706), .B1(new_n748), .B2(new_n749), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT42), .B1(new_n755), .B2(new_n742), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n223), .ZN(G33));
  XOR2_X1   g572(.A(new_n670), .B(KEYINPUT107), .Z(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n755), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  AND2_X1   g575(.A1(new_n657), .A2(new_n655), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n414), .A2(new_n417), .A3(new_n632), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(KEYINPUT43), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n766), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n762), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT109), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n616), .A2(new_n689), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n762), .A2(new_n769), .A3(new_n774), .A4(KEYINPUT44), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT110), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n770), .A2(new_n771), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n581), .B2(new_n593), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n592), .A2(new_n574), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n582), .ZN(new_n782));
  INV_X1    g596(.A(new_n580), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n574), .A3(new_n578), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(KEYINPUT45), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n780), .A2(new_n785), .A3(G469), .ZN(new_n786));
  NAND2_X1  g600(.A1(G469), .A2(G902), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(KEYINPUT46), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n698), .B1(new_n788), .B2(KEYINPUT46), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n558), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n778), .A2(new_n679), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n776), .B2(KEYINPUT110), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n777), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT111), .B(G137), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(G39));
  NAND4_X1  g611(.A1(new_n773), .A2(new_n297), .A3(new_n360), .A4(new_n703), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n792), .A2(KEYINPUT47), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n791), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n798), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(new_n310), .ZN(G42));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n459), .A2(new_n669), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n773), .A2(new_n644), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n804), .B1(new_n666), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n644), .A2(new_n805), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n701), .A2(KEYINPUT113), .A3(new_n773), .A4(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n807), .A2(new_n809), .B1(new_n750), .B2(new_n743), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n760), .B(new_n810), .C1(new_n754), .C2(new_n756), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n711), .B1(new_n635), .B2(new_n646), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n657), .A2(new_n360), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(new_n557), .A3(new_n604), .A4(new_n634), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n605), .A2(new_n659), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n816));
  INV_X1    g630(.A(new_n428), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n616), .A3(new_n460), .A4(new_n462), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n638), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n818), .A2(new_n816), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n819), .A2(new_n820), .B1(new_n717), .B2(new_n718), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n735), .A2(new_n812), .A3(new_n815), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n811), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n704), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n617), .B1(new_n616), .B2(new_n462), .ZN(new_n825));
  AOI211_X1 g639(.A(KEYINPUT96), .B(new_n689), .C1(new_n614), .C2(new_n615), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n731), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n733), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n619), .A2(KEYINPUT102), .A3(new_n731), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n656), .A2(new_n687), .A3(new_n669), .A4(new_n746), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n824), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n739), .A2(new_n655), .A3(new_n724), .A4(new_n740), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n710), .B(new_n833), .C1(new_n607), .C2(new_n618), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n672), .B2(new_n676), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n831), .B1(new_n732), .B2(new_n734), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n835), .A2(KEYINPUT52), .A3(new_n704), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n836), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  AOI211_X1 g654(.A(KEYINPUT114), .B(KEYINPUT52), .C1(new_n832), .C2(new_n835), .ZN(new_n841));
  OAI211_X1 g655(.A(KEYINPUT53), .B(new_n823), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n838), .A2(new_n704), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n619), .A2(KEYINPUT100), .A3(new_n673), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n701), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n671), .A2(KEYINPUT100), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n744), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n844), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n839), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n823), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n842), .A2(new_n843), .A3(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n751), .A2(new_n753), .ZN(new_n856));
  INV_X1    g670(.A(new_n710), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n422), .A2(new_n769), .A3(new_n857), .A4(new_n773), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT48), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n773), .A2(new_n857), .A3(new_n422), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n663), .A2(new_n359), .A3(new_n686), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n861), .A2(KEYINPUT116), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT116), .B1(new_n861), .B2(new_n862), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n633), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n729), .A2(new_n422), .A3(new_n769), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n718), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n419), .A2(new_n860), .A3(new_n865), .A4(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n694), .A2(new_n689), .A3(new_n857), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT50), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n867), .A2(KEYINPUT50), .A3(new_n870), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n873), .A2(new_n874), .B1(new_n743), .B2(new_n858), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n867), .A2(KEYINPUT115), .A3(new_n773), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n799), .B(new_n801), .C1(new_n558), .C2(new_n708), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n878));
  INV_X1    g692(.A(new_n773), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n878), .B1(new_n866), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n620), .A2(new_n632), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n863), .A2(new_n864), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n875), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n875), .A2(new_n881), .A3(KEYINPUT51), .A4(new_n883), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n869), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n851), .A2(new_n823), .A3(KEYINPUT53), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n823), .B1(new_n840), .B2(new_n841), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(new_n890), .B2(new_n853), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n855), .B(new_n888), .C1(new_n891), .C2(new_n843), .ZN(new_n892));
  OR2_X1    g706(.A1(G952), .A2(G953), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n862), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n763), .A2(new_n689), .A3(new_n559), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n708), .B(KEYINPUT49), .Z(new_n897));
  NAND4_X1  g711(.A1(new_n694), .A2(new_n895), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n894), .A2(KEYINPUT117), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(G75));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n531), .B(new_n523), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT118), .Z(new_n907));
  AND2_X1   g721(.A1(new_n842), .A2(new_n854), .ZN(new_n908));
  NAND2_X1  g722(.A1(G210), .A2(G902), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n904), .B(new_n907), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n337), .A2(G952), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n842), .A2(new_n854), .ZN(new_n913));
  INV_X1    g727(.A(new_n909), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT56), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n906), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n910), .B(new_n912), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT119), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n915), .A2(new_n916), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n910), .A4(new_n912), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n918), .A2(new_n921), .ZN(G51));
  XOR2_X1   g736(.A(new_n787), .B(KEYINPUT57), .Z(new_n923));
  NOR2_X1   g737(.A1(new_n908), .A2(new_n843), .ZN(new_n924));
  INV_X1    g738(.A(new_n855), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n597), .A2(new_n598), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OR3_X1    g742(.A1(new_n908), .A2(new_n277), .A3(new_n786), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n911), .B1(new_n928), .B2(new_n929), .ZN(G54));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n913), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n411), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n911), .B1(new_n932), .B2(new_n411), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n932), .A2(new_n931), .A3(new_n411), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(G60));
  XNOR2_X1  g751(.A(new_n626), .B(KEYINPUT59), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n851), .A2(new_n823), .A3(KEYINPUT53), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n856), .A2(KEYINPUT42), .A3(new_n750), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n755), .A2(new_n742), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT42), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI22_X1  g757(.A1(new_n940), .A2(new_n943), .B1(new_n755), .B2(new_n759), .ZN(new_n944));
  AND4_X1   g758(.A1(new_n735), .A2(new_n815), .A3(new_n812), .A4(new_n821), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n945), .A3(new_n810), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n839), .A2(new_n837), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n850), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n939), .B1(new_n950), .B2(KEYINPUT53), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT54), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n938), .B1(new_n952), .B2(new_n855), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n622), .A2(new_n624), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n912), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n938), .B1(new_n622), .B2(new_n624), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n924), .B2(new_n925), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(KEYINPUT121), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT121), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n959), .B(new_n956), .C1(new_n924), .C2(new_n925), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n955), .B1(new_n958), .B2(new_n960), .ZN(G63));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n962));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT122), .Z(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT60), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n348), .B1(new_n908), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n912), .ZN(new_n967));
  INV_X1    g781(.A(new_n653), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n908), .A2(new_n968), .A3(new_n965), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n962), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n969), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(KEYINPUT61), .A3(new_n912), .A4(new_n966), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(G66));
  OAI21_X1  g787(.A(G953), .B1(new_n423), .B2(new_n521), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT123), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n822), .B(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n974), .B1(new_n977), .B2(G953), .ZN(new_n978));
  OAI22_X1  g792(.A1(new_n610), .A2(new_n524), .B1(G898), .B2(new_n337), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(G69));
  AOI21_X1  g794(.A(new_n337), .B1(G227), .B2(G900), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT125), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n944), .B(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n802), .B1(new_n777), .B2(new_n794), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n835), .A2(new_n704), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n830), .A2(new_n856), .A3(new_n679), .A4(new_n792), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n984), .A2(new_n986), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n337), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n667), .A2(G953), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT126), .B1(new_n992), .B2(new_n993), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n244), .A2(new_n246), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(KEYINPUT30), .B2(new_n244), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(new_n390), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n996), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  OR3_X1    g816(.A1(new_n985), .A2(KEYINPUT62), .A3(new_n695), .ZN(new_n1003));
  OAI21_X1  g817(.A(KEYINPUT62), .B1(new_n985), .B2(new_n695), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n414), .A2(new_n460), .A3(new_n417), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1006), .A2(new_n633), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n361), .A2(new_n773), .A3(new_n680), .A4(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1003), .A2(new_n1004), .A3(new_n1008), .A4(new_n984), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1002), .B1(new_n1009), .B2(new_n337), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n981), .B1(new_n1001), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n981), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1010), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n997), .A2(new_n1000), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1012), .B(new_n1013), .C1(new_n1014), .C2(new_n996), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1011), .A2(new_n1015), .ZN(G72));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  OAI21_X1  g832(.A(new_n1018), .B1(new_n1009), .B2(new_n976), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1019), .A2(new_n261), .A3(new_n255), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1018), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n983), .A2(new_n991), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1021), .B1(new_n1022), .B2(new_n977), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n247), .A2(new_n254), .A3(new_n262), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n1020), .B(new_n912), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1021), .B1(new_n263), .B2(new_n290), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1025), .B1(new_n951), .B2(new_n1026), .ZN(G57));
endmodule


