//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  AND2_X1   g0010(.A1(new_n210), .A2(KEYINPUT65), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(KEYINPUT65), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n202), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n201), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n207), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n203), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR4_X1   g0028(.A1(new_n211), .A2(new_n212), .A3(new_n224), .A4(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(G226), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND2_X1  g0045(.A1(G33), .A2(G97), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT68), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n249), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G226), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G1698), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n246), .B1(new_n253), .B2(new_n254), .C1(new_n256), .C2(new_n219), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT13), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n259), .A2(G274), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n266), .A2(G238), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n261), .A2(new_n262), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n262), .B1(new_n261), .B2(new_n271), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G190), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G77), .ZN(new_n279));
  INV_X1    g0079(.A(G50), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n279), .B1(new_n226), .B2(G68), .C1(new_n280), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n227), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(KEYINPUT11), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G13), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(new_n226), .A3(G1), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n202), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT12), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n288), .A2(new_n285), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n263), .A2(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G68), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n286), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT11), .B1(new_n283), .B2(new_n285), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(G200), .B1(new_n273), .B2(new_n274), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n276), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n296), .ZN(new_n300));
  OAI21_X1  g0100(.A(G169), .B1(new_n273), .B2(new_n274), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT14), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n275), .A2(G179), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT14), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(G169), .C1(new_n273), .C2(new_n274), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n299), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n292), .A2(G50), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n291), .A2(new_n309), .B1(new_n280), .B2(new_n288), .ZN(new_n310));
  OAI21_X1  g0110(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT69), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n314), .A2(new_n278), .B1(G150), .B2(new_n281), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n285), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n310), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT9), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n266), .A2(G226), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n270), .A2(new_n259), .A3(G274), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT67), .ZN(new_n324));
  INV_X1    g0124(.A(G223), .ZN(new_n325));
  INV_X1    g0125(.A(G77), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n256), .A2(new_n325), .B1(new_n326), .B2(new_n255), .ZN(new_n327));
  INV_X1    g0127(.A(G222), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n253), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n260), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT67), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n321), .A2(new_n331), .A3(new_n322), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n324), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G200), .ZN(new_n334));
  OAI211_X1 g0134(.A(KEYINPUT9), .B(new_n310), .C1(new_n316), .C2(new_n317), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n324), .A2(new_n330), .A3(G190), .A4(new_n332), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n320), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT10), .ZN(new_n338));
  INV_X1    g0138(.A(new_n333), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n318), .B1(new_n339), .B2(G169), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT70), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n341), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n342), .B(new_n343), .C1(G179), .C2(new_n333), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n251), .A2(new_n252), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G107), .ZN(new_n346));
  OAI221_X1 g0146(.A(new_n346), .B1(new_n253), .B2(new_n219), .C1(new_n214), .C2(new_n256), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n260), .ZN(new_n348));
  INV_X1    g0148(.A(G244), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n322), .B1(new_n349), .B2(new_n265), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT71), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n350), .A2(KEYINPUT71), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  OR2_X1    g0153(.A1(new_n353), .A2(G179), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n291), .A2(G77), .A3(new_n292), .ZN(new_n355));
  INV_X1    g0155(.A(new_n288), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n355), .B1(G77), .B2(new_n356), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT15), .B(G87), .Z(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n278), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n359), .B1(new_n226), .B2(new_n326), .C1(new_n282), .C2(new_n313), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n357), .B1(new_n360), .B2(new_n285), .ZN(new_n361));
  INV_X1    g0161(.A(G169), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n361), .B1(new_n353), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n354), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n353), .A2(G200), .ZN(new_n365));
  INV_X1    g0165(.A(G190), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n365), .B(new_n361), .C1(new_n366), .C2(new_n353), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n338), .A2(new_n344), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT16), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n255), .B2(G20), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n345), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n202), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n201), .A2(new_n202), .ZN(new_n376));
  NOR2_X1   g0176(.A1(G58), .A2(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(G20), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n281), .A2(G159), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n371), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n345), .B2(new_n226), .ZN(new_n382));
  NOR4_X1   g0182(.A1(new_n251), .A2(new_n252), .A3(new_n372), .A4(G20), .ZN(new_n383));
  OAI21_X1  g0183(.A(G68), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n380), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(KEYINPUT16), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n386), .A3(new_n285), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n313), .B1(new_n263), .B2(G20), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(new_n291), .B1(new_n288), .B2(new_n313), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(G226), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n391), .B(new_n392), .C1(new_n253), .C2(new_n325), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n260), .ZN(new_n394));
  INV_X1    g0194(.A(G179), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n322), .B1(new_n265), .B2(new_n219), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(new_n393), .B2(new_n260), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n399), .A2(G169), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n390), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT18), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n394), .A2(new_n366), .A3(new_n397), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G200), .B2(new_n399), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n404), .A2(new_n387), .A3(new_n389), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT17), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n398), .B1(G169), .B2(new_n399), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n387), .B2(new_n389), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n404), .A2(new_n387), .A3(new_n389), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n402), .A2(new_n406), .A3(new_n410), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT72), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n414), .A2(KEYINPUT72), .ZN(new_n416));
  AND4_X1   g0216(.A1(new_n307), .A2(new_n370), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT19), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT73), .B(G97), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n226), .A2(G33), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G87), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n423), .A3(new_n215), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n226), .B1(new_n246), .B2(new_n419), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n226), .B(G68), .C1(new_n251), .C2(new_n252), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n427), .A2(KEYINPUT77), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(KEYINPUT77), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n422), .B(new_n426), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n285), .ZN(new_n431));
  INV_X1    g0231(.A(new_n358), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n288), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n263), .A2(G33), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n291), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n358), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n431), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT78), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT76), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G116), .ZN(new_n442));
  OAI211_X1 g0242(.A(G244), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n442), .B(new_n443), .C1(new_n253), .C2(new_n214), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n260), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n263), .A2(G45), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n446), .A2(G250), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n267), .A2(new_n447), .B1(new_n448), .B2(new_n259), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n441), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n445), .A2(new_n441), .A3(new_n449), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n362), .A3(new_n452), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n445), .A2(new_n441), .A3(new_n449), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n395), .B1(new_n454), .B2(new_n450), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n431), .A2(KEYINPUT78), .A3(new_n433), .A4(new_n437), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n440), .A2(new_n453), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(G190), .B1(new_n454), .B2(new_n450), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n436), .A2(G87), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n431), .A2(new_n433), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n451), .A2(new_n452), .ZN(new_n461));
  INV_X1    g0261(.A(G200), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n458), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT82), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n256), .B2(new_n221), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n255), .A2(KEYINPUT82), .A3(G257), .A4(G1698), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n249), .A2(new_n250), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G250), .A3(new_n255), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G294), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n466), .A2(new_n467), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n260), .ZN(new_n472));
  OR2_X1    g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n446), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n267), .A2(new_n475), .ZN(new_n476));
  OR2_X1    g0276(.A1(new_n475), .A2(new_n260), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(new_n216), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n472), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n362), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n471), .B2(new_n260), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n395), .A3(new_n476), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n442), .A2(G20), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT23), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n226), .B2(G107), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n215), .A2(KEYINPUT23), .A3(G20), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n255), .A2(new_n226), .A3(G87), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n489), .A2(KEYINPUT22), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(KEYINPUT22), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT24), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT24), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n494), .B(new_n488), .C1(new_n490), .C2(new_n491), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n317), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n288), .A2(KEYINPUT25), .A3(new_n215), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT25), .B1(new_n288), .B2(new_n215), .ZN(new_n499));
  OAI22_X1  g0299(.A1(new_n435), .A2(new_n215), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n481), .B(new_n483), .C1(new_n496), .C2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n464), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n477), .A2(new_n221), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n253), .B2(new_n349), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT75), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(KEYINPUT75), .B(new_n505), .C1(new_n253), .C2(new_n349), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n345), .A2(new_n248), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n468), .A2(KEYINPUT4), .A3(G244), .A4(new_n255), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n508), .A2(new_n509), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n504), .B1(new_n513), .B2(new_n260), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(new_n366), .A3(new_n476), .ZN(new_n515));
  INV_X1    g0315(.A(new_n476), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n516), .B(new_n504), .C1(new_n513), .C2(new_n260), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(G200), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n356), .A2(G97), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n436), .B2(G97), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(G107), .B1(new_n382), .B2(new_n383), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT74), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT74), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n524), .B(G107), .C1(new_n382), .C2(new_n383), .ZN(new_n525));
  XOR2_X1   g0325(.A(G97), .B(G107), .Z(new_n526));
  NAND2_X1  g0326(.A1(new_n215), .A2(KEYINPUT6), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n526), .A2(KEYINPUT6), .B1(new_n420), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(G20), .B1(G77), .B2(new_n281), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n523), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n521), .B1(new_n530), .B2(new_n285), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n517), .B2(new_n395), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n514), .A2(new_n476), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n362), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n518), .A2(new_n531), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n356), .A2(G116), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n436), .B2(G116), .ZN(new_n537));
  AOI21_X1  g0337(.A(G20), .B1(G33), .B2(G283), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n420), .B2(G33), .ZN(new_n539));
  INV_X1    g0339(.A(G116), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G20), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n285), .A2(KEYINPUT79), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT79), .B1(new_n285), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT20), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n545), .A2(KEYINPUT80), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(KEYINPUT80), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n285), .A2(new_n541), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT79), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n285), .A2(KEYINPUT79), .A3(new_n541), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n553), .A2(KEYINPUT80), .A3(new_n545), .A4(new_n539), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n537), .A2(new_n548), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n345), .A2(G303), .ZN(new_n556));
  OAI211_X1 g0356(.A(G264), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n556), .B(new_n557), .C1(new_n253), .C2(new_n221), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n260), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n475), .A2(new_n260), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n560), .A2(G270), .B1(new_n267), .B2(new_n475), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n362), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT21), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n555), .A2(KEYINPUT21), .A3(new_n562), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n559), .A2(new_n561), .A3(G179), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT81), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n555), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n568), .B1(new_n555), .B2(new_n567), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n565), .B(new_n566), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n559), .A2(new_n561), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n366), .ZN(new_n573));
  AOI211_X1 g0373(.A(new_n555), .B(new_n573), .C1(G200), .C2(new_n572), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n472), .A2(new_n366), .A3(new_n476), .A4(new_n479), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT83), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n480), .A2(new_n462), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT83), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n482), .A2(new_n579), .A3(new_n366), .A4(new_n476), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n496), .A2(new_n500), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n503), .A2(new_n535), .A3(new_n575), .A4(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n418), .A2(new_n584), .ZN(G372));
  AND2_X1   g0385(.A1(new_n402), .A2(new_n410), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n306), .A2(new_n300), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n299), .B2(new_n364), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n406), .A2(new_n413), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n338), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n344), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT84), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n444), .A2(new_n595), .A3(new_n260), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n444), .B2(new_n260), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n449), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n362), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(new_n455), .A3(new_n438), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(G200), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n458), .A2(new_n602), .A3(new_n460), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n600), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n514), .A2(new_n395), .A3(new_n476), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n530), .A2(new_n285), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n520), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n607), .C1(new_n517), .C2(G169), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT26), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n601), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT26), .B1(new_n464), .B2(new_n608), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT85), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n571), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n555), .A2(new_n567), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT81), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n555), .A2(new_n567), .A3(new_n568), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(KEYINPUT85), .A3(new_n565), .A4(new_n566), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n502), .B1(new_n614), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n603), .A2(new_n600), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n518), .A2(new_n531), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n621), .A2(new_n622), .A3(new_n583), .A4(new_n608), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n611), .B(new_n612), .C1(new_n620), .C2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n594), .B1(new_n418), .B2(new_n625), .ZN(G369));
  NAND3_X1  g0426(.A1(new_n263), .A2(new_n226), .A3(G13), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(G213), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(G343), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n555), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n575), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n614), .A2(new_n619), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(new_n633), .ZN(new_n636));
  XOR2_X1   g0436(.A(new_n636), .B(KEYINPUT86), .Z(new_n637));
  INV_X1    g0437(.A(new_n632), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n582), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n582), .B2(new_n581), .ZN(new_n640));
  MUX2_X1   g0440(.A(new_n632), .B(new_n640), .S(new_n501), .Z(new_n641));
  NAND3_X1  g0441(.A1(new_n637), .A2(G330), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n502), .A2(new_n638), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n640), .A2(new_n571), .A3(new_n501), .A4(new_n638), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(G399));
  INV_X1    g0445(.A(new_n208), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(G41), .ZN(new_n647));
  INV_X1    g0447(.A(new_n225), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n424), .A2(G116), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G1), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT28), .ZN(new_n653));
  INV_X1    g0453(.A(G330), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n514), .A2(new_n567), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT87), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n461), .B2(new_n482), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n482), .B(new_n656), .C1(new_n454), .C2(new_n450), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI211_X1 g0459(.A(KEYINPUT30), .B(new_n655), .C1(new_n657), .C2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n655), .B1(new_n657), .B2(new_n659), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT30), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n480), .A2(new_n395), .A3(new_n572), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n533), .A3(new_n598), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT88), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n661), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n666), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n663), .B2(new_n662), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT88), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT31), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n638), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n584), .A2(KEYINPUT31), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n664), .A2(new_n674), .A3(new_n660), .A4(new_n666), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n632), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n654), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n502), .A2(new_n571), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n623), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n605), .A2(new_n607), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n517), .A2(G169), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(new_n610), .A3(new_n463), .A4(new_n457), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT26), .B1(new_n604), .B2(new_n608), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n600), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n638), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT29), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n624), .A2(new_n638), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n691), .B1(KEYINPUT29), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n681), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n653), .B1(new_n694), .B2(G1), .ZN(G364));
  AND2_X1   g0495(.A1(new_n637), .A2(G330), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n287), .A2(G20), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n263), .B1(new_n697), .B2(G45), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n647), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(G330), .B2(new_n637), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n208), .A2(G355), .A3(new_n255), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(G116), .B2(new_n208), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n208), .A2(new_n345), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n269), .B2(new_n648), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n241), .A2(new_n269), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(G13), .A2(G33), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G20), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n227), .B1(G20), .B2(new_n362), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n700), .B1(new_n708), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n226), .A2(G179), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(G190), .A3(G200), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(new_n366), .A3(G200), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n423), .A2(new_n717), .B1(new_n718), .B2(new_n215), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n226), .A2(new_n395), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G200), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n366), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n719), .B1(G50), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G190), .A2(G200), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n716), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G159), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT32), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n720), .A2(G190), .A3(new_n462), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n255), .B1(new_n729), .B2(new_n201), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n720), .A2(new_n724), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n730), .B1(G77), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n366), .A2(G179), .A3(G200), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n226), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n721), .A2(G190), .ZN(new_n737));
  AOI22_X1  g0537(.A1(G97), .A2(new_n736), .B1(new_n737), .B2(G68), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n723), .A2(new_n728), .A3(new_n733), .A4(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G322), .ZN(new_n740));
  INV_X1    g0540(.A(G311), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n729), .A2(new_n740), .B1(new_n731), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n725), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n255), .B(new_n742), .C1(G329), .C2(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(G294), .A2(new_n736), .B1(new_n722), .B2(G326), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT33), .B(G317), .ZN(new_n746));
  INV_X1    g0546(.A(new_n718), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n737), .A2(new_n746), .B1(new_n747), .B2(G283), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n744), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n717), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n750), .A2(KEYINPUT89), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(KEYINPUT89), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G303), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n739), .B1(new_n749), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n715), .B1(new_n756), .B2(new_n712), .ZN(new_n757));
  INV_X1    g0557(.A(new_n711), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n757), .B1(new_n636), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n702), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(G396));
  NOR2_X1   g0561(.A1(new_n368), .A2(new_n632), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n620), .A2(new_n623), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n609), .A2(new_n610), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(new_n600), .A3(new_n612), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n367), .B1(new_n361), .B2(new_n638), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n364), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n364), .A2(new_n632), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT90), .Z(new_n773));
  AOI21_X1  g0573(.A(new_n767), .B1(new_n692), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n681), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT91), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n700), .B(new_n777), .C1(new_n681), .C2(new_n774), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n776), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n700), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n712), .A2(new_n709), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(new_n326), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n712), .ZN(new_n784));
  INV_X1    g0584(.A(new_n729), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n785), .A2(G294), .B1(new_n743), .B2(G311), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n786), .B(new_n345), .C1(new_n540), .C2(new_n731), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n737), .A2(G283), .B1(new_n747), .B2(G87), .ZN(new_n788));
  INV_X1    g0588(.A(new_n722), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n788), .B1(new_n220), .B2(new_n735), .C1(new_n754), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n753), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n787), .B(new_n790), .C1(G107), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n718), .A2(new_n202), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n345), .B(new_n793), .C1(G132), .C2(new_n743), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n201), .B2(new_n735), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n785), .A2(G143), .B1(new_n732), .B2(G159), .ZN(new_n796));
  INV_X1    g0596(.A(G137), .ZN(new_n797));
  INV_X1    g0597(.A(G150), .ZN(new_n798));
  INV_X1    g0598(.A(new_n737), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n796), .B1(new_n789), .B2(new_n797), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT34), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n795), .B(new_n802), .C1(G50), .C2(new_n791), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n792), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n772), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n783), .B1(new_n784), .B2(new_n805), .C1(new_n806), .C2(new_n710), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n780), .A2(new_n807), .ZN(G384));
  NOR2_X1   g0608(.A1(new_n697), .A2(new_n263), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n306), .A2(new_n300), .A3(new_n638), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n389), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n384), .A2(new_n385), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n317), .B1(new_n813), .B2(new_n371), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(new_n814), .B2(new_n386), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n630), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n414), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n411), .B1(new_n815), .B2(new_n407), .ZN(new_n818));
  OAI21_X1  g0618(.A(KEYINPUT37), .B1(new_n818), .B2(new_n816), .ZN(new_n819));
  INV_X1    g0619(.A(new_n630), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n390), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT37), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n401), .A2(new_n821), .A3(new_n822), .A4(new_n411), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n817), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT38), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n817), .A2(KEYINPUT38), .A3(new_n824), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT39), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n828), .B(KEYINPUT96), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n816), .B1(new_n818), .B2(KEYINPUT93), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT93), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n401), .A2(new_n835), .A3(new_n411), .ZN(new_n836));
  AOI211_X1 g0636(.A(KEYINPUT94), .B(new_n822), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n823), .A2(KEYINPUT94), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT93), .B1(new_n405), .B2(new_n408), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n839), .A2(new_n836), .A3(new_n821), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n838), .B1(new_n840), .B2(KEYINPUT37), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT95), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT94), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n840), .A2(new_n843), .A3(KEYINPUT37), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT95), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n822), .B1(new_n834), .B2(new_n836), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n838), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n842), .A2(new_n847), .A3(new_n817), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n833), .B1(new_n826), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n811), .B(new_n832), .C1(new_n849), .C2(KEYINPUT39), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n300), .A2(new_n632), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n588), .A2(new_n298), .A3(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n300), .B(new_n632), .C1(new_n299), .C2(new_n306), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n766), .B2(new_n771), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n855), .A2(new_n829), .B1(new_n587), .B2(new_n630), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n593), .B1(new_n693), .B2(new_n417), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n848), .A2(new_n826), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n828), .B(KEYINPUT96), .Z(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n675), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n671), .B2(new_n660), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n677), .B2(new_n679), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n852), .A2(new_n853), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n806), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT97), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n772), .B1(new_n852), .B2(new_n853), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT97), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n584), .A2(KEYINPUT31), .B1(new_n678), .B2(new_n632), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n869), .B(new_n870), .C1(new_n871), .C2(new_n864), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n862), .A2(KEYINPUT40), .A3(new_n868), .A4(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n864), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n680), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n829), .A3(new_n869), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n875), .A2(new_n417), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n654), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n809), .B1(new_n859), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n859), .B2(new_n882), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n227), .A2(new_n226), .A3(new_n540), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT36), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n225), .A2(new_n326), .A3(new_n376), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n890), .A2(KEYINPUT92), .B1(new_n280), .B2(G68), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(KEYINPUT92), .B2(new_n890), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(G1), .A3(new_n287), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n884), .A2(new_n889), .A3(new_n893), .ZN(G367));
  INV_X1    g0694(.A(new_n237), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n713), .B1(new_n208), .B2(new_n432), .C1(new_n895), .C2(new_n705), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n700), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n255), .B1(new_n743), .B2(G317), .ZN(new_n898));
  INV_X1    g0698(.A(G283), .ZN(new_n899));
  OAI221_X1 g0699(.A(new_n898), .B1(new_n899), .B2(new_n731), .C1(new_n754), .C2(new_n729), .ZN(new_n900));
  INV_X1    g0700(.A(G294), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n799), .A2(new_n901), .B1(new_n789), .B2(new_n741), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n735), .A2(new_n215), .B1(new_n718), .B2(new_n420), .ZN(new_n903));
  XOR2_X1   g0703(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n750), .B2(G116), .ZN(new_n905));
  NOR4_X1   g0705(.A1(new_n900), .A2(new_n902), .A3(new_n903), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n791), .A2(KEYINPUT46), .A3(G116), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n255), .B1(new_n725), .B2(new_n797), .C1(new_n729), .C2(new_n798), .ZN(new_n909));
  INV_X1    g0709(.A(G143), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n789), .A2(new_n910), .B1(new_n717), .B2(new_n201), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n735), .A2(new_n202), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n718), .A2(new_n326), .ZN(new_n913));
  OR4_X1    g0713(.A1(new_n909), .A2(new_n911), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n737), .A2(G159), .B1(new_n732), .B2(G50), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT108), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n908), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT47), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n897), .B1(new_n918), .B2(new_n712), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n460), .A2(new_n638), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n604), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n601), .A2(new_n920), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n711), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT105), .ZN(new_n925));
  INV_X1    g0725(.A(new_n694), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n571), .A2(new_n638), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n641), .B(new_n927), .Z(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n696), .B2(KEYINPUT104), .ZN(new_n929));
  INV_X1    g0729(.A(new_n928), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n637), .A2(G330), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT104), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n622), .B(new_n608), .C1(new_n531), .C2(new_n638), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n686), .A2(new_n632), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n938));
  NAND4_X1  g0738(.A1(new_n937), .A2(new_n644), .A3(new_n643), .A4(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n938), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n644), .A2(new_n643), .ZN(new_n941));
  INV_X1    g0741(.A(new_n937), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND4_X1   g0743(.A1(KEYINPUT44), .A2(new_n941), .A3(new_n935), .A4(new_n936), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT44), .B1(new_n941), .B2(new_n942), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n939), .B(new_n943), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(new_n642), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n926), .B1(new_n934), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n647), .B(new_n949), .Z(new_n950));
  OAI21_X1  g0750(.A(new_n925), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n946), .B(new_n642), .Z(new_n952));
  NAND2_X1  g0752(.A1(new_n929), .A2(new_n933), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n694), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n950), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(KEYINPUT105), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n699), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n921), .A2(new_n922), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT98), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(KEYINPUT99), .B(KEYINPUT101), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n608), .B1(new_n935), .B2(new_n501), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n638), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n942), .A2(new_n644), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT42), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT100), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n967), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT100), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n971), .B(new_n965), .C1(new_n966), .C2(new_n967), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n637), .A2(G330), .A3(new_n641), .A4(new_n937), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n974), .B1(new_n973), .B2(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n963), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n978), .ZN(new_n980));
  INV_X1    g0780(.A(new_n963), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(new_n976), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n962), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n979), .A2(new_n982), .A3(new_n962), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT106), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n957), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n948), .A2(new_n925), .A3(new_n950), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT105), .B1(new_n954), .B2(new_n955), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n698), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n985), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(new_n983), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT106), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n924), .B1(new_n988), .B2(new_n994), .ZN(G387));
  NAND2_X1  g0795(.A1(new_n934), .A2(new_n694), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n953), .A2(new_n926), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n647), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n234), .A2(G45), .A3(new_n345), .ZN(new_n999));
  OAI21_X1  g0799(.A(KEYINPUT50), .B1(new_n313), .B2(G50), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n1000), .B(new_n269), .C1(new_n202), .C2(new_n326), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n313), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n345), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n650), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n646), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n713), .B1(new_n208), .B2(new_n215), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n700), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n729), .A2(new_n280), .B1(new_n725), .B2(new_n798), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n345), .B(new_n1008), .C1(G68), .C2(new_n732), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n750), .A2(G77), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n737), .A2(new_n314), .B1(new_n747), .B2(G97), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n358), .A2(new_n736), .B1(new_n722), .B2(G159), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n255), .B1(new_n743), .B2(G326), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n735), .A2(new_n899), .B1(new_n717), .B2(new_n901), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n785), .A2(G317), .B1(new_n732), .B2(G303), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n789), .B2(new_n740), .C1(new_n741), .C2(new_n799), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT48), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1018), .B2(new_n1017), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT49), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1014), .B1(new_n540), .B2(new_n718), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1013), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1007), .B1(new_n1024), .B2(new_n712), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n641), .B2(new_n758), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n998), .B(new_n1026), .C1(new_n698), .C2(new_n953), .ZN(G393));
  NAND2_X1  g0827(.A1(new_n996), .A2(new_n952), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n934), .A2(new_n694), .A3(new_n947), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n647), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n942), .A2(new_n711), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n713), .B1(new_n208), .B2(new_n420), .C1(new_n705), .C2(new_n244), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n700), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n789), .A2(new_n798), .B1(new_n726), .B2(new_n729), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT51), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n255), .B1(new_n725), .B2(new_n910), .C1(new_n313), .C2(new_n731), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n737), .A2(G50), .B1(new_n747), .B2(G87), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n735), .A2(new_n326), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G68), .B2(new_n750), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT109), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n345), .B1(new_n731), .B2(new_n901), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n799), .A2(new_n754), .B1(new_n540), .B2(new_n735), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(G107), .C2(new_n747), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G317), .A2(new_n722), .B1(new_n785), .B2(G311), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT52), .Z(new_n1047));
  AOI22_X1  g0847(.A1(new_n750), .A2(G283), .B1(new_n743), .B2(G322), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1048), .A2(KEYINPUT110), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(KEYINPUT110), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1045), .A2(new_n1047), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1041), .A2(KEYINPUT109), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1042), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1033), .B1(new_n1053), .B2(new_n712), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n947), .A2(new_n699), .B1(new_n1031), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1030), .A2(new_n1055), .ZN(G390));
  AOI21_X1  g0856(.A(new_n831), .B1(new_n862), .B2(new_n830), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1057), .A2(new_n710), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n781), .B1(new_n313), .B2(new_n782), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n737), .A2(G107), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n420), .B2(new_n731), .C1(new_n789), .C2(new_n899), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT116), .Z(new_n1062));
  NOR2_X1   g0862(.A1(new_n753), .A2(new_n423), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n345), .B1(new_n725), .B2(new_n901), .C1(new_n729), .C2(new_n540), .ZN(new_n1064));
  NOR4_X1   g0864(.A1(new_n1063), .A2(new_n793), .A3(new_n1039), .A4(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(KEYINPUT54), .B(G143), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n737), .A2(G137), .B1(new_n732), .B2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT115), .Z(new_n1069));
  AOI22_X1  g0869(.A1(G159), .A2(new_n736), .B1(new_n722), .B2(G128), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n280), .B2(new_n718), .ZN(new_n1071));
  INV_X1    g0871(.A(G125), .ZN(new_n1072));
  INV_X1    g0872(.A(G132), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n255), .B1(new_n725), .B2(new_n1072), .C1(new_n729), .C2(new_n1073), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n717), .A2(KEYINPUT53), .A3(new_n798), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT53), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n750), .B2(G150), .ZN(new_n1077));
  NOR4_X1   g0877(.A1(new_n1071), .A2(new_n1074), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1062), .A2(new_n1065), .B1(new_n1069), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1059), .B1(new_n1079), .B2(new_n784), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1058), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n865), .A2(new_n867), .A3(new_n654), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT112), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n855), .B2(new_n811), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n770), .B1(new_n624), .B2(new_n762), .ZN(new_n1086));
  OAI211_X1 g0886(.A(KEYINPUT112), .B(new_n810), .C1(new_n1086), .C2(new_n854), .ZN(new_n1087));
  AOI21_X1  g0887(.A(KEYINPUT39), .B1(new_n860), .B2(new_n861), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1085), .B(new_n1087), .C1(new_n1088), .C2(new_n831), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n638), .B(new_n769), .C1(new_n683), .C2(new_n689), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT111), .B1(new_n1090), .B2(new_n771), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(KEYINPUT111), .A3(new_n771), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1092), .A2(new_n866), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n811), .B1(new_n860), .B2(new_n861), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1083), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT113), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1057), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n681), .A2(new_n806), .A3(new_n866), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n844), .B1(new_n846), .B2(new_n838), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1102), .A2(KEYINPUT95), .B1(new_n414), .B2(new_n816), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT38), .B1(new_n1103), .B2(new_n847), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n810), .B1(new_n1104), .B2(new_n833), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1090), .A2(KEYINPUT111), .A3(new_n771), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n1106), .A2(new_n1091), .A3(new_n854), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1101), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1098), .B1(new_n1100), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n863), .B1(new_n669), .B2(new_n672), .ZN(new_n1110));
  OAI21_X1  g0910(.A(G330), .B1(new_n1110), .B2(new_n871), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1111), .A2(new_n772), .A3(new_n854), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1113), .A2(new_n1089), .A3(KEYINPUT113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1097), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1081), .B1(new_n1115), .B2(new_n699), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n875), .A2(new_n417), .A3(G330), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT114), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n875), .A2(new_n417), .A3(KEYINPUT114), .A4(G330), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n858), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n866), .B1(new_n681), .B2(new_n806), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1123), .A2(new_n1082), .B1(new_n767), .B2(new_n770), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n865), .A2(new_n773), .A3(new_n654), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1101), .B(new_n1125), .C1(new_n866), .C2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1122), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n647), .B1(new_n1115), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1096), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1082), .B1(new_n1100), .B2(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1113), .A2(new_n1089), .A3(KEYINPUT113), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT113), .B1(new_n1113), .B2(new_n1089), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1128), .B(new_n1131), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1116), .B1(new_n1129), .B2(new_n1135), .ZN(G378));
  INV_X1    g0936(.A(new_n1122), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n868), .A2(KEYINPUT40), .A3(new_n872), .ZN(new_n1138));
  OAI211_X1 g0938(.A(G330), .B(new_n878), .C1(new_n1138), .C2(new_n849), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n338), .A2(new_n344), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n318), .A2(new_n820), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1142), .B(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n873), .A2(G330), .A3(new_n878), .A4(new_n1144), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n857), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n857), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1134), .A2(new_n1137), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1152), .A2(KEYINPUT57), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1122), .B1(new_n1115), .B2(new_n1128), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1146), .A2(new_n857), .A3(new_n1147), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n857), .B1(new_n1147), .B2(new_n1146), .ZN(new_n1156));
  OAI21_X1  g0956(.A(KEYINPUT57), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT120), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT120), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1151), .A2(new_n1148), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(KEYINPUT57), .A4(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1153), .A2(new_n1158), .A3(new_n647), .A4(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n698), .B1(new_n1151), .B2(new_n1148), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n799), .A2(new_n1073), .B1(new_n789), .B2(new_n1072), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n785), .A2(G128), .B1(new_n732), .B2(G137), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n717), .B2(new_n1066), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(G150), .C2(new_n736), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n747), .A2(G159), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G33), .B(G41), .C1(new_n743), .C2(G124), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n789), .A2(new_n540), .B1(new_n718), .B2(new_n201), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G97), .B2(new_n737), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n345), .A2(new_n268), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G283), .B2(new_n743), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n785), .A2(G107), .B1(new_n732), .B2(new_n358), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n912), .B1(G77), .B2(new_n750), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1178), .B(new_n280), .C1(G33), .C2(G41), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1175), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n712), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT118), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n781), .B(new_n1189), .C1(new_n280), .C2(new_n782), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1145), .A2(new_n709), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1164), .A2(new_n1165), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n699), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT119), .B1(new_n1195), .B2(new_n1192), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1163), .A2(new_n1197), .ZN(G375));
  INV_X1    g0998(.A(new_n1128), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1122), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(new_n955), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n698), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n854), .A2(new_n709), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n712), .A2(G68), .A3(new_n709), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n791), .A2(G159), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n729), .A2(new_n797), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n255), .B1(new_n731), .B2(new_n798), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G128), .C2(new_n743), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n736), .A2(G50), .B1(new_n747), .B2(G58), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G132), .A2(new_n722), .B1(new_n737), .B2(new_n1067), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1205), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n791), .A2(G97), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n729), .A2(new_n899), .B1(new_n725), .B2(new_n754), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G107), .B2(new_n732), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n737), .A2(G116), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n358), .A2(new_n736), .B1(new_n722), .B2(G294), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n913), .A2(new_n255), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT121), .Z(new_n1219));
  OAI21_X1  g1019(.A(new_n1211), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n781), .B(new_n1204), .C1(new_n1220), .C2(new_n712), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1202), .B1(new_n1203), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1201), .A2(new_n1222), .ZN(G381));
  INV_X1    g1023(.A(G390), .ZN(new_n1224));
  INV_X1    g1024(.A(G384), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  OR4_X1    g1026(.A1(G396), .A2(new_n1226), .A3(G393), .A4(G381), .ZN(new_n1227));
  OR4_X1    g1027(.A1(G387), .A2(new_n1227), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1028(.A(G378), .ZN(new_n1229));
  INV_X1    g1029(.A(G213), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(G343), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G407), .B(G213), .C1(G375), .C2(new_n1232), .ZN(G409));
  OAI21_X1  g1033(.A(new_n987), .B1(new_n957), .B2(new_n986), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n991), .A2(new_n993), .A3(KEYINPUT106), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G390), .B1(new_n1236), .B2(new_n924), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n924), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n1238), .B(new_n1224), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(G393), .B(new_n760), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1237), .A2(new_n1239), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G387), .A2(new_n1224), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1236), .A2(new_n924), .A3(G390), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1240), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT123), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1200), .A2(new_n1249), .A3(KEYINPUT60), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT60), .B1(new_n1200), .B2(new_n1249), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n647), .B(new_n1199), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1222), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1225), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(G384), .A3(new_n1222), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1231), .A2(G2897), .ZN(new_n1257));
  OR3_X1    g1057(.A1(new_n1256), .A2(KEYINPUT124), .A3(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1256), .B2(KEYINPUT124), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1256), .A2(KEYINPUT124), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1164), .B(new_n1193), .C1(new_n1152), .C2(new_n955), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(G378), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1158), .A2(new_n1162), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n647), .B1(new_n1152), .B2(KEYINPUT57), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G378), .B(new_n1197), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT122), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT122), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1163), .A2(new_n1268), .A3(G378), .A4(new_n1197), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1263), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1261), .B1(new_n1270), .B2(new_n1231), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1270), .A2(new_n1231), .A3(new_n1256), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1248), .B(new_n1271), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1263), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1231), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1279), .A2(KEYINPUT62), .A3(new_n1256), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1247), .B1(new_n1274), .B2(new_n1280), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1271), .A2(new_n1248), .A3(new_n1246), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1279), .B2(new_n1256), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1256), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1277), .A2(KEYINPUT63), .A3(new_n1278), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT125), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1272), .A2(new_n1288), .A3(KEYINPUT63), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1282), .A2(new_n1284), .A3(new_n1287), .A4(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1281), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT126), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1281), .A2(new_n1290), .A3(KEYINPUT126), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(G405));
  NAND2_X1  g1095(.A1(G375), .A2(new_n1229), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1275), .A2(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(new_n1285), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1285), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(KEYINPUT127), .B2(new_n1247), .ZN(new_n1302));
  XOR2_X1   g1102(.A(new_n1246), .B(KEYINPUT127), .Z(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1303), .B2(new_n1301), .ZN(G402));
endmodule


