//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G146), .ZN(new_n188));
  NOR2_X1   g002(.A1(G125), .A2(G140), .ZN(new_n189));
  AND2_X1   g003(.A1(G125), .A2(G140), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n194), .A2(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n192), .A2(G119), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT76), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G110), .ZN(new_n202));
  INV_X1    g016(.A(G110), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(KEYINPUT24), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT77), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(KEYINPUT24), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(G110), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n197), .A2(new_n200), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n198), .B2(new_n199), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(new_n193), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n213), .A2(new_n203), .A3(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n191), .B1(new_n210), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G125), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT79), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT79), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G125), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT16), .ZN(new_n224));
  INV_X1    g038(.A(G140), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n189), .B1(new_n223), .B2(G140), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(new_n224), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n187), .B1(new_n218), .B2(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n200), .A2(new_n197), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n205), .A2(new_n209), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n213), .A2(new_n216), .ZN(new_n234));
  OAI22_X1  g048(.A1(new_n232), .A2(new_n233), .B1(G110), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n189), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT79), .B(G125), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(new_n225), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT16), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(G146), .A3(new_n226), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n235), .A2(KEYINPUT80), .A3(new_n240), .A4(new_n191), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n232), .A2(new_n233), .B1(G110), .B2(new_n234), .ZN(new_n242));
  AOI21_X1  g056(.A(G146), .B1(new_n239), .B2(new_n226), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n230), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n231), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT22), .B(G137), .ZN(new_n246));
  INV_X1    g060(.A(G953), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(G221), .A3(G234), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n246), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT75), .B(G902), .Z(new_n252));
  NAND4_X1  g066(.A1(new_n231), .A2(new_n241), .A3(new_n244), .A4(new_n249), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n251), .A2(KEYINPUT25), .A3(new_n252), .A4(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G217), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(new_n252), .B2(G234), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT81), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n251), .A2(new_n253), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n263), .B(KEYINPUT82), .Z(new_n264));
  NOR2_X1   g078(.A1(new_n260), .A2(G902), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT81), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n258), .A2(new_n267), .A3(new_n260), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n262), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  XOR2_X1   g083(.A(KEYINPUT26), .B(G101), .Z(new_n270));
  NOR2_X1   g084(.A1(G237), .A2(G953), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G210), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n270), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  INV_X1    g091(.A(G137), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(G134), .ZN(new_n279));
  INV_X1    g093(.A(G134), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G137), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(KEYINPUT11), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n278), .A2(G134), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT11), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(KEYINPUT65), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT65), .B1(new_n283), .B2(new_n284), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n277), .B(new_n282), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n283), .A2(KEYINPUT66), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n278), .A3(G134), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n289), .B(new_n291), .C1(G134), .C2(new_n278), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G131), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT67), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n288), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n229), .A2(KEYINPUT64), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT64), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G146), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n300), .A3(G143), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n229), .A2(G143), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n301), .A2(new_n302), .A3(G128), .A4(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(G143), .B1(new_n298), .B2(new_n300), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n229), .A2(G143), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n301), .A2(KEYINPUT1), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n192), .B1(new_n311), .B2(KEYINPUT68), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n301), .A2(new_n313), .A3(KEYINPUT1), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n310), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n295), .B(new_n297), .C1(new_n306), .C2(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT0), .B(G128), .Z(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n307), .B2(new_n309), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n301), .A2(KEYINPUT0), .A3(G128), .A4(new_n304), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n288), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT65), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n281), .B2(KEYINPUT11), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n285), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n277), .B1(new_n325), .B2(new_n282), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n321), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n316), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT2), .B(G113), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT69), .ZN(new_n331));
  INV_X1    g145(.A(G116), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(G119), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n194), .A2(KEYINPUT69), .A3(G116), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(G119), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n330), .A2(new_n333), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n329), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n339), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n311), .A2(KEYINPUT68), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(G128), .A3(new_n314), .ZN(new_n343));
  INV_X1    g157(.A(new_n310), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n306), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n327), .B(new_n341), .C1(new_n345), .C2(new_n294), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n276), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n327), .B1(new_n345), .B2(new_n294), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n339), .B1(new_n348), .B2(KEYINPUT71), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n327), .B(new_n350), .C1(new_n345), .C2(new_n294), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT28), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n275), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(KEYINPUT72), .B(new_n275), .C1(new_n347), .C2(new_n352), .ZN(new_n356));
  INV_X1    g170(.A(new_n346), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n348), .A2(KEYINPUT30), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n295), .A2(new_n297), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n359), .B(new_n327), .C1(new_n360), .C2(new_n345), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n357), .B1(new_n362), .B2(new_n339), .ZN(new_n363));
  INV_X1    g177(.A(new_n275), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT31), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n341), .B1(new_n358), .B2(new_n361), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT31), .ZN(new_n367));
  NOR4_X1   g181(.A1(new_n366), .A2(new_n367), .A3(new_n275), .A4(new_n357), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n355), .B(new_n356), .C1(new_n365), .C2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(G472), .A2(G902), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT32), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n348), .A2(new_n339), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT74), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT74), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n348), .A2(new_n376), .A3(new_n339), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT73), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n346), .B(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT28), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n348), .A2(KEYINPUT71), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n341), .A3(new_n351), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n276), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n275), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n341), .B1(new_n316), .B2(new_n327), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT28), .B1(new_n388), .B2(new_n357), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n384), .A2(new_n364), .A3(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n275), .B1(new_n366), .B2(new_n357), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n385), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n387), .A2(new_n392), .A3(new_n252), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n369), .A2(new_n373), .B1(new_n393), .B2(G472), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n356), .B1(new_n365), .B2(new_n368), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n353), .A2(new_n354), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n370), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n372), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n269), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT9), .B(G234), .ZN(new_n400));
  OAI21_X1  g214(.A(G221), .B1(new_n400), .B2(G902), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(KEYINPUT83), .ZN(new_n402));
  INV_X1    g216(.A(G469), .ZN(new_n403));
  INV_X1    g217(.A(G902), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n406));
  INV_X1    g220(.A(G104), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n407), .B2(G107), .ZN(new_n408));
  INV_X1    g222(.A(G107), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(KEYINPUT3), .A3(G104), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G101), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n409), .B2(G104), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n407), .A2(KEYINPUT84), .A3(G107), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n411), .A2(new_n412), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n407), .A2(G107), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n409), .A2(G104), .ZN(new_n418));
  OAI21_X1  g232(.A(G101), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(KEYINPUT10), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n315), .B2(new_n306), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n416), .A2(new_n419), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT85), .ZN(new_n424));
  INV_X1    g238(.A(G143), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n424), .B(KEYINPUT1), .C1(new_n425), .C2(G146), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G128), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n308), .B2(KEYINPUT1), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n303), .B1(new_n188), .B2(G143), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n305), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT10), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n322), .A2(new_n326), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n409), .A2(KEYINPUT3), .A3(G104), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT3), .B1(new_n409), .B2(G104), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n414), .B(new_n415), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G101), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(KEYINPUT4), .A3(new_n416), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT4), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n441), .A3(G101), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n321), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n422), .A2(new_n434), .A3(new_n435), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n416), .A2(new_n419), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n305), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n432), .B1(new_n315), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n435), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n447), .A2(KEYINPUT12), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT12), .B1(new_n447), .B2(new_n448), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n444), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G140), .ZN(new_n452));
  INV_X1    g266(.A(G227), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(G953), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n452), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n444), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n301), .A2(new_n304), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n428), .B2(new_n427), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n445), .B1(new_n305), .B2(new_n459), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n439), .A2(KEYINPUT4), .A3(new_n416), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n442), .A2(new_n319), .A3(new_n318), .ZN(new_n462));
  OAI22_X1  g276(.A1(new_n460), .A2(KEYINPUT10), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n302), .B1(new_n188), .B2(G143), .ZN(new_n464));
  OAI21_X1  g278(.A(G128), .B1(new_n464), .B2(new_n313), .ZN(new_n465));
  INV_X1    g279(.A(new_n314), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n344), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n420), .B1(new_n467), .B2(new_n305), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n448), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n451), .A2(new_n455), .B1(new_n457), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n405), .B1(new_n470), .B2(G469), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n444), .B(new_n456), .C1(new_n449), .C2(new_n450), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n456), .B1(new_n469), .B2(new_n444), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n403), .B(new_n252), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n402), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G214), .B1(G237), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n440), .A2(new_n339), .A3(new_n442), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT86), .B(KEYINPUT5), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(G116), .A3(new_n194), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(G113), .C1(new_n337), .C2(new_n480), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n482), .A2(new_n336), .A3(new_n416), .A4(new_n419), .ZN(new_n483));
  XNOR2_X1  g297(.A(G110), .B(G122), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n479), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n339), .A2(new_n442), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n483), .B1(new_n461), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n484), .B(KEYINPUT87), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n485), .A2(KEYINPUT6), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n414), .A2(new_n415), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n412), .B1(new_n490), .B2(new_n411), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n491), .A2(new_n441), .B1(new_n336), .B2(new_n338), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n336), .A2(new_n416), .A3(new_n419), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n492), .A2(new_n440), .B1(new_n493), .B2(new_n482), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n495));
  INV_X1    g309(.A(new_n488), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n320), .B2(new_n223), .ZN(new_n499));
  AOI211_X1 g313(.A(KEYINPUT88), .B(new_n237), .C1(new_n318), .C2(new_n319), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n467), .A2(new_n305), .A3(new_n237), .ZN(new_n502));
  INV_X1    g316(.A(G224), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(G953), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n501), .B2(new_n502), .ZN(new_n507));
  OAI22_X1  g321(.A1(new_n489), .A2(new_n497), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(KEYINPUT7), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n315), .A2(new_n306), .A3(new_n223), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n321), .A2(new_n237), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT7), .A4(new_n505), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n484), .B(KEYINPUT8), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n336), .A2(new_n416), .A3(new_n419), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n481), .A2(G113), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT5), .A4(new_n335), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n517), .B2(KEYINPUT89), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n517), .A2(KEYINPUT89), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n423), .B1(new_n336), .B2(new_n482), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n514), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n512), .A2(new_n513), .A3(new_n485), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n508), .A2(new_n404), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(G210), .B1(G237), .B2(G902), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT90), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n526), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n508), .A2(new_n404), .A3(new_n528), .A4(new_n523), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n478), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n476), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n228), .A2(new_n229), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT91), .ZN(new_n533));
  OR2_X1    g347(.A1(G237), .A2(G953), .ZN(new_n534));
  NAND2_X1  g348(.A1(G143), .A2(G214), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n277), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(G143), .B1(new_n271), .B2(G214), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G214), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n425), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n271), .A2(G143), .A3(G214), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n540), .A2(KEYINPUT91), .A3(new_n277), .A4(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n534), .A2(new_n535), .ZN(new_n544));
  OAI21_X1  g358(.A(G131), .B1(new_n544), .B2(new_n537), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n538), .A2(new_n542), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n545), .A2(new_n543), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n532), .A2(new_n546), .A3(new_n240), .A4(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G113), .B(G122), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(new_n407), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n544), .A2(new_n537), .ZN(new_n551));
  AND2_X1   g365(.A1(KEYINPUT18), .A2(G131), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n191), .B1(new_n238), .B2(new_n229), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n548), .A2(new_n550), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n550), .B1(new_n548), .B2(new_n555), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n404), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n558), .A2(G475), .ZN(new_n559));
  NOR2_X1   g373(.A1(G475), .A2(G902), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n560), .B(KEYINPUT94), .Z(new_n561));
  INV_X1    g375(.A(KEYINPUT19), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n562), .B1(new_n190), .B2(new_n189), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(new_n227), .B2(KEYINPUT19), .ZN(new_n566));
  OAI211_X1 g380(.A(KEYINPUT19), .B(new_n236), .C1(new_n237), .C2(new_n225), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(new_n564), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n188), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n538), .A2(new_n542), .A3(new_n545), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT92), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n538), .A2(new_n542), .A3(new_n572), .A4(new_n545), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n569), .A2(new_n571), .A3(new_n240), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n550), .B1(new_n574), .B2(new_n555), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n561), .B1(new_n575), .B2(new_n556), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT20), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT20), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n578), .B(new_n561), .C1(new_n575), .C2(new_n556), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n559), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G952), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(G953), .ZN(new_n582));
  NAND2_X1  g396(.A1(G234), .A2(G237), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n252), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(G953), .A3(new_n583), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT21), .B(G898), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G478), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(KEYINPUT15), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n425), .A2(G128), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n192), .A2(G143), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(new_n280), .ZN(new_n598));
  XNOR2_X1  g412(.A(G116), .B(G122), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n409), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n332), .A2(KEYINPUT14), .A3(G122), .ZN(new_n601));
  XOR2_X1   g415(.A(G116), .B(G122), .Z(new_n602));
  OAI211_X1 g416(.A(G107), .B(new_n601), .C1(new_n602), .C2(KEYINPUT14), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n598), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(G107), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n600), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n597), .A2(new_n280), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n425), .A2(KEYINPUT13), .A3(G128), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(KEYINPUT95), .A3(new_n596), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT13), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n595), .ZN(new_n611));
  OAI21_X1  g425(.A(G134), .B1(new_n608), .B2(KEYINPUT95), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n606), .B(new_n607), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n604), .A2(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n400), .A2(new_n259), .A3(G953), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n604), .A2(new_n613), .A3(new_n615), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n594), .B1(new_n619), .B2(new_n252), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n586), .B(new_n593), .C1(new_n617), .C2(new_n618), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n580), .A2(new_n591), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n531), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n399), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  NAND2_X1  g440(.A1(new_n369), .A2(new_n252), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n627), .A2(G472), .B1(new_n370), .B2(new_n369), .ZN(new_n628));
  INV_X1    g442(.A(new_n402), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n469), .A2(new_n444), .A3(new_n456), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n447), .A2(KEYINPUT12), .A3(new_n448), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT12), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n306), .B1(new_n416), .B2(new_n419), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n467), .A2(new_n633), .B1(new_n423), .B2(new_n431), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n632), .B1(new_n634), .B2(new_n435), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n463), .A2(new_n468), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n631), .A2(new_n635), .B1(new_n636), .B2(new_n435), .ZN(new_n637));
  OAI211_X1 g451(.A(G469), .B(new_n630), .C1(new_n637), .C2(new_n456), .ZN(new_n638));
  INV_X1    g452(.A(new_n405), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n462), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n641), .A2(new_n440), .B1(new_n432), .B2(new_n433), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n435), .B1(new_n642), .B2(new_n422), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n463), .A2(new_n468), .A3(new_n448), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n455), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI211_X1 g459(.A(G469), .B(new_n586), .C1(new_n645), .C2(new_n472), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n629), .B1(new_n640), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n269), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n628), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n530), .A2(new_n591), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n619), .B(KEYINPUT33), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n586), .A2(new_n592), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n619), .A2(new_n252), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n651), .A2(new_n652), .B1(new_n653), .B2(new_n592), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n650), .A2(new_n580), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT96), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT34), .B(G104), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  INV_X1    g473(.A(new_n577), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT97), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n559), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n577), .A2(KEYINPUT97), .A3(new_n579), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n650), .A2(new_n622), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n649), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  AOI21_X1  g482(.A(new_n267), .B1(new_n258), .B2(new_n260), .ZN(new_n669));
  INV_X1    g483(.A(new_n260), .ZN(new_n670));
  AOI211_X1 g484(.A(KEYINPUT81), .B(new_n670), .C1(new_n256), .C2(new_n257), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT36), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n249), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT98), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n245), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n245), .A2(new_n674), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(KEYINPUT99), .A3(new_n265), .ZN(new_n679));
  INV_X1    g493(.A(new_n677), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n265), .A3(new_n675), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n669), .A2(new_n671), .A3(new_n684), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n685), .A2(new_n531), .A3(new_n623), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n628), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  NAND2_X1  g503(.A1(new_n394), .A2(new_n398), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n496), .B1(new_n479), .B2(new_n483), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT6), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n495), .B1(new_n494), .B2(new_n484), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n693), .B1(new_n694), .B2(new_n692), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n501), .A2(new_n502), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n504), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(G902), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n528), .B1(new_n700), .B2(new_n523), .ZN(new_n701));
  INV_X1    g515(.A(new_n529), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n477), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n647), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n679), .A2(new_n683), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n262), .A2(new_n268), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n622), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n584), .B(KEYINPUT101), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT100), .ZN(new_n710));
  INV_X1    g524(.A(G900), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n588), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT100), .B1(new_n587), .B2(G900), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AND4_X1   g529(.A1(new_n707), .A2(new_n662), .A3(new_n663), .A4(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n704), .A2(new_n706), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n691), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n192), .ZN(G30));
  NAND2_X1  g533(.A1(new_n527), .A2(new_n529), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT38), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n577), .A2(new_n579), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n558), .A2(G475), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n622), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NOR4_X1   g540(.A1(new_n722), .A2(new_n706), .A3(new_n478), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n346), .B(KEYINPUT73), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n275), .A3(new_n375), .A4(new_n377), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n729), .B(new_n404), .C1(new_n275), .C2(new_n363), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G472), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(KEYINPUT102), .A3(G472), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n733), .A2(new_n734), .B1(new_n369), .B2(new_n373), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n398), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n714), .B(KEYINPUT39), .Z(new_n737));
  NAND2_X1  g551(.A1(new_n476), .A2(new_n737), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT40), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(KEYINPUT40), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n727), .A2(new_n736), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G143), .ZN(G45));
  NAND2_X1  g556(.A1(new_n723), .A2(new_n724), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n653), .A2(new_n592), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n619), .B(KEYINPUT33), .Z(new_n745));
  INV_X1    g559(.A(new_n652), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n743), .A2(new_n747), .A3(new_n715), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT103), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n743), .A2(new_n747), .A3(KEYINPUT103), .A4(new_n715), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n704), .A2(new_n706), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n691), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n229), .ZN(G48));
  NAND2_X1  g568(.A1(new_n635), .A2(new_n631), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n469), .A2(new_n444), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n755), .A2(new_n457), .B1(new_n756), .B2(new_n455), .ZN(new_n757));
  OAI21_X1  g571(.A(G469), .B1(new_n757), .B2(new_n586), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n629), .A3(new_n475), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT104), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(KEYINPUT104), .A3(new_n629), .A4(new_n475), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n399), .A2(new_n655), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT41), .B(G113), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G15));
  NAND3_X1  g581(.A1(new_n399), .A2(new_n665), .A3(new_n764), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G116), .ZN(G18));
  NAND3_X1  g583(.A1(new_n761), .A2(new_n530), .A3(new_n762), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n761), .A2(new_n530), .A3(KEYINPUT105), .A4(new_n762), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n623), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n706), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n398), .B2(new_n394), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G119), .ZN(G21));
  NOR3_X1   g593(.A1(new_n763), .A2(new_n650), .A3(new_n726), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT106), .B(G472), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n369), .B2(new_n252), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n365), .A2(new_n368), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n381), .A2(new_n384), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n275), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n371), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n783), .A2(new_n787), .A3(new_n269), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n780), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G122), .ZN(G24));
  NAND2_X1  g604(.A1(new_n750), .A2(new_n751), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n783), .A2(new_n791), .A3(new_n787), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n774), .A2(new_n706), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G125), .ZN(G27));
  NOR2_X1   g608(.A1(new_n720), .A2(new_n478), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n476), .A2(new_n750), .A3(new_n751), .A4(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(new_n269), .ZN(new_n797));
  AND4_X1   g611(.A1(KEYINPUT42), .A2(new_n690), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT42), .B1(new_n399), .B2(new_n796), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n277), .ZN(G33));
  INV_X1    g615(.A(new_n795), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n647), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(new_n716), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n399), .ZN(new_n805));
  XOR2_X1   g619(.A(KEYINPUT107), .B(G134), .Z(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(G36));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n743), .A2(KEYINPUT43), .A3(new_n654), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n580), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n743), .A2(KEYINPUT109), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n812), .A3(new_n747), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n809), .B1(new_n813), .B2(KEYINPUT43), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n706), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT44), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n815), .A2(new_n628), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n808), .B1(new_n817), .B2(new_n802), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n813), .A2(KEYINPUT43), .ZN(new_n819));
  INV_X1    g633(.A(new_n809), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n819), .A2(new_n706), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n627), .A2(G472), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n397), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(KEYINPUT110), .B(new_n795), .C1(new_n824), .C2(new_n816), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT44), .B1(new_n821), .B2(new_n823), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT46), .ZN(new_n827));
  OAI21_X1  g641(.A(G469), .B1(new_n470), .B2(KEYINPUT45), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n630), .B1(new_n637), .B2(new_n456), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT45), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT108), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT108), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n470), .A2(new_n832), .A3(KEYINPUT45), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n828), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n827), .B1(new_n834), .B2(new_n405), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n475), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n834), .A2(new_n827), .A3(new_n405), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n629), .B(new_n737), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n826), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n818), .A2(new_n825), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(G137), .ZN(G39));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n791), .A2(new_n802), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n691), .A2(new_n842), .A3(new_n269), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n269), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT111), .B1(new_n845), .B2(new_n690), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n834), .A2(new_n405), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT46), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n475), .A3(new_n835), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n849), .A2(KEYINPUT47), .A3(new_n629), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT47), .B1(new_n849), .B2(new_n629), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n844), .B(new_n846), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(G140), .ZN(G42));
  AND2_X1   g667(.A1(new_n814), .A2(new_n709), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n399), .A2(new_n854), .A3(new_n764), .A4(new_n795), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT48), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n788), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n774), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n764), .A2(new_n797), .A3(new_n585), .A4(new_n795), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n736), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n743), .A3(new_n747), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n857), .A2(new_n582), .A3(new_n860), .A4(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n850), .A2(new_n851), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n758), .A2(new_n475), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n629), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n802), .B(new_n858), .C1(new_n865), .C2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT50), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n764), .A2(new_n478), .A3(new_n722), .ZN(new_n871));
  OR3_X1    g685(.A1(new_n858), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n858), .B2(new_n871), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n854), .A2(new_n764), .A3(new_n795), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n783), .A2(new_n685), .A3(new_n787), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n743), .A2(new_n747), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n875), .A2(new_n876), .B1(new_n862), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT51), .B1(new_n869), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n865), .A2(new_n868), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n795), .A3(new_n859), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n882), .A2(new_n883), .A3(new_n874), .A4(new_n878), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n864), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT115), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n774), .A2(new_n706), .A3(new_n792), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n685), .A2(new_n531), .ZN(new_n888));
  INV_X1    g702(.A(new_n791), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n690), .B(new_n888), .C1(new_n716), .C2(new_n889), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n402), .B(new_n714), .C1(new_n471), .C2(new_n475), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n720), .A2(new_n477), .A3(new_n725), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n685), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n736), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT113), .B1(new_n887), .B2(new_n896), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n752), .A2(new_n717), .B1(new_n398), .B2(new_n394), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n893), .B1(new_n398), .B2(new_n735), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT113), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n901), .A3(new_n793), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT52), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT52), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n900), .B2(new_n793), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n774), .A2(new_n777), .B1(new_n788), .B2(new_n780), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n743), .A2(new_n654), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n743), .B2(new_n707), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n650), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n628), .A2(new_n648), .A3(new_n910), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n399), .A2(new_n624), .B1(new_n686), .B2(new_n628), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n399), .B(new_n764), .C1(new_n655), .C2(new_n665), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n907), .A2(new_n911), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n805), .B1(new_n798), .B2(new_n799), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n803), .A2(new_n706), .ZN(new_n916));
  INV_X1    g730(.A(new_n792), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n664), .A2(new_n707), .A3(new_n714), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n690), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n914), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT53), .B1(new_n906), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n900), .A2(new_n901), .A3(new_n793), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n901), .B1(new_n900), .B2(new_n793), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n904), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n897), .A2(KEYINPUT52), .A3(new_n902), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n921), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT53), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT54), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT114), .ZN(new_n931));
  INV_X1    g745(.A(new_n905), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n925), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n778), .A2(new_n789), .A3(new_n911), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n913), .A2(new_n912), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n915), .ZN(new_n937));
  INV_X1    g751(.A(new_n920), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT53), .A4(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n931), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n927), .A2(new_n928), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT54), .ZN(new_n942));
  NOR4_X1   g756(.A1(new_n914), .A2(new_n915), .A3(new_n928), .A4(new_n920), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n943), .A2(KEYINPUT114), .A3(new_n925), .A4(new_n932), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n940), .A2(new_n941), .A3(new_n942), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n930), .A2(new_n945), .ZN(new_n946));
  OAI22_X1  g760(.A1(new_n886), .A2(new_n946), .B1(G952), .B2(G953), .ZN(new_n947));
  INV_X1    g761(.A(new_n736), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n866), .B(KEYINPUT49), .Z(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(new_n722), .A3(new_n949), .ZN(new_n950));
  NOR4_X1   g764(.A1(new_n269), .A2(new_n813), .A3(new_n478), .A4(new_n402), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT112), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n947), .B1(new_n950), .B2(new_n952), .ZN(G75));
  NAND3_X1  g767(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n586), .A3(new_n526), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT56), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n695), .B(new_n699), .ZN(new_n957));
  XNOR2_X1  g771(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n955), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n955), .B2(new_n956), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n247), .A2(G952), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G51));
  XNOR2_X1  g777(.A(new_n405), .B(KEYINPUT57), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n939), .A2(new_n903), .A3(new_n905), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n965), .A2(KEYINPUT114), .B1(new_n928), .B2(new_n927), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n942), .B1(new_n966), .B2(new_n940), .ZN(new_n967));
  INV_X1    g781(.A(new_n945), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n757), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n954), .A2(new_n586), .A3(new_n834), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n962), .B1(new_n971), .B2(new_n972), .ZN(G54));
  NAND4_X1  g787(.A1(new_n954), .A2(KEYINPUT58), .A3(G475), .A4(new_n586), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n575), .A2(new_n556), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n974), .A2(new_n976), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n977), .A2(new_n978), .A3(new_n962), .ZN(G60));
  INV_X1    g793(.A(new_n962), .ZN(new_n980));
  NAND2_X1  g794(.A1(G478), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT59), .Z(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n930), .B2(new_n945), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n980), .B1(new_n983), .B2(new_n651), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n745), .A2(new_n982), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n967), .B2(new_n968), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(KEYINPUT117), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT117), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n988), .B(new_n985), .C1(new_n967), .C2(new_n968), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n984), .B1(new_n987), .B2(new_n989), .ZN(G63));
  NAND2_X1  g804(.A1(G217), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT118), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT60), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n954), .A2(new_n678), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n980), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n264), .B1(new_n954), .B2(new_n993), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n994), .A2(KEYINPUT119), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT61), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n999), .B(new_n998), .C1(new_n995), .C2(new_n996), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(G66));
  OAI21_X1  g817(.A(G953), .B1(new_n589), .B2(new_n503), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n936), .B2(G953), .ZN(new_n1005));
  INV_X1    g819(.A(G898), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n695), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT120), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1005), .B(new_n1008), .ZN(G69));
  OAI21_X1  g823(.A(G953), .B1(new_n453), .B2(new_n711), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n399), .A2(new_n892), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n838), .A2(new_n1011), .ZN(new_n1012));
  NOR4_X1   g826(.A1(new_n1012), .A2(new_n887), .A3(new_n718), .A4(new_n753), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1013), .A2(new_n840), .A3(new_n852), .A4(new_n937), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1014), .A2(G953), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n566), .A2(new_n568), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n362), .B(new_n1016), .Z(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n711), .B2(new_n247), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT124), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1010), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n793), .A2(new_n741), .A3(new_n890), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT62), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n738), .A2(new_n802), .A3(new_n909), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n399), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n840), .A2(new_n852), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(KEYINPUT122), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT62), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1022), .B(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT122), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n852), .A2(new_n1025), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n840), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n247), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1017), .B(KEYINPUT121), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1019), .B1(new_n1036), .B2(KEYINPUT123), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT123), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1034), .A2(new_n1038), .A3(new_n1035), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1021), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1019), .ZN(new_n1041));
  AOI21_X1  g855(.A(G953), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1035), .ZN(new_n1043));
  OAI21_X1  g857(.A(KEYINPUT123), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AND4_X1   g858(.A1(new_n1041), .A2(new_n1039), .A3(new_n1021), .A4(new_n1044), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1040), .A2(new_n1045), .ZN(G72));
  NAND2_X1  g860(.A1(G472), .A2(G902), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(KEYINPUT63), .Z(new_n1048));
  XNOR2_X1  g862(.A(new_n1048), .B(KEYINPUT125), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1049), .B1(new_n1014), .B2(new_n914), .ZN(new_n1050));
  NOR3_X1   g864(.A1(new_n366), .A2(new_n364), .A3(new_n357), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n962), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g866(.A(new_n1052), .B(KEYINPUT126), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1049), .B1(new_n1033), .B2(new_n914), .ZN(new_n1054));
  OAI211_X1 g868(.A(new_n1054), .B(new_n364), .C1(new_n357), .C2(new_n366), .ZN(new_n1055));
  INV_X1    g869(.A(KEYINPUT127), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1056), .B1(new_n363), .B2(new_n364), .ZN(new_n1057));
  XOR2_X1   g871(.A(new_n1057), .B(new_n391), .Z(new_n1058));
  OAI211_X1 g872(.A(new_n1048), .B(new_n1058), .C1(new_n922), .C2(new_n929), .ZN(new_n1059));
  AND3_X1   g873(.A1(new_n1053), .A2(new_n1055), .A3(new_n1059), .ZN(G57));
endmodule


