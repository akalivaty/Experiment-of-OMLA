//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  OR2_X1    g001(.A1(G43gat), .A2(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G43gat), .A2(G50gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n206), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT14), .B(G29gat), .Z(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(G36gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT93), .B(G43gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n202), .B(new_n204), .C1(new_n210), .C2(G50gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n205), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(new_n205), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n215), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT17), .B1(new_n217), .B2(new_n212), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  INV_X1    g018(.A(G1gat), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(KEYINPUT16), .A3(new_n220), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT94), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(G8gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(new_n223), .A3(G8gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(G8gat), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n221), .A2(new_n222), .A3(new_n227), .A4(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n216), .A2(new_n218), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n217), .A2(new_n212), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(new_n228), .A3(new_n226), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT18), .A4(new_n233), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n229), .B1(new_n212), .B2(new_n217), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n232), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(new_n233), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n237), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G197gat), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT11), .B(G169gat), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(KEYINPUT12), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n248), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n250), .A2(new_n236), .A3(new_n237), .A4(new_n242), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT35), .ZN(new_n254));
  XNOR2_X1  g053(.A(G78gat), .B(G106gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n255), .B(G50gat), .Z(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(G228gat), .A2(G233gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(G155gat), .B(G162gat), .ZN(new_n259));
  INV_X1    g058(.A(G148gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G141gat), .ZN(new_n261));
  INV_X1    g060(.A(G141gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G148gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n259), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT2), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT79), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(KEYINPUT79), .A3(KEYINPUT2), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n259), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n262), .A2(KEYINPUT78), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT78), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G141gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n276), .A3(G148gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n261), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n266), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(G211gat), .A2(G218gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(G211gat), .A2(G218gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g081(.A1(G197gat), .A2(G204gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(G197gat), .A2(G204gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G211gat), .B(G218gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(G197gat), .B(G204gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n286), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(new_n291), .A3(KEYINPUT88), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT88), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n288), .A2(new_n289), .A3(new_n294), .A4(new_n290), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n279), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n287), .A2(new_n291), .ZN(new_n299));
  XOR2_X1   g098(.A(G155gat), .B(G162gat), .Z(new_n300));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT77), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT77), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT2), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G141gat), .B(G148gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n300), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n261), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT78), .B(G141gat), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(G148gat), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n307), .B(new_n297), .C1(new_n272), .C2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n299), .B1(new_n311), .B2(new_n293), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n258), .B1(new_n298), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT89), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT89), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n315), .B(new_n258), .C1(new_n298), .C2(new_n312), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT3), .B1(new_n299), .B2(new_n293), .ZN(new_n318));
  OAI211_X1 g117(.A(G228gat), .B(G233gat), .C1(new_n318), .C2(new_n279), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(new_n312), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n257), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  AOI211_X1 g121(.A(G22gat), .B(new_n320), .C1(new_n314), .C2(new_n316), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n256), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n311), .A2(new_n293), .ZN(new_n325));
  INV_X1    g124(.A(new_n297), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n295), .A2(new_n293), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(new_n292), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n325), .A2(new_n299), .B1(new_n328), .B2(new_n279), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n315), .B1(new_n329), .B2(new_n258), .ZN(new_n330));
  INV_X1    g129(.A(new_n316), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n321), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G22gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n256), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n257), .A3(new_n321), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n324), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n336), .A3(new_n338), .ZN(new_n341));
  INV_X1    g140(.A(G183gat), .ZN(new_n342));
  INV_X1    g141(.A(G190gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n343), .A3(KEYINPUT65), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT65), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(G183gat), .B2(G190gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT24), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT24), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(G183gat), .A3(G190gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT66), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT66), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n347), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(G169gat), .B2(G176gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n357), .A2(G169gat), .A3(G176gat), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT67), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT23), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT67), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n358), .A4(new_n359), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n354), .A2(new_n356), .A3(new_n362), .A4(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT25), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n349), .A2(new_n351), .B1(new_n342), .B2(new_n343), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n364), .A2(new_n359), .A3(new_n358), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n370), .A2(new_n371), .A3(new_n368), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G113gat), .B(G120gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G127gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G134gat), .ZN(new_n379));
  INV_X1    g178(.A(G134gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(G127gat), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n375), .A2(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G120gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G113gat), .ZN(new_n384));
  INV_X1    g183(.A(G113gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G120gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G127gat), .B(G134gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n376), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT27), .B(G183gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n343), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT28), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(G169gat), .B2(G176gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n363), .A2(KEYINPUT26), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n396), .A2(new_n348), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n374), .A2(new_n390), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G227gat), .ZN(new_n401));
  INV_X1    g200(.A(G233gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n382), .A2(new_n389), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n372), .B1(new_n367), .B2(new_n368), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n394), .A2(new_n398), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n400), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT34), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT70), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT69), .B(G71gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G99gat), .ZN(new_n414));
  XOR2_X1   g213(.A(G15gat), .B(G43gat), .Z(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  XOR2_X1   g215(.A(new_n403), .B(KEYINPUT64), .Z(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n400), .B2(new_n408), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n416), .B1(new_n419), .B2(KEYINPUT33), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT32), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n417), .A2(KEYINPUT34), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n400), .A2(new_n408), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n420), .A2(new_n422), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n412), .A2(new_n423), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n410), .A2(new_n411), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT70), .B1(new_n409), .B2(KEYINPUT34), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n426), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n420), .A2(new_n422), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n340), .A2(new_n341), .A3(new_n427), .A4(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G226gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(new_n402), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(KEYINPUT29), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n374), .B2(new_n399), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT72), .B1(new_n406), .B2(new_n407), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT72), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n347), .A2(new_n352), .A3(new_n355), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n355), .B1(new_n347), .B2(new_n352), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n362), .A2(new_n366), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT25), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n399), .B(new_n441), .C1(new_n446), .C2(new_n372), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n439), .B1(new_n448), .B2(new_n436), .ZN(new_n449));
  INV_X1    g248(.A(new_n299), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT73), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n440), .A2(new_n447), .A3(new_n437), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n374), .A2(new_n399), .A3(new_n436), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT73), .ZN(new_n455));
  INV_X1    g254(.A(new_n436), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n456), .B1(new_n440), .B2(new_n447), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n455), .B(new_n299), .C1(new_n457), .C2(new_n439), .ZN(new_n458));
  XOR2_X1   g257(.A(G8gat), .B(G36gat), .Z(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT75), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n460), .B(KEYINPUT76), .Z(new_n461));
  XNOR2_X1  g260(.A(G64gat), .B(G92gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n451), .A2(new_n454), .A3(new_n458), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT30), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n458), .A2(new_n454), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT30), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n451), .A4(new_n463), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT74), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n448), .A2(new_n436), .ZN(new_n471));
  INV_X1    g270(.A(new_n439), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n455), .B1(new_n473), .B2(new_n299), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n454), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n451), .A2(KEYINPUT74), .A3(new_n454), .A4(new_n458), .ZN(new_n477));
  INV_X1    g276(.A(new_n463), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n469), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n434), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G1gat), .B(G29gat), .Z(new_n482));
  XNOR2_X1  g281(.A(G57gat), .B(G85gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT6), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n307), .B1(new_n272), .B2(new_n310), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT82), .B1(new_n491), .B2(new_n405), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n278), .A2(new_n259), .A3(new_n271), .A4(new_n270), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT82), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n390), .A2(new_n493), .A3(new_n494), .A4(new_n307), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n491), .A2(KEYINPUT3), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n382), .A2(new_n389), .A3(KEYINPUT80), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT80), .B1(new_n382), .B2(new_n389), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n498), .B(new_n311), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n279), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n497), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n491), .B1(new_n499), .B2(new_n500), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n507), .A2(new_n492), .A3(new_n495), .ZN(new_n508));
  INV_X1    g307(.A(new_n502), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT83), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n508), .A2(KEYINPUT83), .A3(new_n509), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(KEYINPUT5), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT5), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n510), .B2(new_n511), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(KEYINPUT84), .A3(new_n513), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n506), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT4), .B1(new_n279), .B2(new_n390), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n501), .A2(new_n517), .A3(new_n502), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT86), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n488), .B(new_n490), .C1(new_n520), .C2(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n518), .A2(KEYINPUT84), .A3(new_n513), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT84), .B1(new_n518), .B2(new_n513), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n505), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT86), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n526), .B(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n531), .A2(new_n533), .A3(new_n489), .A4(new_n486), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT92), .B1(new_n481), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n476), .A2(KEYINPUT37), .A3(new_n477), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT37), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n451), .A2(new_n538), .A3(new_n454), .A4(new_n458), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n539), .A2(new_n478), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT38), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n452), .A2(new_n299), .A3(new_n453), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n543), .A2(KEYINPUT37), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n450), .B1(new_n457), .B2(new_n439), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT38), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(new_n539), .A3(new_n478), .ZN(new_n547));
  AND4_X1   g346(.A1(new_n534), .A2(new_n547), .A3(new_n528), .A4(new_n464), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n340), .A2(new_n341), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT90), .B(KEYINPUT40), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n522), .B1(new_n496), .B2(KEYINPUT4), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n502), .B1(new_n552), .B2(new_n501), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT39), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n486), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n521), .A2(new_n523), .A3(new_n501), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n509), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n507), .A2(new_n492), .A3(new_n495), .A4(new_n502), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT39), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  AOI211_X1 g360(.A(KEYINPUT91), .B(new_n551), .C1(new_n555), .C2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT91), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n556), .A2(new_n554), .A3(new_n509), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(new_n487), .C1(new_n553), .C2(new_n559), .ZN(new_n565));
  INV_X1    g364(.A(new_n551), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n487), .B1(new_n531), .B2(new_n533), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n555), .A2(KEYINPUT40), .A3(new_n561), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n550), .B1(new_n571), .B2(new_n480), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n549), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n535), .A2(new_n479), .A3(new_n469), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n427), .A2(new_n433), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT36), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n576), .A2(KEYINPUT71), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n576), .A2(KEYINPUT71), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n427), .B(new_n433), .C1(new_n580), .C2(new_n577), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n574), .A2(new_n550), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n254), .A2(new_n536), .B1(new_n573), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT92), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n469), .A2(new_n479), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n340), .A2(new_n341), .ZN(new_n586));
  INV_X1    g385(.A(new_n575), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n528), .A2(new_n534), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR3_X1   g389(.A1(new_n434), .A2(new_n480), .A3(new_n589), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT92), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n590), .A2(KEYINPUT35), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n253), .B1(new_n583), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n594), .A2(new_n589), .ZN(new_n595));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596));
  OR2_X1    g395(.A1(G57gat), .A2(G64gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(G57gat), .A2(G64gat), .ZN(new_n598));
  AND2_X1   g397(.A1(G71gat), .A2(G78gat), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(KEYINPUT9), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT96), .ZN(new_n601));
  NOR2_X1   g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n600), .B(KEYINPUT96), .C1(new_n599), .C2(new_n602), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G231gat), .A2(G233gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT98), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(G231gat), .A3(G233gat), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n609), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n611), .B1(new_n609), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n596), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n609), .A2(new_n613), .ZN(new_n617));
  INV_X1    g416(.A(new_n611), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n596), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n609), .A2(new_n611), .A3(new_n613), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n604), .A2(new_n605), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT21), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n229), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(new_n229), .B2(new_n624), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n616), .A2(new_n622), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n616), .B2(new_n622), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G134gat), .B(G162gat), .Z(new_n633));
  AND2_X1   g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(KEYINPUT41), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT100), .ZN(new_n637));
  NAND2_X1  g436(.A1(G85gat), .A2(G92gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT7), .ZN(new_n639));
  NAND2_X1  g438(.A1(G99gat), .A2(G106gat), .ZN(new_n640));
  INV_X1    g439(.A(G85gat), .ZN(new_n641));
  INV_X1    g440(.A(G92gat), .ZN(new_n642));
  AOI22_X1  g441(.A1(KEYINPUT8), .A2(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G99gat), .B(G106gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n644), .A2(KEYINPUT99), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n639), .A2(new_n645), .A3(new_n643), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(KEYINPUT99), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n216), .A2(new_n218), .A3(new_n647), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n647), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n652), .A2(new_n231), .B1(KEYINPUT41), .B2(new_n634), .ZN(new_n653));
  XOR2_X1   g452(.A(G190gat), .B(G218gat), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n651), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n655), .B1(new_n651), .B2(new_n653), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n637), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n651), .A2(new_n653), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n654), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n636), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n651), .A2(new_n653), .A3(new_n655), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n632), .A2(KEYINPUT101), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT101), .B1(new_n632), .B2(new_n665), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(G230gat), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n402), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT10), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n649), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n648), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n644), .A2(new_n676), .A3(new_n646), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n606), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n623), .B1(new_n650), .B2(new_n647), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n675), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n652), .A2(KEYINPUT10), .A3(new_n623), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n674), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n674), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n680), .A2(new_n681), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n672), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n652), .A2(new_n606), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n678), .A2(new_n679), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n623), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT10), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n683), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n685), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n686), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n671), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n687), .A2(new_n695), .A3(KEYINPUT103), .ZN(new_n696));
  AOI21_X1  g495(.A(KEYINPUT103), .B1(new_n687), .B2(new_n695), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n668), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n595), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G1gat), .ZN(G1324gat));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n594), .A2(new_n700), .A3(new_n480), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT16), .B(G8gat), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n706), .A2(KEYINPUT42), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(G8gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(KEYINPUT42), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(G1325gat));
  NAND2_X1  g509(.A1(new_n594), .A2(new_n700), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n579), .A2(new_n581), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G15gat), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n575), .A2(G15gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n711), .B2(new_n715), .ZN(G1326gat));
  NOR2_X1   g515(.A1(new_n711), .A2(new_n586), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT43), .B(G22gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1327gat));
  INV_X1    g518(.A(new_n698), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n632), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n658), .A2(new_n664), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n595), .A2(new_n206), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT45), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n571), .A2(new_n480), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n586), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n547), .A2(new_n528), .A3(new_n534), .A4(new_n464), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(KEYINPUT38), .B2(new_n541), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n582), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n584), .B(new_n254), .C1(new_n588), .C2(new_n589), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT35), .B1(new_n591), .B2(KEYINPUT92), .ZN(new_n738));
  NOR4_X1   g537(.A1(new_n434), .A2(new_n480), .A3(new_n589), .A4(new_n584), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n736), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n731), .B1(new_n740), .B2(new_n722), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n665), .B1(new_n583), .B2(new_n593), .ZN(new_n743));
  INV_X1    g542(.A(new_n729), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n721), .A2(new_n252), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G29gat), .B1(new_n749), .B2(new_n535), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n726), .A2(new_n750), .ZN(G1328gat));
  NOR2_X1   g550(.A1(new_n723), .A2(G36gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n594), .A2(new_n480), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT106), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(KEYINPUT107), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n755), .A2(KEYINPUT107), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G36gat), .B1(new_n749), .B2(new_n585), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n758), .B(new_n759), .C1(new_n754), .C2(new_n756), .ZN(G1329gat));
  OAI21_X1  g559(.A(new_n210), .B1(new_n749), .B2(new_n713), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n723), .A2(new_n210), .A3(new_n575), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n594), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT47), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n210), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n747), .B1(new_n742), .B2(new_n745), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(new_n712), .ZN(new_n770));
  INV_X1    g569(.A(new_n763), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n765), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n767), .A2(new_n772), .ZN(G1330gat));
  AND3_X1   g572(.A1(new_n740), .A2(new_n722), .A3(new_n744), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n550), .B(new_n748), .C1(new_n774), .C2(new_n741), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G50gat), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT110), .A2(KEYINPUT48), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n586), .A2(G50gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n724), .B1(new_n778), .B2(KEYINPUT109), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(KEYINPUT109), .B2(new_n778), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n777), .B1(new_n594), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(KEYINPUT110), .A2(KEYINPUT48), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1331gat));
  AND4_X1   g583(.A1(new_n668), .A2(new_n740), .A3(new_n720), .A4(new_n253), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n589), .ZN(new_n786));
  XOR2_X1   g585(.A(KEYINPUT111), .B(G57gat), .Z(new_n787));
  XNOR2_X1  g586(.A(new_n786), .B(new_n787), .ZN(G1332gat));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n480), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n790));
  XOR2_X1   g589(.A(KEYINPUT49), .B(G64gat), .Z(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(G1333gat));
  NAND2_X1  g591(.A1(new_n785), .A2(new_n712), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n575), .A2(G71gat), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n793), .A2(G71gat), .B1(new_n785), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g595(.A1(new_n785), .A2(new_n550), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g597(.A1(new_n252), .A2(new_n632), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n698), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n746), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G85gat), .B1(new_n802), .B2(new_n535), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT51), .B1(new_n743), .B2(new_n799), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  AND4_X1   g604(.A1(KEYINPUT51), .A2(new_n740), .A3(new_n722), .A4(new_n799), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n808), .A2(new_n641), .A3(new_n720), .A4(new_n589), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n803), .A2(new_n809), .ZN(G1336gat));
  OAI21_X1  g609(.A(G92gat), .B1(new_n802), .B2(new_n585), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n585), .A2(G92gat), .A3(new_n698), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n805), .B2(new_n807), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n811), .A2(new_n812), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n801), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n742), .B2(new_n745), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n642), .B1(new_n819), .B2(new_n480), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT52), .B1(new_n820), .B2(new_n815), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n821), .ZN(G1337gat));
  OAI21_X1  g621(.A(G99gat), .B1(new_n802), .B2(new_n713), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n575), .A2(G99gat), .A3(new_n698), .ZN(new_n824));
  XOR2_X1   g623(.A(new_n824), .B(KEYINPUT112), .Z(new_n825));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(G1338gat));
  NOR3_X1   g626(.A1(new_n586), .A2(G106gat), .A3(new_n698), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n804), .B2(new_n806), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(KEYINPUT113), .B(new_n828), .C1(new_n804), .C2(new_n806), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n550), .B(new_n801), .C1(new_n774), .C2(new_n741), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(G106gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT53), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n808), .A2(new_n837), .A3(new_n828), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n829), .A2(KEYINPUT114), .ZN(new_n839));
  XNOR2_X1  g638(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n834), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n836), .A2(new_n841), .ZN(G1339gat));
  NAND4_X1  g641(.A1(new_n668), .A2(KEYINPUT116), .A3(new_n698), .A4(new_n253), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT101), .ZN(new_n844));
  INV_X1    g643(.A(new_n631), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n616), .A2(new_n622), .A3(new_n629), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n844), .B1(new_n847), .B2(new_n722), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n632), .A2(KEYINPUT101), .A3(new_n665), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n848), .A2(new_n698), .A3(new_n849), .A4(new_n253), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n682), .A2(new_n674), .A3(new_n683), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n693), .A2(KEYINPUT54), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g654(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n684), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n672), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT55), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n855), .A2(KEYINPUT55), .A3(new_n672), .A4(new_n857), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n860), .A2(new_n695), .A3(new_n252), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n239), .A2(new_n241), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n233), .B1(new_n230), .B2(new_n232), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n247), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n251), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n696), .B2(new_n697), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n722), .B1(new_n862), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n860), .A2(new_n695), .A3(new_n861), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n722), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n847), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n550), .B1(new_n853), .B2(new_n872), .ZN(new_n873));
  AND4_X1   g672(.A1(new_n589), .A2(new_n873), .A3(new_n587), .A4(new_n585), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n385), .B1(new_n874), .B2(new_n252), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT118), .Z(new_n876));
  AOI21_X1  g675(.A(new_n535), .B1(new_n853), .B2(new_n872), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n481), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(new_n385), .A3(new_n252), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n876), .A2(new_n879), .ZN(G1340gat));
  AOI21_X1  g679(.A(G120gat), .B1(new_n878), .B2(new_n720), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n698), .A2(new_n383), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n874), .B2(new_n882), .ZN(G1341gat));
  NAND3_X1  g682(.A1(new_n878), .A2(new_n378), .A3(new_n632), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n874), .A2(new_n632), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n378), .ZN(G1342gat));
  AND2_X1   g685(.A1(new_n874), .A2(new_n722), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(new_n380), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n878), .A2(new_n380), .A3(new_n722), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(KEYINPUT56), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(KEYINPUT56), .B2(new_n889), .ZN(G1343gat));
  NOR3_X1   g690(.A1(new_n712), .A2(new_n586), .A3(new_n480), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(G141gat), .A3(new_n253), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(KEYINPUT58), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n712), .A2(new_n535), .A3(new_n480), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n853), .A2(new_n872), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT57), .B1(new_n897), .B2(new_n550), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n899), .B(new_n586), .C1(new_n853), .C2(new_n872), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n896), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n901), .A2(new_n253), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n895), .B1(new_n903), .B2(new_n309), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT119), .B(new_n896), .C1(new_n898), .C2(new_n900), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n252), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n909));
  INV_X1    g708(.A(new_n309), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n911), .A2(new_n912), .A3(new_n894), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n904), .B1(new_n913), .B2(new_n914), .ZN(G1344gat));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n916));
  INV_X1    g715(.A(new_n893), .ZN(new_n917));
  AOI211_X1 g716(.A(new_n916), .B(G148gat), .C1(new_n917), .C2(new_n720), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n906), .A2(new_n907), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n916), .A3(new_n720), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n872), .A2(new_n850), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT57), .B1(new_n921), .B2(new_n550), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n720), .B(new_n896), .C1(new_n900), .C2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n260), .B1(new_n923), .B2(KEYINPUT59), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n918), .B1(new_n920), .B2(new_n924), .ZN(G1345gat));
  INV_X1    g724(.A(G155gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n917), .A2(new_n926), .A3(new_n632), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n919), .A2(new_n632), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n926), .ZN(G1346gat));
  AOI21_X1  g728(.A(G162gat), .B1(new_n917), .B2(new_n722), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n722), .A2(G162gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n919), .B2(new_n931), .ZN(G1347gat));
  AOI21_X1  g731(.A(new_n589), .B1(new_n853), .B2(new_n872), .ZN(new_n933));
  AND4_X1   g732(.A1(new_n586), .A2(new_n933), .A3(new_n587), .A4(new_n480), .ZN(new_n934));
  AOI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n252), .ZN(new_n935));
  AND4_X1   g734(.A1(new_n535), .A2(new_n873), .A3(new_n587), .A4(new_n480), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n252), .A2(G169gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(G1348gat));
  INV_X1    g737(.A(G176gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n934), .A2(new_n939), .A3(new_n720), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n936), .A2(new_n720), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n939), .ZN(G1349gat));
  NAND3_X1  g741(.A1(new_n934), .A2(new_n632), .A3(new_n391), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n936), .A2(new_n632), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n342), .ZN(new_n945));
  XOR2_X1   g744(.A(KEYINPUT121), .B(KEYINPUT60), .Z(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(G1350gat));
  AOI21_X1  g746(.A(new_n343), .B1(new_n936), .B2(new_n722), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT61), .Z(new_n949));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n343), .A3(new_n722), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT122), .Z(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1351gat));
  AND4_X1   g751(.A1(new_n550), .A2(new_n933), .A3(new_n480), .A4(new_n713), .ZN(new_n953));
  XOR2_X1   g752(.A(KEYINPUT123), .B(G197gat), .Z(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n252), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n900), .A2(new_n922), .ZN(new_n956));
  NOR4_X1   g755(.A1(new_n956), .A2(new_n589), .A3(new_n585), .A4(new_n712), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n252), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(KEYINPUT124), .ZN(new_n959));
  INV_X1    g758(.A(new_n954), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(new_n958), .B2(KEYINPUT124), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n955), .B1(new_n959), .B2(new_n961), .ZN(G1352gat));
  XOR2_X1   g761(.A(KEYINPUT125), .B(G204gat), .Z(new_n963));
  NAND3_X1  g762(.A1(new_n953), .A2(new_n720), .A3(new_n963), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n966), .B1(new_n965), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n957), .A2(new_n720), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  OAI22_X1  g770(.A1(new_n968), .A2(new_n969), .B1(new_n963), .B2(new_n971), .ZN(G1353gat));
  INV_X1    g771(.A(G211gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n953), .A2(new_n973), .A3(new_n632), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n632), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  INV_X1    g777(.A(G218gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n953), .A2(new_n979), .A3(new_n722), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n957), .A2(new_n722), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n980), .B1(new_n982), .B2(new_n979), .ZN(G1355gat));
endmodule


