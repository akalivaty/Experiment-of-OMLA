

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U554 ( .A(n604), .Z(n798) );
  AND2_X2 U555 ( .A1(n545), .A2(n544), .ZN(n613) );
  NOR2_X1 U556 ( .A1(n1023), .A2(n629), .ZN(n630) );
  XNOR2_X1 U557 ( .A(n528), .B(n527), .ZN(n702) );
  NOR2_X2 U558 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  AND2_X2 U559 ( .A1(G2105), .A2(G2104), .ZN(n999) );
  NOR2_X2 U560 ( .A1(n663), .A2(n662), .ZN(n664) );
  AND2_X2 U561 ( .A1(n631), .A2(n1023), .ZN(n633) );
  XNOR2_X2 U562 ( .A(n628), .B(KEYINPUT26), .ZN(n631) );
  XNOR2_X2 U563 ( .A(n537), .B(n536), .ZN(G160) );
  NOR2_X2 U564 ( .A1(n535), .A2(n534), .ZN(n537) );
  AND2_X1 U565 ( .A1(n726), .A2(n522), .ZN(n727) );
  NAND2_X1 U566 ( .A1(n640), .A2(n639), .ZN(n642) );
  XNOR2_X1 U567 ( .A(n548), .B(n547), .ZN(n604) );
  NOR2_X1 U568 ( .A1(G543), .A2(n551), .ZN(n548) );
  NAND2_X1 U569 ( .A1(n743), .A2(n523), .ZN(n744) );
  XOR2_X1 U570 ( .A(KEYINPUT0), .B(G543), .Z(n587) );
  XNOR2_X1 U571 ( .A(n526), .B(n525), .ZN(n530) );
  XNOR2_X1 U572 ( .A(n524), .B(KEYINPUT66), .ZN(n525) );
  AND2_X2 U573 ( .A1(n700), .A2(n616), .ZN(n636) );
  OR2_X1 U574 ( .A1(n739), .A2(n725), .ZN(n522) );
  XNOR2_X1 U575 ( .A(n614), .B(KEYINPUT64), .ZN(n700) );
  AND2_X1 U576 ( .A1(n742), .A2(n741), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n633), .A2(n632), .ZN(n635) );
  XNOR2_X1 U578 ( .A(n635), .B(n634), .ZN(n640) );
  INV_X1 U579 ( .A(KEYINPUT100), .ZN(n641) );
  INV_X1 U580 ( .A(KEYINPUT102), .ZN(n651) );
  INV_X1 U581 ( .A(n636), .ZN(n675) );
  NOR2_X2 U582 ( .A1(n613), .A2(G1384), .ZN(n614) );
  NAND2_X1 U583 ( .A1(n604), .A2(G66), .ZN(n606) );
  INV_X1 U584 ( .A(KEYINPUT17), .ZN(n527) );
  INV_X1 U585 ( .A(G651), .ZN(n551) );
  INV_X1 U586 ( .A(KEYINPUT1), .ZN(n547) );
  NOR2_X1 U587 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X2 U588 ( .A1(G651), .A2(n587), .ZN(n799) );
  BUF_X1 U589 ( .A(n702), .Z(n1003) );
  NOR2_X1 U590 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U591 ( .A1(n625), .A2(n624), .ZN(n1022) );
  BUF_X1 U592 ( .A(n613), .Z(G164) );
  INV_X1 U593 ( .A(G2104), .ZN(n531) );
  NOR2_X2 U594 ( .A1(G2105), .A2(n531), .ZN(n705) );
  NAND2_X1 U595 ( .A1(G101), .A2(n705), .ZN(n526) );
  INV_X1 U596 ( .A(KEYINPUT23), .ZN(n524) );
  NAND2_X1 U597 ( .A1(G137), .A2(n702), .ZN(n529) );
  NAND2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n535) );
  NAND2_X1 U599 ( .A1(G113), .A2(n999), .ZN(n533) );
  AND2_X2 U600 ( .A1(n531), .A2(G2105), .ZN(n1000) );
  NAND2_X1 U601 ( .A1(G125), .A2(n1000), .ZN(n532) );
  NAND2_X1 U602 ( .A1(n533), .A2(n532), .ZN(n534) );
  INV_X1 U603 ( .A(KEYINPUT65), .ZN(n536) );
  NAND2_X1 U604 ( .A1(G114), .A2(n999), .ZN(n538) );
  XNOR2_X1 U605 ( .A(KEYINPUT87), .B(n538), .ZN(n542) );
  NAND2_X1 U606 ( .A1(G102), .A2(n705), .ZN(n540) );
  NAND2_X1 U607 ( .A1(G126), .A2(n1000), .ZN(n539) );
  NAND2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n702), .A2(G138), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n543), .B(KEYINPUT88), .ZN(n544) );
  NAND2_X1 U612 ( .A1(G53), .A2(n799), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT70), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G65), .A2(n798), .ZN(n550) );
  NOR2_X2 U615 ( .A1(G651), .A2(G543), .ZN(n802) );
  NAND2_X1 U616 ( .A1(G91), .A2(n802), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n554) );
  NOR2_X2 U618 ( .A1(n587), .A2(n551), .ZN(n803) );
  NAND2_X1 U619 ( .A1(G78), .A2(n803), .ZN(n552) );
  XNOR2_X1 U620 ( .A(KEYINPUT69), .B(n552), .ZN(n553) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(G299) );
  NAND2_X1 U623 ( .A1(G64), .A2(n798), .ZN(n558) );
  NAND2_X1 U624 ( .A1(G52), .A2(n799), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n564) );
  NAND2_X1 U626 ( .A1(n803), .A2(G77), .ZN(n559) );
  XOR2_X1 U627 ( .A(KEYINPUT67), .B(n559), .Z(n561) );
  NAND2_X1 U628 ( .A1(n802), .A2(G90), .ZN(n560) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U630 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U631 ( .A1(n564), .A2(n563), .ZN(G171) );
  INV_X1 U632 ( .A(G171), .ZN(G301) );
  NAND2_X1 U633 ( .A1(n802), .A2(G89), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n565), .B(KEYINPUT4), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G76), .A2(n803), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n568), .B(KEYINPUT5), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G63), .A2(n798), .ZN(n570) );
  NAND2_X1 U639 ( .A1(G51), .A2(n799), .ZN(n569) );
  NAND2_X1 U640 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U641 ( .A(KEYINPUT6), .B(n571), .Z(n572) );
  NAND2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n574), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U644 ( .A(G168), .B(KEYINPUT8), .ZN(n575) );
  XNOR2_X1 U645 ( .A(n575), .B(KEYINPUT73), .ZN(G286) );
  NAND2_X1 U646 ( .A1(G62), .A2(n798), .ZN(n577) );
  NAND2_X1 U647 ( .A1(G50), .A2(n799), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U649 ( .A(KEYINPUT80), .B(n578), .ZN(n581) );
  NAND2_X1 U650 ( .A1(G75), .A2(n803), .ZN(n579) );
  XNOR2_X1 U651 ( .A(KEYINPUT81), .B(n579), .ZN(n580) );
  NOR2_X1 U652 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n802), .A2(G88), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(G303) );
  INV_X1 U655 ( .A(G303), .ZN(G166) );
  NAND2_X1 U656 ( .A1(G49), .A2(n799), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G74), .A2(G651), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U659 ( .A1(n798), .A2(n586), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n587), .A2(G87), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(G288) );
  NAND2_X1 U662 ( .A1(n799), .A2(G48), .ZN(n596) );
  NAND2_X1 U663 ( .A1(G61), .A2(n798), .ZN(n591) );
  NAND2_X1 U664 ( .A1(G86), .A2(n802), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n803), .A2(G73), .ZN(n592) );
  XOR2_X1 U667 ( .A(KEYINPUT2), .B(n592), .Z(n593) );
  NOR2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U670 ( .A(KEYINPUT79), .B(n597), .Z(G305) );
  NAND2_X1 U671 ( .A1(G85), .A2(n802), .ZN(n599) );
  NAND2_X1 U672 ( .A1(G72), .A2(n803), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G60), .A2(n798), .ZN(n601) );
  NAND2_X1 U675 ( .A1(G47), .A2(n799), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n602) );
  OR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(G290) );
  NAND2_X1 U678 ( .A1(G92), .A2(n802), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U680 ( .A(KEYINPUT72), .B(n607), .ZN(n611) );
  NAND2_X1 U681 ( .A1(G79), .A2(n803), .ZN(n609) );
  NAND2_X1 U682 ( .A1(G54), .A2(n799), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X2 U684 ( .A(KEYINPUT15), .B(n612), .Z(n1023) );
  NAND2_X1 U685 ( .A1(G160), .A2(G40), .ZN(n701) );
  INV_X1 U686 ( .A(n701), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n675), .A2(G1341), .ZN(n627) );
  NAND2_X1 U688 ( .A1(G56), .A2(n798), .ZN(n617) );
  XOR2_X1 U689 ( .A(KEYINPUT14), .B(n617), .Z(n623) );
  NAND2_X1 U690 ( .A1(n802), .A2(G81), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n618), .B(KEYINPUT12), .ZN(n620) );
  NAND2_X1 U692 ( .A1(G68), .A2(n803), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U694 ( .A(KEYINPUT13), .B(n621), .Z(n622) );
  NAND2_X1 U695 ( .A1(n799), .A2(G43), .ZN(n624) );
  INV_X1 U696 ( .A(n1022), .ZN(n626) );
  AND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n632) );
  NAND2_X1 U698 ( .A1(n636), .A2(G1996), .ZN(n628) );
  AND2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n629) );
  XOR2_X1 U700 ( .A(KEYINPUT101), .B(n630), .Z(n644) );
  INV_X1 U701 ( .A(KEYINPUT99), .ZN(n634) );
  NOR2_X1 U702 ( .A1(n636), .A2(G1348), .ZN(n638) );
  NOR2_X1 U703 ( .A1(G2067), .A2(n675), .ZN(n637) );
  NOR2_X1 U704 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U705 ( .A(n642), .B(n641), .ZN(n643) );
  NOR2_X1 U706 ( .A1(n644), .A2(n643), .ZN(n650) );
  NAND2_X1 U707 ( .A1(n675), .A2(G1956), .ZN(n647) );
  NAND2_X1 U708 ( .A1(n636), .A2(G2072), .ZN(n645) );
  XOR2_X1 U709 ( .A(KEYINPUT27), .B(n645), .Z(n646) );
  NAND2_X1 U710 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U711 ( .A(n648), .B(KEYINPUT98), .ZN(n653) );
  NOR2_X1 U712 ( .A1(n653), .A2(G299), .ZN(n649) );
  NOR2_X1 U713 ( .A1(n650), .A2(n649), .ZN(n652) );
  XNOR2_X1 U714 ( .A(n652), .B(n651), .ZN(n656) );
  NAND2_X1 U715 ( .A1(n653), .A2(G299), .ZN(n654) );
  XNOR2_X1 U716 ( .A(KEYINPUT28), .B(n654), .ZN(n655) );
  NAND2_X1 U717 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U718 ( .A(n657), .B(KEYINPUT29), .ZN(n663) );
  XOR2_X1 U719 ( .A(G1961), .B(KEYINPUT95), .Z(n947) );
  NOR2_X1 U720 ( .A1(n636), .A2(n947), .ZN(n658) );
  XOR2_X1 U721 ( .A(KEYINPUT96), .B(n658), .Z(n660) );
  XNOR2_X1 U722 ( .A(G2078), .B(KEYINPUT25), .ZN(n854) );
  NAND2_X1 U723 ( .A1(n636), .A2(n854), .ZN(n659) );
  NAND2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U725 ( .A(KEYINPUT97), .B(n661), .ZN(n668) );
  NOR2_X1 U726 ( .A1(G301), .A2(n668), .ZN(n662) );
  XNOR2_X1 U727 ( .A(n664), .B(KEYINPUT103), .ZN(n673) );
  NAND2_X1 U728 ( .A1(G8), .A2(n675), .ZN(n739) );
  NOR2_X1 U729 ( .A1(G1966), .A2(n739), .ZN(n688) );
  NOR2_X1 U730 ( .A1(G2084), .A2(n675), .ZN(n686) );
  NOR2_X1 U731 ( .A1(n688), .A2(n686), .ZN(n665) );
  NAND2_X1 U732 ( .A1(G8), .A2(n665), .ZN(n666) );
  XNOR2_X1 U733 ( .A(KEYINPUT30), .B(n666), .ZN(n667) );
  NOR2_X1 U734 ( .A1(G168), .A2(n667), .ZN(n670) );
  AND2_X1 U735 ( .A1(G301), .A2(n668), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U737 ( .A(KEYINPUT31), .B(n671), .Z(n672) );
  NAND2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X2 U739 ( .A(n674), .B(KEYINPUT104), .ZN(n690) );
  NAND2_X1 U740 ( .A1(n690), .A2(G286), .ZN(n683) );
  INV_X1 U741 ( .A(G8), .ZN(n681) );
  NOR2_X1 U742 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U743 ( .A(KEYINPUT105), .B(n676), .ZN(n679) );
  NOR2_X1 U744 ( .A1(G1971), .A2(n739), .ZN(n677) );
  NOR2_X1 U745 ( .A1(G166), .A2(n677), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  OR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n685) );
  INV_X1 U749 ( .A(KEYINPUT32), .ZN(n684) );
  XNOR2_X1 U750 ( .A(n685), .B(n684), .ZN(n729) );
  AND2_X1 U751 ( .A1(G8), .A2(n686), .ZN(n687) );
  NOR2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n730) );
  NAND2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n924) );
  AND2_X1 U755 ( .A1(n730), .A2(n924), .ZN(n691) );
  NAND2_X1 U756 ( .A1(n729), .A2(n691), .ZN(n698) );
  INV_X1 U757 ( .A(KEYINPUT33), .ZN(n696) );
  INV_X1 U758 ( .A(n924), .ZN(n693) );
  NOR2_X1 U759 ( .A1(G1976), .A2(G288), .ZN(n724) );
  NOR2_X1 U760 ( .A1(G1971), .A2(G303), .ZN(n692) );
  NOR2_X1 U761 ( .A1(n724), .A2(n692), .ZN(n925) );
  OR2_X1 U762 ( .A1(n693), .A2(n925), .ZN(n694) );
  OR2_X1 U763 ( .A1(n739), .A2(n694), .ZN(n695) );
  AND2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U766 ( .A(n699), .B(KEYINPUT106), .ZN(n728) );
  XOR2_X1 U767 ( .A(G1981), .B(G305), .Z(n914) );
  NOR2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n770) );
  XNOR2_X1 U769 ( .A(n770), .B(KEYINPUT94), .ZN(n721) );
  NAND2_X1 U770 ( .A1(G107), .A2(n999), .ZN(n704) );
  NAND2_X1 U771 ( .A1(G131), .A2(n1003), .ZN(n703) );
  NAND2_X1 U772 ( .A1(n704), .A2(n703), .ZN(n709) );
  BUF_X1 U773 ( .A(n705), .Z(n1005) );
  NAND2_X1 U774 ( .A1(G95), .A2(n1005), .ZN(n707) );
  NAND2_X1 U775 ( .A1(G119), .A2(n1000), .ZN(n706) );
  NAND2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U778 ( .A(KEYINPUT92), .B(n710), .Z(n994) );
  NAND2_X1 U779 ( .A1(G1991), .A2(n994), .ZN(n720) );
  NAND2_X1 U780 ( .A1(n1000), .A2(G129), .ZN(n717) );
  NAND2_X1 U781 ( .A1(G117), .A2(n999), .ZN(n712) );
  NAND2_X1 U782 ( .A1(G141), .A2(n1003), .ZN(n711) );
  NAND2_X1 U783 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U784 ( .A1(n1005), .A2(G105), .ZN(n713) );
  XOR2_X1 U785 ( .A(KEYINPUT38), .B(n713), .Z(n714) );
  NOR2_X1 U786 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U787 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U788 ( .A(KEYINPUT93), .B(n718), .Z(n996) );
  NAND2_X1 U789 ( .A1(G1996), .A2(n996), .ZN(n719) );
  NAND2_X1 U790 ( .A1(n720), .A2(n719), .ZN(n888) );
  NAND2_X1 U791 ( .A1(n721), .A2(n888), .ZN(n759) );
  XNOR2_X1 U792 ( .A(G1986), .B(G290), .ZN(n919) );
  NAND2_X1 U793 ( .A1(n770), .A2(n919), .ZN(n722) );
  XOR2_X1 U794 ( .A(KEYINPUT89), .B(n722), .Z(n723) );
  AND2_X1 U795 ( .A1(n759), .A2(n723), .ZN(n741) );
  AND2_X1 U796 ( .A1(n914), .A2(n741), .ZN(n726) );
  NAND2_X1 U797 ( .A1(n724), .A2(KEYINPUT33), .ZN(n725) );
  NAND2_X1 U798 ( .A1(n728), .A2(n727), .ZN(n745) );
  NAND2_X1 U799 ( .A1(n730), .A2(n729), .ZN(n738) );
  NAND2_X1 U800 ( .A1(G8), .A2(G166), .ZN(n731) );
  NOR2_X1 U801 ( .A1(G2090), .A2(n731), .ZN(n732) );
  XNOR2_X1 U802 ( .A(n732), .B(KEYINPUT107), .ZN(n736) );
  NOR2_X1 U803 ( .A1(G1981), .A2(G305), .ZN(n733) );
  XOR2_X1 U804 ( .A(n733), .B(KEYINPUT24), .Z(n734) );
  NOR2_X1 U805 ( .A1(n739), .A2(n734), .ZN(n740) );
  INV_X1 U806 ( .A(n740), .ZN(n735) );
  AND2_X1 U807 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n743) );
  OR2_X1 U809 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U810 ( .A1(n745), .A2(n744), .ZN(n757) );
  XNOR2_X1 U811 ( .A(G2067), .B(KEYINPUT37), .ZN(n746) );
  XNOR2_X1 U812 ( .A(n746), .B(KEYINPUT90), .ZN(n767) );
  NAND2_X1 U813 ( .A1(G104), .A2(n1005), .ZN(n748) );
  NAND2_X1 U814 ( .A1(G140), .A2(n1003), .ZN(n747) );
  NAND2_X1 U815 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U816 ( .A(KEYINPUT34), .B(n749), .ZN(n755) );
  NAND2_X1 U817 ( .A1(n1000), .A2(G128), .ZN(n750) );
  XOR2_X1 U818 ( .A(KEYINPUT91), .B(n750), .Z(n752) );
  NAND2_X1 U819 ( .A1(n999), .A2(G116), .ZN(n751) );
  NAND2_X1 U820 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U821 ( .A(KEYINPUT35), .B(n753), .Z(n754) );
  NOR2_X1 U822 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U823 ( .A(KEYINPUT36), .B(n756), .ZN(n1011) );
  NOR2_X1 U824 ( .A1(n767), .A2(n1011), .ZN(n896) );
  NAND2_X1 U825 ( .A1(n770), .A2(n896), .ZN(n765) );
  NAND2_X1 U826 ( .A1(n757), .A2(n765), .ZN(n758) );
  XNOR2_X1 U827 ( .A(n758), .B(KEYINPUT108), .ZN(n772) );
  NOR2_X1 U828 ( .A1(G1996), .A2(n996), .ZN(n893) );
  INV_X1 U829 ( .A(n759), .ZN(n762) );
  NOR2_X1 U830 ( .A1(G1986), .A2(G290), .ZN(n760) );
  NOR2_X1 U831 ( .A1(G1991), .A2(n994), .ZN(n898) );
  NOR2_X1 U832 ( .A1(n760), .A2(n898), .ZN(n761) );
  NOR2_X1 U833 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U834 ( .A1(n893), .A2(n763), .ZN(n764) );
  XNOR2_X1 U835 ( .A(n764), .B(KEYINPUT39), .ZN(n766) );
  NAND2_X1 U836 ( .A1(n766), .A2(n765), .ZN(n768) );
  NAND2_X1 U837 ( .A1(n767), .A2(n1011), .ZN(n887) );
  NAND2_X1 U838 ( .A1(n768), .A2(n887), .ZN(n769) );
  NAND2_X1 U839 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U840 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U841 ( .A(n773), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U842 ( .A(G120), .ZN(G236) );
  INV_X1 U843 ( .A(G69), .ZN(G235) );
  INV_X1 U844 ( .A(G108), .ZN(G238) );
  NAND2_X1 U845 ( .A1(G94), .A2(G452), .ZN(n774) );
  XOR2_X1 U846 ( .A(KEYINPUT68), .B(n774), .Z(G173) );
  XOR2_X1 U847 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n776) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n775) );
  XNOR2_X1 U849 ( .A(n776), .B(n775), .ZN(G223) );
  INV_X1 U850 ( .A(G223), .ZN(n841) );
  NAND2_X1 U851 ( .A1(n841), .A2(G567), .ZN(n777) );
  XOR2_X1 U852 ( .A(KEYINPUT11), .B(n777), .Z(G234) );
  INV_X1 U853 ( .A(G860), .ZN(n810) );
  OR2_X1 U854 ( .A1(n1022), .A2(n810), .ZN(G153) );
  NAND2_X1 U855 ( .A1(G868), .A2(G301), .ZN(n779) );
  OR2_X1 U856 ( .A1(n1023), .A2(G868), .ZN(n778) );
  NAND2_X1 U857 ( .A1(n779), .A2(n778), .ZN(G284) );
  INV_X1 U858 ( .A(G868), .ZN(n822) );
  NOR2_X1 U859 ( .A1(G286), .A2(n822), .ZN(n781) );
  NOR2_X1 U860 ( .A1(G868), .A2(G299), .ZN(n780) );
  NOR2_X1 U861 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U862 ( .A(KEYINPUT74), .B(n782), .ZN(G297) );
  NAND2_X1 U863 ( .A1(G559), .A2(n810), .ZN(n783) );
  XOR2_X1 U864 ( .A(KEYINPUT75), .B(n783), .Z(n784) );
  NAND2_X1 U865 ( .A1(n784), .A2(n1023), .ZN(n785) );
  XNOR2_X1 U866 ( .A(n785), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U867 ( .A1(G868), .A2(n1022), .ZN(n788) );
  NAND2_X1 U868 ( .A1(n1023), .A2(G868), .ZN(n786) );
  NOR2_X1 U869 ( .A1(G559), .A2(n786), .ZN(n787) );
  NOR2_X1 U870 ( .A1(n788), .A2(n787), .ZN(G282) );
  XOR2_X1 U871 ( .A(G2100), .B(KEYINPUT76), .Z(n797) );
  NAND2_X1 U872 ( .A1(G111), .A2(n999), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G135), .A2(n1003), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U875 ( .A1(n1000), .A2(G123), .ZN(n791) );
  XOR2_X1 U876 ( .A(KEYINPUT18), .B(n791), .Z(n792) );
  NOR2_X1 U877 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U878 ( .A1(n1005), .A2(G99), .ZN(n794) );
  NAND2_X1 U879 ( .A1(n795), .A2(n794), .ZN(n1016) );
  XOR2_X1 U880 ( .A(G2096), .B(n1016), .Z(n796) );
  NAND2_X1 U881 ( .A1(n797), .A2(n796), .ZN(G156) );
  NAND2_X1 U882 ( .A1(G67), .A2(n798), .ZN(n801) );
  NAND2_X1 U883 ( .A1(G55), .A2(n799), .ZN(n800) );
  NAND2_X1 U884 ( .A1(n801), .A2(n800), .ZN(n808) );
  NAND2_X1 U885 ( .A1(G93), .A2(n802), .ZN(n805) );
  NAND2_X1 U886 ( .A1(G80), .A2(n803), .ZN(n804) );
  NAND2_X1 U887 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U888 ( .A(KEYINPUT77), .B(n806), .Z(n807) );
  OR2_X1 U889 ( .A1(n808), .A2(n807), .ZN(n823) );
  XNOR2_X1 U890 ( .A(n823), .B(KEYINPUT78), .ZN(n812) );
  NAND2_X1 U891 ( .A1(G559), .A2(n1023), .ZN(n809) );
  XOR2_X1 U892 ( .A(n1022), .B(n809), .Z(n819) );
  NAND2_X1 U893 ( .A1(n819), .A2(n810), .ZN(n811) );
  XNOR2_X1 U894 ( .A(n812), .B(n811), .ZN(G145) );
  XNOR2_X1 U895 ( .A(KEYINPUT19), .B(G303), .ZN(n813) );
  XNOR2_X1 U896 ( .A(n813), .B(G288), .ZN(n814) );
  XNOR2_X1 U897 ( .A(KEYINPUT82), .B(n814), .ZN(n816) );
  XOR2_X1 U898 ( .A(G305), .B(n823), .Z(n815) );
  XNOR2_X1 U899 ( .A(n816), .B(n815), .ZN(n817) );
  XNOR2_X1 U900 ( .A(n817), .B(G290), .ZN(n818) );
  XNOR2_X1 U901 ( .A(n818), .B(G299), .ZN(n1021) );
  XNOR2_X1 U902 ( .A(n819), .B(n1021), .ZN(n820) );
  XNOR2_X1 U903 ( .A(KEYINPUT83), .B(n820), .ZN(n821) );
  NOR2_X1 U904 ( .A1(n822), .A2(n821), .ZN(n825) );
  NOR2_X1 U905 ( .A1(G868), .A2(n823), .ZN(n824) );
  NOR2_X1 U906 ( .A1(n825), .A2(n824), .ZN(G295) );
  NAND2_X1 U907 ( .A1(G2078), .A2(G2084), .ZN(n826) );
  XOR2_X1 U908 ( .A(KEYINPUT20), .B(n826), .Z(n827) );
  NAND2_X1 U909 ( .A1(G2090), .A2(n827), .ZN(n828) );
  XNOR2_X1 U910 ( .A(KEYINPUT21), .B(n828), .ZN(n829) );
  NAND2_X1 U911 ( .A1(n829), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U912 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U913 ( .A1(G132), .A2(G82), .ZN(n830) );
  XNOR2_X1 U914 ( .A(n830), .B(KEYINPUT84), .ZN(n831) );
  XNOR2_X1 U915 ( .A(n831), .B(KEYINPUT22), .ZN(n832) );
  NOR2_X1 U916 ( .A1(G218), .A2(n832), .ZN(n833) );
  NAND2_X1 U917 ( .A1(G96), .A2(n833), .ZN(n969) );
  NAND2_X1 U918 ( .A1(n969), .A2(G2106), .ZN(n839) );
  NOR2_X1 U919 ( .A1(G235), .A2(G236), .ZN(n834) );
  XNOR2_X1 U920 ( .A(n834), .B(KEYINPUT85), .ZN(n835) );
  NOR2_X1 U921 ( .A1(G238), .A2(n835), .ZN(n836) );
  NAND2_X1 U922 ( .A1(n836), .A2(G57), .ZN(n837) );
  XNOR2_X1 U923 ( .A(n837), .B(KEYINPUT86), .ZN(n970) );
  NAND2_X1 U924 ( .A1(n970), .A2(G567), .ZN(n838) );
  NAND2_X1 U925 ( .A1(n839), .A2(n838), .ZN(n971) );
  NAND2_X1 U926 ( .A1(G483), .A2(G661), .ZN(n840) );
  NOR2_X1 U927 ( .A1(n971), .A2(n840), .ZN(n843) );
  NAND2_X1 U928 ( .A1(n843), .A2(G36), .ZN(G176) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n841), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n842) );
  NAND2_X1 U931 ( .A1(G661), .A2(n842), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U933 ( .A1(n844), .A2(n843), .ZN(n845) );
  XOR2_X1 U934 ( .A(KEYINPUT109), .B(n845), .Z(G188) );
  NAND2_X1 U936 ( .A1(G124), .A2(n1000), .ZN(n846) );
  XNOR2_X1 U937 ( .A(n846), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U938 ( .A1(n999), .A2(G112), .ZN(n847) );
  NAND2_X1 U939 ( .A1(n848), .A2(n847), .ZN(n852) );
  NAND2_X1 U940 ( .A1(G100), .A2(n1005), .ZN(n850) );
  NAND2_X1 U941 ( .A1(G136), .A2(n1003), .ZN(n849) );
  NAND2_X1 U942 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U943 ( .A1(n852), .A2(n851), .ZN(G162) );
  XNOR2_X1 U944 ( .A(G2090), .B(G35), .ZN(n868) );
  XOR2_X1 U945 ( .A(KEYINPUT119), .B(G27), .Z(n853) );
  XNOR2_X1 U946 ( .A(n854), .B(n853), .ZN(n861) );
  XOR2_X1 U947 ( .A(G2067), .B(G26), .Z(n857) );
  XOR2_X1 U948 ( .A(G32), .B(KEYINPUT120), .Z(n855) );
  XNOR2_X1 U949 ( .A(G1996), .B(n855), .ZN(n856) );
  NAND2_X1 U950 ( .A1(n857), .A2(n856), .ZN(n859) );
  XNOR2_X1 U951 ( .A(G33), .B(G2072), .ZN(n858) );
  NOR2_X1 U952 ( .A1(n859), .A2(n858), .ZN(n860) );
  NAND2_X1 U953 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U954 ( .A(KEYINPUT121), .B(n862), .ZN(n863) );
  NAND2_X1 U955 ( .A1(n863), .A2(G28), .ZN(n865) );
  XNOR2_X1 U956 ( .A(G25), .B(G1991), .ZN(n864) );
  NOR2_X1 U957 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U958 ( .A(KEYINPUT53), .B(n866), .ZN(n867) );
  NOR2_X1 U959 ( .A1(n868), .A2(n867), .ZN(n871) );
  XOR2_X1 U960 ( .A(G2084), .B(KEYINPUT54), .Z(n869) );
  XNOR2_X1 U961 ( .A(G34), .B(n869), .ZN(n870) );
  NAND2_X1 U962 ( .A1(n871), .A2(n870), .ZN(n908) );
  NOR2_X1 U963 ( .A1(G29), .A2(KEYINPUT55), .ZN(n872) );
  NAND2_X1 U964 ( .A1(n908), .A2(n872), .ZN(n873) );
  NAND2_X1 U965 ( .A1(G11), .A2(n873), .ZN(n913) );
  XOR2_X1 U966 ( .A(G164), .B(G2078), .Z(n874) );
  XNOR2_X1 U967 ( .A(KEYINPUT118), .B(n874), .ZN(n885) );
  NAND2_X1 U968 ( .A1(G103), .A2(n1005), .ZN(n876) );
  NAND2_X1 U969 ( .A1(G139), .A2(n1003), .ZN(n875) );
  NAND2_X1 U970 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U971 ( .A(KEYINPUT114), .B(n877), .ZN(n883) );
  NAND2_X1 U972 ( .A1(n999), .A2(G115), .ZN(n878) );
  XOR2_X1 U973 ( .A(KEYINPUT115), .B(n878), .Z(n880) );
  NAND2_X1 U974 ( .A1(n1000), .A2(G127), .ZN(n879) );
  NAND2_X1 U975 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U976 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U977 ( .A1(n883), .A2(n882), .ZN(n1015) );
  XOR2_X1 U978 ( .A(G2072), .B(n1015), .Z(n884) );
  NOR2_X1 U979 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U980 ( .A(KEYINPUT50), .B(n886), .ZN(n891) );
  INV_X1 U981 ( .A(n887), .ZN(n889) );
  NOR2_X1 U982 ( .A1(n889), .A2(n888), .ZN(n890) );
  NAND2_X1 U983 ( .A1(n891), .A2(n890), .ZN(n904) );
  XOR2_X1 U984 ( .A(G2090), .B(G162), .Z(n892) );
  NOR2_X1 U985 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U986 ( .A(n894), .B(KEYINPUT51), .ZN(n895) );
  NOR2_X1 U987 ( .A1(n896), .A2(n895), .ZN(n902) );
  XNOR2_X1 U988 ( .A(G160), .B(G2084), .ZN(n897) );
  NAND2_X1 U989 ( .A1(n897), .A2(n1016), .ZN(n899) );
  NOR2_X1 U990 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U991 ( .A(KEYINPUT117), .B(n900), .Z(n901) );
  NAND2_X1 U992 ( .A1(n902), .A2(n901), .ZN(n903) );
  NOR2_X1 U993 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U994 ( .A(KEYINPUT52), .B(n905), .ZN(n906) );
  INV_X1 U995 ( .A(KEYINPUT55), .ZN(n909) );
  NAND2_X1 U996 ( .A1(n906), .A2(n909), .ZN(n907) );
  NAND2_X1 U997 ( .A1(n907), .A2(G29), .ZN(n911) );
  OR2_X1 U998 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U999 ( .A1(n911), .A2(n910), .ZN(n912) );
  NOR2_X1 U1000 ( .A1(n913), .A2(n912), .ZN(n967) );
  XNOR2_X1 U1001 ( .A(G16), .B(KEYINPUT56), .ZN(n937) );
  XNOR2_X1 U1002 ( .A(G1966), .B(G168), .ZN(n915) );
  NAND2_X1 U1003 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1004 ( .A(n916), .B(KEYINPUT57), .ZN(n935) );
  XNOR2_X1 U1005 ( .A(G1348), .B(n1023), .ZN(n917) );
  XNOR2_X1 U1006 ( .A(n917), .B(KEYINPUT122), .ZN(n921) );
  XNOR2_X1 U1007 ( .A(G1956), .B(G299), .ZN(n918) );
  NOR2_X1 U1008 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1009 ( .A1(n921), .A2(n920), .ZN(n923) );
  XNOR2_X1 U1010 ( .A(G1341), .B(n1022), .ZN(n922) );
  NOR2_X1 U1011 ( .A1(n923), .A2(n922), .ZN(n931) );
  NAND2_X1 U1012 ( .A1(n925), .A2(n924), .ZN(n928) );
  INV_X1 U1013 ( .A(G1971), .ZN(n926) );
  NOR2_X1 U1014 ( .A1(G166), .A2(n926), .ZN(n927) );
  NOR2_X1 U1015 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1016 ( .A(KEYINPUT123), .B(n929), .Z(n930) );
  NAND2_X1 U1017 ( .A1(n931), .A2(n930), .ZN(n933) );
  XNOR2_X1 U1018 ( .A(G1961), .B(G301), .ZN(n932) );
  NOR2_X1 U1019 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1020 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1021 ( .A1(n937), .A2(n936), .ZN(n964) );
  INV_X1 U1022 ( .A(G16), .ZN(n962) );
  XNOR2_X1 U1023 ( .A(G1348), .B(KEYINPUT59), .ZN(n938) );
  XNOR2_X1 U1024 ( .A(n938), .B(G4), .ZN(n942) );
  XNOR2_X1 U1025 ( .A(G1956), .B(G20), .ZN(n940) );
  XNOR2_X1 U1026 ( .A(G1981), .B(G6), .ZN(n939) );
  NOR2_X1 U1027 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1028 ( .A1(n942), .A2(n941), .ZN(n945) );
  XOR2_X1 U1029 ( .A(KEYINPUT125), .B(G1341), .Z(n943) );
  XNOR2_X1 U1030 ( .A(G19), .B(n943), .ZN(n944) );
  NOR2_X1 U1031 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1032 ( .A(KEYINPUT60), .B(n946), .ZN(n957) );
  XNOR2_X1 U1033 ( .A(n947), .B(G5), .ZN(n948) );
  XNOR2_X1 U1034 ( .A(n948), .B(KEYINPUT124), .ZN(n955) );
  XNOR2_X1 U1035 ( .A(G1986), .B(G24), .ZN(n950) );
  XNOR2_X1 U1036 ( .A(G1971), .B(G22), .ZN(n949) );
  NOR2_X1 U1037 ( .A1(n950), .A2(n949), .ZN(n952) );
  XOR2_X1 U1038 ( .A(G1976), .B(G23), .Z(n951) );
  NAND2_X1 U1039 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1040 ( .A(KEYINPUT58), .B(n953), .ZN(n954) );
  NOR2_X1 U1041 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1042 ( .A1(n957), .A2(n956), .ZN(n959) );
  XNOR2_X1 U1043 ( .A(G21), .B(G1966), .ZN(n958) );
  NOR2_X1 U1044 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1045 ( .A(KEYINPUT61), .B(n960), .ZN(n961) );
  NAND2_X1 U1046 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1047 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1048 ( .A(KEYINPUT126), .B(n965), .Z(n966) );
  NAND2_X1 U1049 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1050 ( .A(KEYINPUT62), .B(n968), .Z(G311) );
  XNOR2_X1 U1051 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1052 ( .A(G132), .ZN(G219) );
  INV_X1 U1053 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1054 ( .A1(n970), .A2(n969), .ZN(G325) );
  INV_X1 U1055 ( .A(G325), .ZN(G261) );
  INV_X1 U1056 ( .A(n971), .ZN(G319) );
  XOR2_X1 U1057 ( .A(G2096), .B(G2100), .Z(n973) );
  XNOR2_X1 U1058 ( .A(G2072), .B(G2090), .ZN(n972) );
  XNOR2_X1 U1059 ( .A(n973), .B(n972), .ZN(n977) );
  XOR2_X1 U1060 ( .A(G2678), .B(KEYINPUT42), .Z(n975) );
  XNOR2_X1 U1061 ( .A(G2067), .B(KEYINPUT43), .ZN(n974) );
  XNOR2_X1 U1062 ( .A(n975), .B(n974), .ZN(n976) );
  XOR2_X1 U1063 ( .A(n977), .B(n976), .Z(n979) );
  XNOR2_X1 U1064 ( .A(G2078), .B(G2084), .ZN(n978) );
  XNOR2_X1 U1065 ( .A(n979), .B(n978), .ZN(G227) );
  XOR2_X1 U1066 ( .A(KEYINPUT41), .B(G2474), .Z(n981) );
  XNOR2_X1 U1067 ( .A(G1961), .B(G1976), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(n981), .B(n980), .ZN(n991) );
  XOR2_X1 U1069 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n983) );
  XNOR2_X1 U1070 ( .A(G1996), .B(G1966), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(n983), .B(n982), .ZN(n987) );
  XOR2_X1 U1072 ( .A(G1981), .B(G1971), .Z(n985) );
  XNOR2_X1 U1073 ( .A(G1991), .B(G1956), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(n985), .B(n984), .ZN(n986) );
  XOR2_X1 U1075 ( .A(n987), .B(n986), .Z(n989) );
  XNOR2_X1 U1076 ( .A(G1986), .B(KEYINPUT112), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(n989), .B(n988), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(n991), .B(n990), .ZN(G229) );
  XOR2_X1 U1079 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n993) );
  XNOR2_X1 U1080 ( .A(G162), .B(KEYINPUT116), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n993), .B(n992), .ZN(n998) );
  XOR2_X1 U1082 ( .A(G160), .B(n994), .Z(n995) );
  XNOR2_X1 U1083 ( .A(n996), .B(n995), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(n998), .B(n997), .ZN(n1014) );
  NAND2_X1 U1085 ( .A1(G118), .A2(n999), .ZN(n1002) );
  NAND2_X1 U1086 ( .A1(G130), .A2(n1000), .ZN(n1001) );
  NAND2_X1 U1087 ( .A1(n1002), .A2(n1001), .ZN(n1010) );
  NAND2_X1 U1088 ( .A1(n1003), .A2(G142), .ZN(n1004) );
  XOR2_X1 U1089 ( .A(KEYINPUT113), .B(n1004), .Z(n1007) );
  NAND2_X1 U1090 ( .A1(n1005), .A2(G106), .ZN(n1006) );
  NAND2_X1 U1091 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1092 ( .A(n1008), .B(KEYINPUT45), .Z(n1009) );
  NOR2_X1 U1093 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1094 ( .A(n1012), .B(n1011), .ZN(n1013) );
  XNOR2_X1 U1095 ( .A(n1014), .B(n1013), .ZN(n1019) );
  XNOR2_X1 U1096 ( .A(G164), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1097 ( .A(n1017), .B(n1016), .ZN(n1018) );
  XOR2_X1 U1098 ( .A(n1019), .B(n1018), .Z(n1020) );
  NOR2_X1 U1099 ( .A1(G37), .A2(n1020), .ZN(G395) );
  XNOR2_X1 U1100 ( .A(n1022), .B(n1021), .ZN(n1025) );
  XNOR2_X1 U1101 ( .A(G171), .B(n1023), .ZN(n1024) );
  XNOR2_X1 U1102 ( .A(n1025), .B(n1024), .ZN(n1026) );
  XOR2_X1 U1103 ( .A(G286), .B(n1026), .Z(n1027) );
  NOR2_X1 U1104 ( .A1(G37), .A2(n1027), .ZN(G397) );
  XOR2_X1 U1105 ( .A(G2446), .B(G2451), .Z(n1029) );
  XNOR2_X1 U1106 ( .A(G1348), .B(G2430), .ZN(n1028) );
  XNOR2_X1 U1107 ( .A(n1029), .B(n1028), .ZN(n1035) );
  XOR2_X1 U1108 ( .A(G2443), .B(G2438), .Z(n1031) );
  XNOR2_X1 U1109 ( .A(G2454), .B(G2435), .ZN(n1030) );
  XNOR2_X1 U1110 ( .A(n1031), .B(n1030), .ZN(n1033) );
  XOR2_X1 U1111 ( .A(G1341), .B(G2427), .Z(n1032) );
  XNOR2_X1 U1112 ( .A(n1033), .B(n1032), .ZN(n1034) );
  XOR2_X1 U1113 ( .A(n1035), .B(n1034), .Z(n1036) );
  NAND2_X1 U1114 ( .A1(G14), .A2(n1036), .ZN(n1042) );
  NAND2_X1 U1115 ( .A1(G319), .A2(n1042), .ZN(n1039) );
  NOR2_X1 U1116 ( .A1(G227), .A2(G229), .ZN(n1037) );
  XNOR2_X1 U1117 ( .A(KEYINPUT49), .B(n1037), .ZN(n1038) );
  NOR2_X1 U1118 ( .A1(n1039), .A2(n1038), .ZN(n1041) );
  NOR2_X1 U1119 ( .A1(G395), .A2(G397), .ZN(n1040) );
  NAND2_X1 U1120 ( .A1(n1041), .A2(n1040), .ZN(G225) );
  INV_X1 U1121 ( .A(G225), .ZN(G308) );
  INV_X1 U1122 ( .A(G57), .ZN(G237) );
  INV_X1 U1123 ( .A(G96), .ZN(G221) );
  INV_X1 U1124 ( .A(n1042), .ZN(G401) );
endmodule

