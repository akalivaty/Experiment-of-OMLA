//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1300, new_n1301, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n207), .B1(new_n213), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n207), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n221), .B(new_n224), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT65), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n215), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT68), .B(G50), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n245), .B(KEYINPUT71), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT69), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT70), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n226), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n226), .A2(new_n256), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n253), .A2(new_n254), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n258), .B1(G20), .B2(new_n203), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n225), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G13), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n264), .A2(new_n226), .A3(G1), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n261), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(G50), .A3(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n264), .A2(G1), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G20), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n269), .B1(G50), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n273), .B(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n282), .A3(G1698), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT73), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT73), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(G1698), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n279), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n285), .A2(G222), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G77), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n285), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n278), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n277), .A2(G274), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n277), .A2(new_n295), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT72), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT72), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n277), .A2(new_n299), .A3(new_n295), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n296), .B1(new_n301), .B2(G226), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n293), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G190), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n275), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT79), .ZN(new_n307));
  XNOR2_X1  g0107(.A(KEYINPUT78), .B(G200), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT10), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n275), .A2(new_n305), .ZN(new_n314));
  INV_X1    g0114(.A(new_n310), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n273), .B1(new_n303), .B2(new_n319), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n320), .A2(KEYINPUT74), .ZN(new_n321));
  INV_X1    g0121(.A(G179), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n304), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(KEYINPUT74), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n216), .A2(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(G226), .B2(G1698), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n280), .A2(new_n282), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n327), .A2(new_n328), .B1(new_n256), .B2(new_n217), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n278), .ZN(new_n330));
  INV_X1    g0130(.A(new_n295), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(new_n277), .A3(G274), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n210), .B1(new_n298), .B2(new_n300), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT13), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n334), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n296), .B1(new_n329), .B2(new_n278), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT13), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT14), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT80), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n333), .B2(new_n334), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT80), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT13), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(G179), .A3(new_n339), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT14), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n340), .A2(new_n348), .A3(G169), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n342), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT77), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n262), .A2(new_n271), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT77), .B1(new_n265), .B2(new_n261), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n267), .B2(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G68), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G20), .A2(G33), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(G50), .B1(G20), .B2(new_n209), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n291), .B2(new_n254), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n359), .A2(new_n261), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n360), .A2(KEYINPUT11), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n265), .A2(new_n209), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT12), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(KEYINPUT11), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n356), .A2(new_n361), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n350), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(G200), .B2(new_n340), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n346), .A2(G190), .A3(new_n339), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n318), .A2(new_n325), .A3(new_n366), .A4(new_n369), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n253), .A2(new_n257), .B1(new_n226), .B2(new_n291), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT15), .B(G87), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n254), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n261), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n265), .A2(new_n291), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n355), .B2(G77), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n301), .A2(G244), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT75), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n332), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n210), .B1(new_n284), .B2(new_n287), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n285), .A2(G232), .A3(new_n289), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n211), .B2(new_n285), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n278), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G244), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n298), .B2(new_n300), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT75), .B1(new_n386), .B2(new_n296), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n380), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT76), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT76), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n380), .A2(new_n387), .A3(new_n390), .A4(new_n384), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n377), .B1(new_n392), .B2(new_n308), .ZN(new_n393));
  INV_X1    g0193(.A(G190), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n394), .B1(new_n389), .B2(new_n391), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n377), .B1(new_n392), .B2(new_n322), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n389), .A2(new_n319), .A3(new_n391), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n253), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n268), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n403), .A2(new_n266), .B1(new_n265), .B2(new_n253), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  INV_X1    g0206(.A(G159), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT81), .B1(new_n257), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT81), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n357), .A2(new_n409), .A3(G159), .ZN(new_n410));
  XNOR2_X1  g0210(.A(G58), .B(G68), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n408), .A2(new_n410), .B1(new_n411), .B2(G20), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT82), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n280), .A2(new_n282), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(G20), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n256), .A2(KEYINPUT82), .A3(KEYINPUT3), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n415), .B1(new_n285), .B2(G20), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n209), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n412), .B1(new_n420), .B2(KEYINPUT83), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT83), .ZN(new_n422));
  AOI211_X1 g0222(.A(new_n422), .B(new_n209), .C1(new_n418), .C2(new_n419), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n406), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n408), .A2(new_n410), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n411), .A2(G20), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n226), .A2(KEYINPUT7), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n419), .B1(new_n285), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n427), .B1(new_n429), .B2(G68), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n262), .B1(new_n430), .B2(KEYINPUT16), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n405), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n279), .A2(new_n289), .ZN(new_n433));
  INV_X1    g0233(.A(G226), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G1698), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n280), .A2(new_n433), .A3(new_n282), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G87), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n278), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n277), .A2(G232), .A3(new_n295), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n439), .A2(new_n394), .A3(new_n332), .A4(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G200), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n332), .A2(new_n440), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n277), .B1(new_n436), .B2(new_n437), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n441), .A2(KEYINPUT84), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT84), .B1(new_n441), .B2(new_n445), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n432), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT17), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n443), .A2(new_n444), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G179), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n319), .B2(new_n452), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT18), .B1(new_n432), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT18), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n428), .B1(new_n280), .B2(new_n282), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n328), .A2(new_n226), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(new_n415), .ZN(new_n460));
  OAI211_X1 g0260(.A(KEYINPUT16), .B(new_n412), .C1(new_n460), .C2(new_n209), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n261), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n417), .A2(new_n416), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n459), .A2(new_n415), .B1(new_n463), .B2(new_n414), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n422), .B1(new_n464), .B2(new_n209), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n420), .A2(KEYINPUT83), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n466), .A3(new_n412), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n462), .B1(new_n467), .B2(new_n406), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n457), .B(new_n454), .C1(new_n468), .C2(new_n405), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n432), .A2(KEYINPUT17), .A3(new_n448), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n451), .A2(new_n456), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n400), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n370), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n267), .A2(G45), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n225), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n475), .A2(new_n477), .B1(new_n478), .B2(new_n276), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G257), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n475), .A2(new_n477), .A3(G274), .A4(new_n277), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n280), .A2(new_n282), .A3(G250), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G1698), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G1698), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(new_n280), .A3(new_n282), .A4(G244), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G283), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n280), .A2(new_n282), .A3(G244), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n486), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n485), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n277), .B1(new_n493), .B2(KEYINPUT87), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT87), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n485), .A2(new_n490), .A3(new_n495), .A4(new_n492), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n482), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(KEYINPUT88), .A3(G190), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT88), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n492), .A2(new_n488), .A3(new_n489), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n289), .B1(new_n483), .B2(KEYINPUT4), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT87), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(new_n496), .A3(new_n278), .ZN(new_n503));
  INV_X1    g0303(.A(new_n482), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n499), .B1(new_n505), .B2(new_n394), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(G200), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n267), .A2(G33), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT86), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n266), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT85), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n265), .B2(new_n217), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n271), .A2(KEYINPUT85), .A3(G97), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n510), .A2(new_n217), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n418), .A2(new_n419), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n257), .A2(new_n291), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n217), .A2(new_n211), .ZN(new_n519));
  NOR2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n211), .A2(KEYINPUT6), .A3(G97), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n517), .B1(new_n523), .B2(G20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n514), .B1(new_n525), .B2(new_n261), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n498), .A2(new_n506), .A3(new_n507), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n526), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n503), .A2(new_n322), .A3(new_n504), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n528), .B(new_n529), .C1(new_n497), .C2(G169), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n210), .A2(G1698), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(new_n280), .A3(new_n282), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT89), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n280), .A2(new_n282), .A3(G244), .A4(G1698), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT89), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n531), .A2(new_n280), .A3(new_n282), .A4(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n278), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n476), .A2(G250), .ZN(new_n540));
  OAI22_X1  g0340(.A1(new_n294), .A2(new_n476), .B1(new_n278), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n226), .ZN(new_n545));
  INV_X1    g0345(.A(G87), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n520), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n280), .A2(new_n282), .A3(new_n226), .A4(G68), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n254), .B2(new_n217), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n261), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n372), .A2(new_n265), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n510), .ZN(new_n556));
  INV_X1    g0356(.A(new_n372), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n543), .A2(new_n319), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n541), .B1(new_n538), .B2(new_n278), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n322), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n543), .A2(new_n309), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n509), .A2(G87), .A3(new_n266), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n553), .A2(new_n554), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n560), .B2(G190), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n559), .A2(new_n561), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n527), .A2(new_n530), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n475), .A2(new_n477), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(G270), .A3(new_n277), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n481), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(G303), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n283), .A2(new_n212), .B1(new_n285), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT90), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n289), .A2(G257), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n328), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n285), .A2(KEYINPUT90), .A3(G257), .A4(new_n289), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n571), .B1(new_n578), .B2(new_n277), .ZN(new_n579));
  INV_X1    g0379(.A(G116), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n270), .A2(G20), .A3(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n260), .A2(new_n225), .B1(G20), .B2(new_n580), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n489), .B(new_n226), .C1(G33), .C2(new_n217), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n582), .A2(KEYINPUT20), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT20), .B1(new_n582), .B2(new_n583), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n509), .A2(G116), .ZN(new_n586));
  OAI221_X1 g0386(.A(new_n581), .B1(new_n584), .B2(new_n585), .C1(new_n354), .C2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n579), .A2(new_n587), .A3(G169), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n576), .A2(new_n577), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n280), .A2(new_n282), .A3(G1698), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n591), .A2(G264), .B1(G303), .B2(new_n328), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n277), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n593), .A2(new_n322), .A3(new_n570), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n587), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT91), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT91), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n597), .A3(new_n587), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n587), .B1(new_n579), .B2(G200), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n394), .B2(new_n579), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n589), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g0402(.A(KEYINPUT92), .B(KEYINPUT22), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n280), .A2(new_n282), .A3(new_n226), .A4(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n285), .A2(new_n603), .A3(new_n226), .A4(G87), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT24), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n534), .A2(G20), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT23), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n226), .B2(G107), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n211), .A2(KEYINPUT23), .A3(G20), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n609), .B1(new_n608), .B2(new_n614), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n261), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n271), .A2(G107), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n618), .A2(KEYINPUT25), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(KEYINPUT25), .ZN(new_n620));
  AOI22_X1  g0420(.A1(G107), .A2(new_n556), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n218), .A2(G1698), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(G250), .B2(G1698), .ZN(new_n624));
  INV_X1    g0424(.A(G294), .ZN(new_n625));
  OAI22_X1  g0425(.A1(new_n624), .A2(new_n328), .B1(new_n256), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n278), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n479), .A2(G264), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n481), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G200), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n394), .B2(new_n629), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n622), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n626), .A2(new_n278), .B1(new_n479), .B2(G264), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n319), .B1(new_n634), .B2(new_n481), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(KEYINPUT93), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n629), .A2(KEYINPUT93), .A3(G169), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(G179), .A3(new_n481), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n622), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n602), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n474), .A2(new_n567), .A3(new_n642), .ZN(G372));
  INV_X1    g0443(.A(new_n325), .ZN(new_n644));
  INV_X1    g0444(.A(new_n369), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n366), .B1(new_n399), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n451), .A2(new_n470), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n456), .A2(new_n469), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT95), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n456), .A2(KEYINPUT95), .A3(new_n469), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n644), .B1(new_n654), .B2(new_n318), .ZN(new_n655));
  INV_X1    g0455(.A(new_n474), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n589), .A2(new_n640), .A3(new_n599), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n633), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n527), .A2(new_n530), .A3(new_n566), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n553), .B(new_n554), .C1(new_n510), .C2(new_n372), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n560), .B2(G169), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n560), .A2(new_n322), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n503), .A2(new_n322), .A3(new_n504), .ZN(new_n666));
  AOI21_X1  g0466(.A(G169), .B1(new_n503), .B2(new_n504), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n666), .A2(new_n667), .A3(new_n526), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT26), .B1(new_n668), .B2(new_n566), .ZN(new_n669));
  INV_X1    g0469(.A(new_n564), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n543), .B2(new_n394), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n560), .A2(new_n308), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n671), .A2(new_n672), .B1(new_n662), .B2(new_n663), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n530), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n665), .B1(new_n669), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT94), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n674), .B1(new_n530), .B2(new_n673), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n526), .B1(new_n505), .B2(new_n319), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n566), .A2(KEYINPUT26), .A3(new_n529), .A4(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n664), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT94), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n660), .B1(new_n678), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n655), .B1(new_n656), .B2(new_n684), .ZN(G369));
  INV_X1    g0485(.A(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n270), .A2(new_n226), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n587), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n602), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n589), .A2(new_n599), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n693), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n686), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n639), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n635), .A2(KEYINPUT93), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n698), .A2(new_n699), .B1(new_n617), .B2(new_n621), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n632), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n622), .A2(new_n692), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n692), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n692), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n695), .A2(new_n701), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n700), .A2(new_n707), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT96), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n708), .A2(KEYINPUT96), .A3(new_n709), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n706), .B1(new_n710), .B2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n222), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n520), .A2(new_n546), .A3(new_n580), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n714), .A2(new_n267), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n229), .B2(new_n714), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT28), .Z(new_n718));
  NAND3_X1  g0518(.A1(new_n567), .A2(new_n633), .A3(new_n657), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n692), .B1(new_n719), .B2(new_n682), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n684), .A2(new_n692), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(KEYINPUT29), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n579), .A2(new_n322), .A3(new_n543), .A4(new_n629), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n497), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n539), .A2(new_n634), .A3(KEYINPUT97), .A4(new_n542), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n590), .A2(new_n592), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n570), .B1(new_n729), .B2(new_n278), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(G179), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT97), .B1(new_n560), .B2(new_n634), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n727), .B1(new_n733), .B2(new_n497), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n539), .A2(new_n542), .A3(new_n634), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT97), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n594), .A3(new_n728), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n738), .A2(KEYINPUT30), .A3(new_n505), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n726), .B1(new_n734), .B2(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n692), .A2(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n642), .A2(new_n567), .A3(new_n707), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT98), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT30), .B1(new_n738), .B2(new_n505), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n728), .A2(G179), .A3(new_n730), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n746), .A2(new_n727), .A3(new_n497), .A4(new_n737), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n744), .B1(new_n748), .B2(new_n726), .ZN(new_n749));
  AOI211_X1 g0549(.A(KEYINPUT98), .B(new_n725), .C1(new_n745), .C2(new_n747), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n749), .A2(new_n750), .A3(new_n707), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n742), .B(new_n743), .C1(new_n751), .C2(KEYINPUT31), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G330), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n723), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n718), .B1(new_n754), .B2(G1), .ZN(G364));
  NOR2_X1   g0555(.A1(new_n264), .A2(G20), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G45), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(KEYINPUT99), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n267), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(KEYINPUT99), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n714), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n697), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n694), .A2(new_n696), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(G330), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n713), .A2(new_n328), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G355), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G116), .B2(new_n222), .ZN(new_n768));
  INV_X1    g0568(.A(G45), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n245), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n713), .A2(new_n285), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n769), .B2(new_n229), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n768), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  OR3_X1    g0574(.A1(KEYINPUT100), .A2(G13), .A3(G33), .ZN(new_n775));
  OAI21_X1  g0575(.A(KEYINPUT100), .B1(G13), .B2(G33), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n225), .B1(G20), .B2(new_n319), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n762), .B1(new_n774), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n226), .A2(G179), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n309), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G190), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G107), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n785), .A2(new_n394), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G87), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n787), .A2(new_n789), .A3(new_n285), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT101), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n226), .A2(new_n322), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(new_n394), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G190), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n793), .A2(new_n209), .B1(new_n795), .B2(new_n291), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT32), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n784), .A2(new_n794), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n407), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n394), .A2(G179), .A3(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n226), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n217), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n792), .A2(G190), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n806), .A2(new_n215), .B1(new_n797), .B2(new_n799), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n804), .A2(new_n442), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n803), .B(new_n807), .C1(G50), .C2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n791), .A2(new_n800), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n806), .A2(new_n811), .B1(new_n625), .B2(new_n802), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G326), .B2(new_n808), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n786), .A2(G283), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n788), .A2(G303), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n328), .B1(new_n795), .B2(new_n816), .ZN(new_n817));
  XOR2_X1   g0617(.A(KEYINPUT33), .B(G317), .Z(new_n818));
  NOR2_X1   g0618(.A1(new_n793), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n798), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n817), .B(new_n819), .C1(G329), .C2(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n810), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n783), .B1(new_n823), .B2(new_n780), .ZN(new_n824));
  INV_X1    g0624(.A(new_n779), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n764), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n765), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT102), .ZN(G396));
  NAND3_X1  g0628(.A1(new_n397), .A2(new_n398), .A3(new_n707), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n377), .A2(new_n707), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n393), .B2(new_n395), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n830), .B1(new_n399), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n396), .A2(new_n399), .A3(new_n707), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n722), .A2(new_n833), .B1(new_n684), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n762), .B1(new_n836), .B2(new_n753), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n753), .B2(new_n836), .ZN(new_n838));
  INV_X1    g0638(.A(new_n762), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n777), .A2(new_n780), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(new_n291), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n780), .ZN(new_n842));
  INV_X1    g0642(.A(new_n793), .ZN(new_n843));
  INV_X1    g0643(.A(new_n795), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n843), .A2(G150), .B1(new_n844), .B2(G159), .ZN(new_n845));
  INV_X1    g0645(.A(G143), .ZN(new_n846));
  INV_X1    g0646(.A(G137), .ZN(new_n847));
  INV_X1    g0647(.A(new_n808), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n845), .B1(new_n806), .B2(new_n846), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n786), .A2(G68), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n788), .A2(G50), .ZN(new_n853));
  INV_X1    g0653(.A(new_n802), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(G58), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n328), .B1(new_n820), .B2(G132), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n852), .A2(new_n853), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n849), .A2(new_n850), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n848), .A2(new_n572), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n803), .B(new_n860), .C1(G294), .C2(new_n805), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n786), .A2(G87), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n285), .B1(new_n843), .B2(G283), .ZN(new_n863));
  AOI22_X1  g0663(.A1(G116), .A2(new_n844), .B1(new_n820), .B2(G311), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(G107), .B2(new_n788), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n858), .A2(new_n859), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n841), .B1(new_n842), .B2(new_n867), .C1(new_n833), .C2(new_n778), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n838), .A2(new_n868), .ZN(G384));
  OR2_X1    g0669(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(G116), .A3(new_n227), .A4(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT36), .Z(new_n873));
  OAI211_X1 g0673(.A(new_n229), .B(G77), .C1(new_n215), .C2(new_n209), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n202), .A2(G68), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n267), .B(G13), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n412), .B1(new_n460), .B2(new_n209), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT16), .B1(new_n879), .B2(KEYINPUT105), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT105), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n430), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n462), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n454), .B1(new_n883), .B2(new_n405), .ZN(new_n884));
  INV_X1    g0684(.A(new_n690), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n883), .B2(new_n405), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n449), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n424), .A2(new_n431), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n404), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n454), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n885), .B1(new_n468), .B2(new_n405), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n891), .A2(new_n892), .A3(new_n449), .A4(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n888), .A2(KEYINPUT106), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n886), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n471), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT106), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n887), .A2(new_n898), .A3(KEYINPUT37), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n895), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n406), .B1(new_n430), .B2(new_n881), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n879), .A2(KEYINPUT105), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n431), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n404), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n906), .A2(new_n885), .B1(new_n432), .B2(new_n448), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n892), .B1(new_n907), .B2(new_n884), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n908), .A2(new_n898), .B1(new_n471), .B2(new_n896), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n902), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n740), .A2(KEYINPUT98), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n748), .A2(new_n744), .A3(new_n726), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n913), .A3(new_n741), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n743), .B(new_n914), .C1(new_n751), .C2(KEYINPUT31), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n365), .A2(new_n692), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT103), .ZN(new_n917));
  INV_X1    g0717(.A(new_n365), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n348), .B1(new_n340), .B2(G169), .ZN(new_n919));
  AOI211_X1 g0719(.A(KEYINPUT14), .B(new_n319), .C1(new_n335), .C2(new_n339), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n918), .B1(new_n921), .B2(new_n347), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n917), .B1(new_n922), .B2(new_n645), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n832), .A2(new_n399), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n916), .B(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n366), .A2(new_n926), .A3(new_n369), .ZN(new_n927));
  AND4_X1   g0727(.A1(new_n829), .A2(new_n923), .A3(new_n924), .A4(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n911), .A2(new_n915), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n893), .B1(new_n653), .B2(new_n647), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n891), .A2(new_n449), .A3(new_n893), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT37), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n894), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n930), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n878), .B1(new_n936), .B2(new_n910), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n833), .A2(new_n927), .A3(new_n923), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n749), .A2(new_n750), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT31), .B1(new_n939), .B2(new_n692), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n914), .A2(new_n743), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n878), .A2(new_n929), .B1(new_n937), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n474), .A3(new_n915), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(G330), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n944), .B1(new_n474), .B2(new_n915), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n829), .B1(new_n684), .B2(new_n835), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT104), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n923), .A2(new_n927), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n679), .A2(new_n681), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT94), .B1(new_n954), .B2(new_n665), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n677), .B(new_n664), .C1(new_n679), .C2(new_n681), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n719), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n830), .B1(new_n957), .B2(new_n834), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT104), .B1(new_n958), .B2(new_n951), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n953), .A2(new_n959), .A3(new_n911), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n651), .A2(new_n652), .A3(new_n690), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT39), .ZN(new_n962));
  INV_X1    g0762(.A(new_n930), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n456), .A2(KEYINPUT95), .A3(new_n469), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT95), .B1(new_n456), .B2(new_n469), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n647), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n893), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n963), .B1(new_n968), .B2(new_n934), .ZN(new_n969));
  AND4_X1   g0769(.A1(KEYINPUT38), .A2(new_n895), .A3(new_n899), .A4(new_n897), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n962), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n366), .A2(new_n692), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n902), .A2(new_n910), .A3(KEYINPUT39), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n960), .A2(new_n961), .A3(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n474), .B(new_n721), .C1(new_n722), .C2(KEYINPUT29), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n655), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n975), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n948), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n267), .B2(new_n756), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n948), .A2(new_n978), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n877), .B1(new_n980), .B2(new_n981), .ZN(G367));
  NAND2_X1  g0782(.A1(new_n692), .A2(new_n564), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n566), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n665), .B2(new_n983), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n527), .B(new_n530), .C1(new_n526), .C2(new_n707), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n530), .B1(new_n987), .B2(new_n640), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n707), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n668), .A2(new_n692), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n708), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(new_n992), .A3(KEYINPUT42), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT42), .B1(new_n991), .B2(new_n992), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n986), .B(new_n989), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT108), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT109), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n989), .B1(new_n994), .B2(new_n995), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n997), .A2(new_n998), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n998), .B1(new_n997), .B2(new_n1002), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n991), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n1004), .A2(new_n1005), .B1(new_n706), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1005), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n706), .A2(new_n1006), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n1009), .A3(new_n1003), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n714), .B(KEYINPUT41), .Z(new_n1011));
  INV_X1    g0811(.A(new_n695), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(new_n692), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n708), .B1(new_n1013), .B2(new_n705), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(new_n697), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT29), .B1(new_n957), .B2(new_n707), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n721), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1015), .B(new_n753), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(KEYINPUT110), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n991), .B1(new_n711), .B2(new_n710), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(KEYINPUT45), .B(new_n991), .C1(new_n711), .C2(new_n710), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n708), .A2(new_n709), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT96), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n708), .A2(KEYINPUT96), .A3(new_n709), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(new_n1028), .A3(new_n1006), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT44), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(KEYINPUT44), .A3(new_n1028), .A4(new_n1006), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1024), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n706), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT110), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n723), .A2(new_n1037), .A3(new_n753), .A4(new_n1015), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1024), .A2(new_n1033), .A3(new_n706), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1019), .A2(new_n1036), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1011), .B1(new_n1040), .B2(new_n754), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1007), .B(new_n1010), .C1(new_n1041), .C2(new_n761), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n240), .A2(new_n772), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n781), .B1(new_n222), .B2(new_n372), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n762), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n806), .A2(new_n572), .B1(new_n848), .B2(new_n816), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G107), .B2(new_n854), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n786), .A2(G97), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n285), .B1(new_n843), .B2(G294), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G283), .A2(new_n844), .B1(new_n820), .B2(G317), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n788), .A2(G116), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT46), .Z(new_n1053));
  NOR2_X1   g0853(.A1(new_n802), .A2(new_n209), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G143), .B2(new_n808), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n255), .B2(new_n806), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n786), .A2(G77), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n788), .A2(G58), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n328), .B1(new_n843), .B2(G159), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G50), .A2(new_n844), .B1(new_n820), .B2(G137), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n1051), .A2(new_n1053), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT47), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1045), .B1(new_n1063), .B2(new_n780), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n825), .B2(new_n985), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1042), .A2(new_n1065), .ZN(G387));
  NAND3_X1  g0866(.A1(new_n703), .A2(new_n704), .A3(new_n779), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n253), .A2(G50), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT50), .ZN(new_n1069));
  AOI211_X1 g0869(.A(G45), .B(new_n715), .C1(G68), .C2(G77), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n772), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n236), .B2(new_n769), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n766), .A2(new_n715), .B1(new_n211), .B2(new_n713), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1072), .B1(KEYINPUT111), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(KEYINPUT111), .B2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n762), .B1(new_n1075), .B2(new_n782), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n285), .B1(new_n795), .B2(new_n209), .C1(new_n253), .C2(new_n793), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n854), .A2(new_n557), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n806), .B2(new_n202), .C1(new_n407), .C2(new_n848), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1077), .B(new_n1079), .C1(G97), .C2(new_n786), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n788), .A2(G77), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n255), .B2(new_n798), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1082), .A2(KEYINPUT112), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(KEYINPUT112), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1080), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT113), .Z(new_n1086));
  INV_X1    g0886(.A(new_n788), .ZN(new_n1087));
  INV_X1    g0887(.A(G283), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1087), .A2(new_n625), .B1(new_n1088), .B2(new_n802), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n843), .A2(G311), .B1(new_n844), .B2(G303), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n805), .A2(G317), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(new_n811), .C2(new_n848), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT48), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1089), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n1093), .B2(new_n1092), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT49), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n285), .B1(new_n820), .B2(G326), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n786), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1098), .B1(new_n580), .B2(new_n1099), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1086), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1076), .B1(new_n1101), .B2(new_n780), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1015), .A2(new_n761), .B1(new_n1067), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n754), .A2(new_n1015), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1018), .A2(new_n714), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(G393));
  NAND2_X1  g0906(.A1(new_n1006), .A2(new_n779), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G311), .A2(new_n805), .B1(new_n808), .B2(G317), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT52), .Z(new_n1109));
  OAI21_X1  g0909(.A(new_n328), .B1(new_n795), .B2(new_n625), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n793), .A2(new_n572), .B1(new_n798), .B2(new_n811), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(G116), .C2(new_n854), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n788), .A2(G283), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1109), .A2(new_n787), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G150), .A2(new_n808), .B1(new_n805), .B2(G159), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT51), .Z(new_n1116));
  OAI21_X1  g0916(.A(new_n285), .B1(new_n798), .B2(new_n846), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n793), .A2(new_n202), .B1(new_n795), .B2(new_n253), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(G77), .C2(new_n854), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n788), .A2(G68), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1116), .A2(new_n862), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n842), .B1(new_n1114), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n781), .B1(new_n217), .B2(new_n222), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n251), .B2(new_n771), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n1122), .A2(new_n1124), .A3(new_n839), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1107), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n761), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n714), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n1127), .B2(new_n1018), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT114), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n1040), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1132), .B2(new_n1040), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1130), .B1(new_n1134), .B2(new_n1135), .ZN(G390));
  NAND2_X1  g0936(.A1(new_n914), .A2(new_n743), .ZN(new_n1137));
  OAI211_X1 g0937(.A(G330), .B(new_n928), .C1(new_n940), .C2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(KEYINPUT115), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n743), .A2(new_n742), .ZN(new_n1140));
  OAI211_X1 g0940(.A(G330), .B(new_n833), .C1(new_n940), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n951), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT115), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n915), .A2(new_n1143), .A3(G330), .A4(new_n928), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1139), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n949), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n752), .A2(new_n952), .A3(G330), .A4(new_n833), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n707), .B(new_n924), .C1(new_n660), .C2(new_n676), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n829), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n915), .A2(G330), .A3(new_n833), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n951), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1146), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n971), .A2(new_n973), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n972), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n958), .B2(new_n951), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n972), .B1(new_n936), .B2(new_n910), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1149), .A2(new_n952), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1159), .A2(new_n1162), .A3(new_n1147), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n949), .A2(new_n952), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1165), .A2(new_n1157), .B1(new_n971), .B2(new_n973), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1162), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1164), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n474), .A2(G330), .A3(new_n915), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n976), .A2(new_n655), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1155), .A2(new_n1163), .A3(new_n1168), .A4(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n714), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT116), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT116), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1172), .A2(new_n1175), .A3(new_n714), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1168), .A2(new_n1163), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT117), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT118), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1145), .A2(new_n949), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(new_n1170), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1155), .A2(KEYINPUT118), .A3(new_n1171), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1168), .A2(KEYINPUT117), .A3(new_n1163), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1179), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1174), .A2(new_n1176), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1177), .A2(new_n1128), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1156), .A2(new_n777), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n840), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n762), .B1(new_n401), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n789), .A2(new_n328), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT119), .Z(new_n1192));
  OAI22_X1  g0992(.A1(new_n795), .A2(new_n217), .B1(new_n798), .B2(new_n625), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G107), .B2(new_n843), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n808), .A2(G283), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G77), .A2(new_n854), .B1(new_n805), .B2(G116), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n852), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n786), .A2(G50), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n328), .B1(new_n843), .B2(G137), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(KEYINPUT54), .B(G143), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n844), .A2(new_n1201), .B1(new_n820), .B2(G125), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1198), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G159), .A2(new_n854), .B1(new_n805), .B2(G132), .ZN(new_n1204));
  INV_X1    g1004(.A(G128), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1204), .C1(new_n1205), .C2(new_n848), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n788), .A2(G150), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT53), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1192), .A2(new_n1197), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1190), .B1(new_n1209), .B2(new_n780), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1187), .B1(new_n1188), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1186), .A2(new_n1211), .ZN(G378));
  NAND3_X1  g1012(.A1(new_n311), .A2(new_n325), .A3(new_n316), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n273), .A2(new_n690), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1215), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n944), .B2(G330), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n902), .A2(new_n910), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n928), .B1(new_n940), .B2(new_n1137), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n878), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n937), .A2(new_n943), .ZN(new_n1227));
  AND4_X1   g1027(.A1(G330), .A2(new_n1226), .A3(new_n1227), .A4(new_n1222), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n975), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(G330), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1222), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n974), .A2(new_n961), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1226), .A2(new_n1227), .A3(new_n1222), .A4(G330), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1232), .A2(new_n960), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1229), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n761), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1222), .A2(new_n778), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G150), .A2(new_n854), .B1(new_n808), .B2(G125), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT121), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n843), .A2(G132), .B1(new_n844), .B2(G137), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n1205), .B2(new_n806), .C1(new_n1087), .C2(new_n1200), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(KEYINPUT59), .ZN(new_n1245));
  OR2_X1    g1045(.A1(KEYINPUT122), .A2(G124), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(KEYINPUT122), .A2(G124), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n820), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(G33), .A2(G41), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT120), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1248), .B(new_n1250), .C1(new_n1099), .C2(new_n407), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1244), .A2(new_n1245), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G41), .ZN(new_n1253));
  AOI211_X1 g1053(.A(G50), .B(new_n1250), .C1(new_n1253), .C2(new_n328), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n806), .A2(new_n211), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1054), .B(new_n1255), .C1(G116), .C2(new_n808), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n786), .A2(G58), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n793), .A2(new_n217), .B1(new_n795), .B2(new_n372), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1253), .B(new_n328), .C1(new_n798), .C2(new_n1088), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1256), .A2(new_n1081), .A3(new_n1257), .A4(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT58), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1254), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1262), .B2(new_n1261), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n780), .B1(new_n1252), .B2(new_n1264), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1265), .B(new_n762), .C1(G50), .C2(new_n1189), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1238), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1237), .A2(KEYINPUT123), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT123), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1128), .B1(new_n1229), .B2(new_n1235), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1270), .B1(new_n1271), .B2(new_n1267), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1172), .A2(new_n1171), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(KEYINPUT57), .A3(new_n1236), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1171), .A2(new_n1172), .B1(new_n1229), .B2(new_n1235), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1275), .B(new_n714), .C1(KEYINPUT57), .C2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(new_n1277), .ZN(G375));
  INV_X1    g1078(.A(new_n1011), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1181), .A2(new_n1170), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1183), .A2(new_n1182), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n762), .B1(G68), .B2(new_n1189), .ZN(new_n1282));
  OAI22_X1  g1082(.A1(new_n793), .A2(new_n1200), .B1(new_n798), .B2(new_n1205), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n328), .B(new_n1283), .C1(G150), .C2(new_n844), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1284), .B(new_n1257), .C1(new_n407), .C2(new_n1087), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(G50), .A2(new_n854), .B1(new_n808), .B2(G132), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n847), .B2(new_n806), .ZN(new_n1287));
  OAI221_X1 g1087(.A(new_n1078), .B1(new_n806), .B2(new_n1088), .C1(new_n625), .C2(new_n848), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n788), .A2(G97), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n285), .B1(new_n843), .B2(G116), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(G107), .A2(new_n844), .B1(new_n820), .B2(G303), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1057), .A2(new_n1289), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n1285), .A2(new_n1287), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1282), .B1(new_n1293), .B2(new_n780), .ZN(new_n1294));
  XOR2_X1   g1094(.A(new_n1294), .B(KEYINPUT124), .Z(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n952), .B2(new_n778), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1181), .B2(new_n1128), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1281), .A2(new_n1298), .ZN(G381));
  OR2_X1    g1099(.A1(G393), .A2(G396), .ZN(new_n1300));
  OR4_X1    g1100(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1300), .ZN(new_n1301));
  OR4_X1    g1101(.A1(G387), .A2(new_n1301), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1102(.A(G378), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n691), .A2(G213), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1303), .A2(new_n1277), .A3(new_n1273), .A4(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(G407), .A2(G213), .A3(new_n1306), .ZN(G409));
  NAND3_X1  g1107(.A1(G378), .A2(new_n1277), .A3(new_n1273), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1223), .A2(new_n1228), .A3(new_n975), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1232), .A2(new_n1234), .B1(new_n1233), .B2(new_n960), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT125), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT125), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1229), .A2(new_n1235), .A3(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(new_n761), .A3(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1274), .A2(new_n1279), .A3(new_n1236), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1314), .A2(new_n1268), .A3(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1316), .A2(new_n1186), .A3(new_n1211), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1308), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(G384), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1181), .A2(KEYINPUT60), .A3(new_n1170), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n714), .ZN(new_n1321));
  OAI21_X1  g1121(.A(KEYINPUT60), .B1(new_n1181), .B2(new_n1170), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1321), .B1(new_n1280), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1319), .B1(new_n1323), .B2(new_n1297), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1321), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1322), .A2(new_n1280), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1327), .A2(G384), .A3(new_n1298), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1324), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1318), .A2(new_n1304), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT62), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1318), .A2(new_n1304), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1305), .A2(G2897), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1329), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1324), .A2(new_n1328), .A3(new_n1334), .ZN(new_n1337));
  AND2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1333), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT61), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1305), .B1(new_n1308), .B2(new_n1317), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT62), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1330), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1332), .A2(new_n1339), .A3(new_n1340), .A4(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1132), .A2(new_n1040), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(KEYINPUT114), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1132), .A2(new_n1133), .A3(new_n1040), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1129), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(G387), .A2(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(G390), .A2(new_n1042), .A3(new_n1065), .ZN(new_n1350));
  XOR2_X1   g1150(.A(G393), .B(G396), .Z(new_n1351));
  AND3_X1   g1151(.A1(new_n1349), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1351), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1344), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1354), .B(new_n1340), .C1(new_n1341), .C2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1358), .ZN(new_n1359));
  AOI211_X1 g1159(.A(new_n1305), .B(new_n1329), .C1(new_n1308), .C2(new_n1317), .ZN(new_n1360));
  OAI21_X1  g1160(.A(KEYINPUT126), .B1(new_n1360), .B2(KEYINPUT63), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1360), .A2(KEYINPUT63), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT126), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT63), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1331), .A2(new_n1363), .A3(new_n1364), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1359), .A2(new_n1361), .A3(new_n1362), .A4(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1356), .A2(new_n1366), .ZN(G405));
  OR2_X1    g1167(.A1(new_n1330), .A2(KEYINPUT127), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1330), .A2(KEYINPUT127), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1308), .ZN(new_n1370));
  AOI21_X1  g1170(.A(G378), .B1(new_n1277), .B2(new_n1273), .ZN(new_n1371));
  OAI211_X1 g1171(.A(new_n1368), .B(new_n1369), .C1(new_n1370), .C2(new_n1371), .ZN(new_n1372));
  NOR2_X1   g1172(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1373), .A2(KEYINPUT127), .A3(new_n1330), .ZN(new_n1374));
  AND3_X1   g1174(.A1(new_n1372), .A2(new_n1354), .A3(new_n1374), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1354), .B1(new_n1372), .B2(new_n1374), .ZN(new_n1376));
  NOR2_X1   g1176(.A1(new_n1375), .A2(new_n1376), .ZN(G402));
endmodule


