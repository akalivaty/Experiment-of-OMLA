//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n586, new_n589, new_n590,
    new_n592, new_n593, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n454), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT64), .Z(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT65), .ZN(G160));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n466), .ZN(new_n476));
  INV_X1    g051(.A(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n466), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI22_X1  g054(.A1(new_n476), .A2(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n464), .A2(new_n466), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT66), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n480), .B1(new_n482), .B2(G124), .ZN(G162));
  OAI211_X1 g058(.A(G138), .B(new_n466), .C1(new_n462), .C2(new_n463), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n486), .A2(new_n466), .A3(G138), .ZN(new_n487));
  NOR3_X1   g062(.A1(new_n464), .A2(KEYINPUT67), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n490), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n489), .B1(new_n475), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n485), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G50), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n502), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n504), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n509), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  XNOR2_X1  g089(.A(new_n506), .B(KEYINPUT68), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n516));
  INV_X1    g091(.A(G51), .ZN(new_n517));
  INV_X1    g092(.A(new_n503), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n519), .A2(KEYINPUT69), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(KEYINPUT69), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n505), .A2(new_n506), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n522), .A2(G89), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n520), .A2(new_n521), .A3(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  AOI22_X1  g103(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n511), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n503), .A2(G52), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n507), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  NAND2_X1  g109(.A1(new_n515), .A2(G56), .ZN(new_n535));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n522), .A2(G81), .B1(G43), .B2(new_n503), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  NAND2_X1  g120(.A1(new_n522), .A2(G91), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n503), .A2(G53), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n548), .A2(KEYINPUT9), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(KEYINPUT9), .ZN(new_n550));
  OAI221_X1 g125(.A(new_n546), .B1(new_n511), .B2(new_n547), .C1(new_n549), .C2(new_n550), .ZN(G299));
  INV_X1    g126(.A(G171), .ZN(G301));
  NAND3_X1  g127(.A1(new_n522), .A2(KEYINPUT70), .A3(G87), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n554));
  INV_X1    g129(.A(G87), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n507), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n553), .A2(new_n556), .B1(G49), .B2(new_n503), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(G288));
  AOI22_X1  g134(.A1(new_n522), .A2(G86), .B1(G48), .B2(new_n503), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n506), .A2(G61), .ZN(new_n561));
  NAND2_X1  g136(.A1(G73), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(KEYINPUT71), .B1(new_n563), .B2(G651), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n565));
  AOI211_X1 g140(.A(new_n565), .B(new_n511), .C1(new_n561), .C2(new_n562), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n560), .B1(new_n564), .B2(new_n566), .ZN(G305));
  AOI22_X1  g142(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n511), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n522), .A2(G85), .B1(G47), .B2(new_n503), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(G290));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n572));
  INV_X1    g147(.A(G868), .ZN(new_n573));
  NOR2_X1   g148(.A1(G171), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n522), .A2(G92), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT10), .Z(new_n576));
  NAND2_X1  g151(.A1(new_n503), .A2(G54), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n511), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT73), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  AOI211_X1 g157(.A(new_n572), .B(new_n574), .C1(new_n573), .C2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n572), .B2(new_n574), .ZN(G284));
  AOI21_X1  g159(.A(new_n583), .B1(new_n572), .B2(new_n574), .ZN(G321));
  NAND2_X1  g160(.A1(G299), .A2(new_n573), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n586), .B1(G168), .B2(new_n573), .ZN(G297));
  OAI21_X1  g162(.A(new_n586), .B1(G168), .B2(new_n573), .ZN(G280));
  INV_X1    g163(.A(G860), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n582), .B1(G559), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT74), .ZN(G148));
  OR2_X1    g166(.A1(new_n582), .A2(G559), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G868), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(G868), .B2(new_n540), .ZN(G323));
  XOR2_X1   g169(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n595));
  XNOR2_X1  g170(.A(G323), .B(new_n595), .ZN(G282));
  NAND2_X1  g171(.A1(new_n475), .A2(new_n467), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT12), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT13), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(G2100), .ZN(new_n601));
  OAI21_X1  g176(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n602));
  INV_X1    g177(.A(G111), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G2105), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n465), .B2(G135), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n482), .B2(G123), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(G2096), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n600), .A2(G2100), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(G2096), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n601), .A2(new_n609), .A3(new_n610), .A4(new_n611), .ZN(G156));
  XOR2_X1   g187(.A(KEYINPUT15), .B(G2435), .Z(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT77), .B(G2438), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(G2427), .B(G2430), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT78), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(KEYINPUT76), .B(KEYINPUT14), .Z(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n617), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT79), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G1341), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G1348), .ZN(new_n624));
  XOR2_X1   g199(.A(G2451), .B(G2454), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n626), .B(new_n627), .Z(new_n628));
  OR2_X1    g203(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G14), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n624), .B2(new_n628), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(G401));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2072), .B(G2078), .Z(new_n636));
  XNOR2_X1  g211(.A(G2067), .B(G2678), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  NOR3_X1   g213(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT18), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n636), .A2(KEYINPUT80), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n636), .A2(KEYINPUT80), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(new_n642), .A3(new_n638), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n636), .B(KEYINPUT17), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n643), .B(new_n635), .C1(new_n644), .C2(new_n638), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(new_n638), .A3(new_n634), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n640), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2096), .B(G2100), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT81), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(G227));
  XNOR2_X1  g225(.A(G1971), .B(G1976), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1956), .B(G2474), .Z(new_n654));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  AND2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT20), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n654), .A2(new_n655), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  MUX2_X1   g236(.A(new_n661), .B(new_n660), .S(new_n653), .Z(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G229));
  INV_X1    g245(.A(G288), .ZN(new_n671));
  INV_X1    g246(.A(G16), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n672), .B2(G23), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT33), .B(G1976), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(G6), .A2(G16), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G305), .B2(new_n672), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT32), .B(G1981), .Z(new_n679));
  AOI22_X1  g254(.A1(new_n674), .A2(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n672), .A2(G22), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G166), .B2(new_n672), .ZN(new_n683));
  INV_X1    g258(.A(G1971), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND4_X1  g260(.A1(new_n676), .A2(new_n680), .A3(new_n681), .A4(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT83), .B(KEYINPUT34), .Z(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G25), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n482), .A2(G119), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n694));
  INV_X1    g269(.A(G107), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(G2105), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n465), .B2(G131), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n692), .B1(new_n699), .B2(new_n691), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n672), .A2(G24), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT82), .ZN(new_n704));
  INV_X1    g279(.A(G290), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n672), .ZN(new_n706));
  INV_X1    g281(.A(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n689), .A2(new_n690), .A3(new_n702), .A4(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(KEYINPUT84), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n709), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n672), .A2(G21), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G168), .B2(new_n672), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(G1966), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(G1966), .ZN(new_n716));
  NAND3_X1  g291(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT26), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n467), .A2(G105), .ZN(new_n719));
  INV_X1    g294(.A(G141), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n718), .B(new_n719), .C1(new_n720), .C2(new_n476), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n482), .B2(G129), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(new_n691), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n691), .B2(G32), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT27), .B(G1996), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT92), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n691), .A2(G27), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G164), .B2(new_n691), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2078), .ZN(new_n731));
  NOR4_X1   g306(.A1(new_n715), .A2(new_n716), .A3(new_n728), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(G160), .A2(G29), .ZN(new_n733));
  INV_X1    g308(.A(G34), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(KEYINPUT24), .ZN(new_n735));
  AOI21_X1  g310(.A(G29), .B1(new_n734), .B2(KEYINPUT24), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(KEYINPUT91), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(KEYINPUT91), .B2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(new_n466), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT25), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G139), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(new_n476), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(KEYINPUT90), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(KEYINPUT90), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n743), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G29), .ZN(new_n752));
  NOR2_X1   g327(.A1(G29), .A2(G33), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT89), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(new_n442), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n724), .A2(new_n727), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT31), .B(G11), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT30), .B(G28), .Z(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(G29), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n607), .B2(G29), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n672), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n672), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n757), .B(new_n761), .C1(new_n763), .C2(G1961), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n756), .B(new_n764), .C1(G1961), .C2(new_n763), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n739), .A2(new_n740), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n442), .B2(new_n755), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n732), .A2(new_n741), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT93), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(G29), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G2090), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT95), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n672), .A2(G20), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT23), .Z(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G299), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT96), .ZN(new_n779));
  INV_X1    g354(.A(G1956), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n775), .B(new_n781), .C1(G2090), .C2(new_n773), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n672), .A2(G4), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n581), .B2(new_n672), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1348), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n672), .A2(G19), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT85), .Z(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n540), .B2(new_n672), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1341), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n691), .A2(G26), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT28), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n482), .A2(G128), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(G116), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G2105), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT86), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n465), .A2(G140), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n793), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT87), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n793), .A2(KEYINPUT87), .A3(new_n797), .A4(new_n798), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n792), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2067), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n790), .A2(KEYINPUT88), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(KEYINPUT88), .B1(new_n790), .B2(new_n805), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n782), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n712), .A2(new_n769), .A3(new_n808), .ZN(G150));
  INV_X1    g384(.A(G150), .ZN(G311));
  NAND2_X1  g385(.A1(new_n581), .A2(G559), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT98), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n522), .A2(G93), .B1(G55), .B2(new_n503), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n515), .A2(G67), .ZN(new_n815));
  NAND2_X1  g390(.A1(G80), .A2(G543), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n511), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT97), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g394(.A(KEYINPUT97), .B(new_n511), .C1(new_n815), .C2(new_n816), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(new_n540), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n813), .B(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(new_n589), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n821), .A2(new_n589), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(G145));
  XOR2_X1   g404(.A(G160), .B(G162), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT99), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n608), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n751), .A2(KEYINPUT102), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n835));
  NAND2_X1  g410(.A1(G126), .A2(G2105), .ZN(new_n836));
  OR2_X1    g411(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n837));
  NAND2_X1  g412(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n466), .A2(G114), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n835), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n494), .A2(new_n497), .A3(KEYINPUT100), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n846), .A3(new_n493), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT67), .B1(new_n464), .B2(new_n487), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n475), .A2(new_n489), .A3(new_n491), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n848), .A2(new_n849), .B1(KEYINPUT4), .B2(new_n484), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n843), .A2(new_n844), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT101), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n834), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n466), .B2(G118), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n856), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n855), .A2(new_n466), .A3(G118), .ZN(new_n858));
  INV_X1    g433(.A(G142), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n857), .A2(new_n858), .B1(new_n476), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(new_n482), .B2(G130), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n598), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n854), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n722), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n803), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n722), .B1(new_n801), .B2(new_n802), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n699), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OR3_X1    g442(.A1(new_n865), .A2(new_n699), .A3(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n863), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n863), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n867), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n833), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n869), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n874), .B2(new_n832), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(G395));
  OAI21_X1  g453(.A(new_n573), .B1(new_n819), .B2(new_n820), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n581), .B(G299), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT41), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n822), .B(new_n592), .ZN(new_n882));
  MUX2_X1   g457(.A(new_n881), .B(new_n880), .S(new_n882), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(G290), .B(G166), .ZN(new_n885));
  XNOR2_X1  g460(.A(G288), .B(G305), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n884), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n879), .B1(new_n889), .B2(new_n573), .ZN(G295));
  OAI21_X1  g465(.A(new_n879), .B1(new_n889), .B2(new_n573), .ZN(G331));
  NAND2_X1  g466(.A1(G286), .A2(G301), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n520), .A2(G171), .A3(new_n521), .A4(new_n526), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n822), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n895), .A2(new_n880), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n822), .B2(new_n894), .ZN(new_n898));
  OR3_X1    g473(.A1(new_n822), .A2(new_n894), .A3(new_n897), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n822), .A2(new_n894), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n895), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n881), .A2(new_n902), .A3(KEYINPUT105), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT105), .B1(new_n881), .B2(new_n902), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n888), .B(new_n900), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n881), .A2(new_n902), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n881), .A2(new_n902), .A3(KEYINPUT105), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n888), .B1(new_n912), .B2(new_n900), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n899), .A2(new_n895), .A3(new_n898), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n915), .A2(new_n881), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n896), .A2(new_n901), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n887), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n918), .A2(new_n905), .A3(new_n919), .A4(new_n906), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(new_n905), .A3(new_n906), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n924), .B2(KEYINPUT43), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n905), .A2(new_n906), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n912), .A2(new_n900), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n887), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n928), .A3(new_n919), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n925), .A2(new_n929), .A3(KEYINPUT107), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT107), .B1(new_n925), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(G397));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n933), .B1(new_n853), .B2(G1384), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n468), .A2(G40), .A3(new_n472), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n803), .B(G2067), .ZN(new_n937));
  INV_X1    g512(.A(G1996), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n722), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n936), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n936), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n698), .B(new_n701), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n936), .A2(new_n938), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n943), .B(new_n944), .ZN(new_n945));
  OAI221_X1 g520(.A(new_n940), .B1(new_n941), .B2(new_n942), .C1(new_n945), .C2(new_n864), .ZN(new_n946));
  NOR2_X1   g521(.A1(G290), .A2(G1986), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT108), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n707), .B2(new_n705), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n936), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n951));
  INV_X1    g526(.A(G8), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(G168), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n493), .A2(new_n843), .A3(new_n844), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT45), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT114), .B1(new_n956), .B2(new_n935), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n494), .A2(new_n497), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n955), .B1(new_n850), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n960), .B2(new_n933), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n498), .A2(KEYINPUT115), .A3(KEYINPUT45), .A4(new_n955), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n955), .B1(new_n850), .B2(new_n851), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n933), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n966));
  INV_X1    g541(.A(new_n935), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n957), .A2(new_n963), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1966), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n954), .A2(new_n972), .A3(new_n955), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n974));
  AND4_X1   g549(.A1(new_n740), .A2(new_n973), .A3(new_n974), .A4(new_n967), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n953), .B1(new_n977), .B2(G8), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n966), .B1(new_n965), .B2(new_n967), .ZN(new_n979));
  AOI211_X1 g554(.A(KEYINPUT114), .B(new_n935), .C1(new_n964), .C2(new_n933), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(G1966), .B1(new_n981), .B2(new_n963), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT120), .B1(new_n982), .B2(new_n975), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT120), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n971), .A2(new_n984), .A3(new_n976), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(G168), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n951), .A2(new_n952), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n978), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(G168), .A2(new_n952), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n984), .B1(new_n971), .B2(new_n976), .ZN(new_n990));
  AOI211_X1 g565(.A(KEYINPUT120), .B(new_n975), .C1(new_n969), .C2(new_n970), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT62), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT62), .ZN(new_n995));
  INV_X1    g570(.A(new_n987), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n990), .A2(new_n991), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n996), .B1(new_n997), .B2(G168), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n995), .B(new_n992), .C1(new_n998), .C2(new_n978), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT124), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G303), .A2(G8), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT55), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n845), .B2(new_n493), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(new_n972), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n967), .B1(new_n960), .B2(KEYINPUT50), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1004), .A2(new_n1005), .A3(G2090), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n847), .A2(new_n852), .A3(KEYINPUT45), .A4(new_n955), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n935), .B1(new_n960), .B2(new_n933), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1006), .B1(new_n684), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1002), .B1(new_n1010), .B2(new_n952), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n952), .B1(new_n1003), .B2(new_n967), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G305), .A2(G1981), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT111), .B(G1981), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n560), .B(new_n1015), .C1(new_n564), .C2(new_n566), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT112), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT49), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1013), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g594(.A(KEYINPUT112), .B(KEYINPUT49), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1012), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(KEYINPUT113), .A3(new_n1026), .A4(new_n1013), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1021), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n973), .A2(new_n974), .A3(new_n967), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT110), .B1(new_n1029), .B2(G2090), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1009), .A2(new_n684), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n935), .B1(new_n1003), .B2(new_n972), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n1033));
  INV_X1    g608(.A(G2090), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n974), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1030), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1002), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(G8), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n671), .B2(G1976), .ZN(new_n1040));
  INV_X1    g615(.A(G1976), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1013), .B1(new_n1041), .B2(G288), .ZN(new_n1042));
  MUX2_X1   g617(.A(new_n1040), .B(new_n1039), .S(new_n1042), .Z(new_n1043));
  AND4_X1   g618(.A1(new_n1011), .A2(new_n1028), .A3(new_n1038), .A4(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n1009), .B2(G2078), .ZN(new_n1046));
  INV_X1    g621(.A(G1961), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1029), .A2(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n957), .A2(new_n963), .A3(new_n968), .A4(new_n443), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT53), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1054), .A2(G171), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1044), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n994), .A2(new_n999), .A3(new_n1000), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1036), .A2(G8), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1037), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1059), .B2(new_n1058), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n952), .B(G286), .C1(new_n971), .C2(new_n976), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1062), .A2(KEYINPUT63), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1028), .A2(new_n1043), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1061), .A2(new_n1063), .A3(new_n1038), .A4(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1028), .A2(new_n1011), .A3(new_n1038), .A4(new_n1043), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1062), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT117), .B(KEYINPUT63), .Z(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1067), .A2(new_n1068), .A3(new_n1066), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1065), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n1074));
  XNOR2_X1  g649(.A(G299), .B(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n780), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1007), .A2(new_n1008), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1348), .B1(new_n1032), .B2(new_n974), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1003), .A2(new_n967), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(G2067), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(new_n582), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1075), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1079), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  NAND2_X1  g662(.A1(new_n1081), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1009), .B2(G1996), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n540), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(KEYINPUT59), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n540), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1079), .A2(KEYINPUT61), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1075), .A2(new_n1076), .A3(new_n1097), .A4(new_n1078), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1348), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1029), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(KEYINPUT60), .C1(G2067), .C2(new_n1081), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(new_n1104), .A3(new_n581), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1083), .A2(KEYINPUT60), .A3(new_n582), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1086), .B1(new_n1099), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n934), .A2(new_n967), .A3(new_n1007), .A4(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1029), .A2(KEYINPUT123), .A3(new_n1047), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT123), .B1(new_n1029), .B2(new_n1047), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1046), .B(new_n1111), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1109), .B1(new_n1114), .B2(G171), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1054), .B2(G171), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1108), .A2(new_n1044), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n992), .B1(new_n998), .B2(new_n978), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1114), .A2(G171), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1109), .B1(new_n1055), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1028), .A2(new_n1041), .A3(new_n671), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1016), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1038), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1123), .A2(new_n1013), .B1(new_n1064), .B2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1057), .A2(new_n1073), .A3(new_n1121), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1044), .A2(new_n1055), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n1118), .B2(KEYINPUT62), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1000), .B1(new_n1128), .B2(new_n999), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n950), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n936), .B1(new_n937), .B2(new_n864), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n945), .A2(KEYINPUT46), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n945), .A2(KEYINPUT46), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT47), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n946), .A2(KEYINPUT125), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n946), .A2(KEYINPUT125), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n948), .A2(new_n941), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1138), .B(KEYINPUT48), .Z(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n940), .B1(new_n945), .B2(new_n864), .ZN(new_n1141));
  INV_X1    g716(.A(new_n701), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1141), .A2(new_n1142), .A3(new_n698), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n803), .A2(G2067), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n936), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1135), .A2(new_n1140), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1130), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT126), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1130), .A2(new_n1149), .A3(new_n1146), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n1153));
  INV_X1    g727(.A(G319), .ZN(new_n1154));
  NOR2_X1   g728(.A1(new_n1154), .A2(G227), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n669), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g730(.A(new_n1156), .B1(new_n629), .B2(new_n631), .ZN(new_n1157));
  NAND2_X1  g731(.A1(new_n876), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g732(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g733(.A(new_n1153), .B1(new_n921), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g734(.A(KEYINPUT127), .B(new_n1158), .C1(new_n914), .C2(new_n920), .ZN(new_n1161));
  NOR2_X1   g735(.A1(new_n1160), .A2(new_n1161), .ZN(G308));
  AOI21_X1  g736(.A(new_n919), .B1(new_n926), .B2(new_n928), .ZN(new_n1163));
  INV_X1    g737(.A(new_n920), .ZN(new_n1164));
  OAI21_X1  g738(.A(new_n1159), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n1165), .A2(KEYINPUT127), .ZN(new_n1166));
  NAND3_X1  g740(.A1(new_n921), .A2(new_n1153), .A3(new_n1159), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1167), .ZN(G225));
endmodule


