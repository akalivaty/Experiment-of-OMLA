//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G101), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT77), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n189), .A2(new_n192), .A3(new_n198), .A4(new_n193), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n199), .A2(KEYINPUT4), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(KEYINPUT77), .A3(G101), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT64), .B1(new_n203), .B2(G146), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n205), .A3(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n205), .B2(G143), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n203), .A2(KEYINPUT65), .A3(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n207), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n210), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n194), .A2(new_n223), .A3(G101), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n202), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G137), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT11), .A3(G134), .ZN(new_n227));
  INV_X1    g041(.A(G134), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G137), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n231));
  INV_X1    g045(.A(G131), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n228), .B2(G137), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n230), .A2(new_n231), .A3(new_n232), .A4(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n234), .A2(new_n227), .A3(new_n232), .A4(new_n229), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n229), .A3(new_n227), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n235), .A2(new_n237), .B1(G131), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n188), .A2(G107), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n191), .A2(G104), .ZN(new_n241));
  OAI21_X1  g055(.A(G101), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n199), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT1), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n214), .A2(new_n218), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n244), .B1(new_n206), .B2(KEYINPUT1), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(new_n218), .B2(new_n214), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n243), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n214), .A2(new_n218), .A3(new_n245), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n203), .A2(G146), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  OAI21_X1  g068(.A(G128), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n204), .A2(new_n206), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT10), .A3(new_n243), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n225), .A2(new_n239), .A3(new_n251), .A4(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G110), .B(G140), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G227), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n261), .B(new_n263), .ZN(new_n264));
  XOR2_X1   g078(.A(KEYINPUT75), .B(KEYINPUT76), .Z(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n238), .A2(G131), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n199), .A2(new_n242), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n219), .A2(new_n255), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(new_n274), .B2(new_n252), .ZN(new_n275));
  INV_X1    g089(.A(new_n250), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n259), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n194), .A2(KEYINPUT77), .A3(G101), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT77), .B1(new_n194), .B2(G101), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n199), .A2(KEYINPUT4), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n207), .B1(new_n214), .B2(new_n218), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n224), .B1(new_n282), .B2(new_n210), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n272), .B1(new_n277), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n268), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n260), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n273), .A2(new_n252), .A3(new_n257), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n235), .A2(new_n237), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n249), .A2(new_n288), .B1(new_n289), .B2(new_n269), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT80), .B1(new_n290), .B2(KEYINPUT12), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n273), .A2(new_n252), .A3(new_n257), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n272), .B1(new_n275), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT80), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT12), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(KEYINPUT12), .B(new_n272), .C1(new_n275), .C2(new_n292), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT79), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT79), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n290), .A2(new_n300), .A3(KEYINPUT12), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n287), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(G469), .B(new_n286), .C1(new_n303), .C2(new_n266), .ZN(new_n304));
  INV_X1    g118(.A(G469), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n267), .B1(new_n297), .B2(new_n302), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n266), .B1(new_n285), .B2(new_n260), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(G469), .A2(G902), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n304), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT9), .B(G234), .ZN(new_n312));
  OAI21_X1  g126(.A(G221), .B1(new_n312), .B2(G902), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT89), .ZN(new_n315));
  XNOR2_X1  g129(.A(G113), .B(G122), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(new_n188), .ZN(new_n317));
  INV_X1    g131(.A(G237), .ZN(new_n318));
  AND4_X1   g132(.A1(G143), .A2(new_n318), .A3(new_n262), .A4(G214), .ZN(new_n319));
  NOR2_X1   g133(.A1(G237), .A2(G953), .ZN(new_n320));
  AOI21_X1  g134(.A(G143), .B1(new_n320), .B2(G214), .ZN(new_n321));
  OAI21_X1  g135(.A(G131), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT17), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n318), .A2(new_n262), .A3(G214), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n203), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n320), .A2(G143), .A3(G214), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n232), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n322), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G125), .B(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n331), .A2(KEYINPUT16), .A3(G140), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n205), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n332), .B1(new_n329), .B2(KEYINPUT16), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G146), .ZN(new_n337));
  OAI211_X1 g151(.A(KEYINPUT17), .B(G131), .C1(new_n319), .C2(new_n321), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n328), .A2(new_n335), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT18), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(new_n232), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n319), .B2(new_n321), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT86), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n329), .B(new_n205), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT86), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n345), .B(new_n341), .C1(new_n319), .C2(new_n321), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n325), .B(new_n326), .C1(new_n340), .C2(new_n232), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n343), .A2(new_n344), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n317), .B1(new_n339), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n339), .A2(new_n317), .A3(new_n348), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT88), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT88), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n339), .A2(new_n352), .A3(new_n348), .A4(new_n317), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n349), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G475), .B1(new_n354), .B2(G902), .ZN(new_n355));
  XOR2_X1   g169(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n353), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n322), .A2(new_n327), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT87), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n329), .A2(new_n359), .A3(KEYINPUT19), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT19), .B1(new_n329), .B2(new_n359), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n205), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n336), .A2(KEYINPUT73), .A3(G146), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT73), .B1(new_n336), .B2(G146), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n358), .B(new_n362), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n317), .B1(new_n365), .B2(new_n348), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n357), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(G475), .A2(G902), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n356), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n366), .B1(new_n351), .B2(new_n353), .ZN(new_n371));
  INV_X1    g185(.A(new_n369), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n371), .A2(KEYINPUT20), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n315), .B(new_n355), .C1(new_n370), .C2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT20), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n368), .A2(new_n376), .A3(new_n369), .ZN(new_n377));
  INV_X1    g191(.A(new_n356), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n378), .B1(new_n371), .B2(new_n372), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n315), .B1(new_n380), .B2(new_n355), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G478), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(KEYINPUT15), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT90), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n203), .A2(G128), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n203), .A2(G128), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT13), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n385), .B(new_n386), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n244), .A2(G143), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n244), .A2(G143), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n390), .B1(KEYINPUT13), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT90), .B1(new_n386), .B2(new_n388), .ZN(new_n393));
  OAI211_X1 g207(.A(G134), .B(new_n389), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n390), .A2(new_n387), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n228), .ZN(new_n396));
  XNOR2_X1  g210(.A(G116), .B(G122), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(new_n191), .ZN(new_n398));
  INV_X1    g212(.A(G122), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G116), .ZN(new_n400));
  INV_X1    g214(.A(G116), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G122), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G107), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n394), .B(new_n396), .C1(new_n398), .C2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G134), .B1(new_n390), .B2(new_n387), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n396), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n397), .A2(new_n191), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n401), .A2(KEYINPUT14), .A3(G122), .ZN(new_n409));
  OAI211_X1 g223(.A(G107), .B(new_n409), .C1(new_n403), .C2(KEYINPUT14), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G217), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n312), .A2(new_n412), .A3(G953), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n405), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n413), .B1(new_n405), .B2(new_n411), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n384), .B1(new_n417), .B2(G902), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n405), .A2(new_n411), .ZN(new_n419));
  INV_X1    g233(.A(new_n413), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n414), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n422), .B(new_n306), .C1(KEYINPUT15), .C2(new_n383), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n418), .A2(new_n423), .A3(KEYINPUT91), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT91), .B1(new_n418), .B2(new_n423), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(G234), .A2(G237), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(G952), .A3(new_n262), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT92), .Z(new_n429));
  AND3_X1   g243(.A1(new_n427), .A2(G902), .A3(G953), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(G898), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n426), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n314), .A2(new_n382), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G214), .B1(G237), .B2(G902), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT6), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n438));
  INV_X1    g252(.A(G119), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(G116), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G116), .B(G119), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n440), .B(G113), .C1(new_n442), .C2(new_n438), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT2), .ZN(new_n444));
  INV_X1    g258(.A(G113), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT67), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(KEYINPUT2), .B2(G113), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(KEYINPUT2), .A2(G113), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n441), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n443), .A2(new_n243), .A3(new_n451), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n449), .A2(new_n450), .A3(new_n441), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n441), .B1(new_n449), .B2(new_n450), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n224), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n452), .B1(new_n281), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G110), .B(G122), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n437), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n454), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n194), .A2(G101), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n460), .A2(new_n451), .B1(new_n461), .B2(new_n223), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n453), .A2(new_n273), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n462), .A2(new_n202), .B1(new_n443), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT82), .B1(new_n464), .B2(new_n457), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n457), .B(new_n452), .C1(new_n281), .C2(new_n455), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT82), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n459), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n456), .A2(new_n437), .A3(new_n458), .ZN(new_n470));
  INV_X1    g284(.A(G224), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(G953), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n258), .A2(new_n331), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT83), .ZN(new_n475));
  OAI21_X1  g289(.A(G125), .B1(new_n282), .B2(new_n210), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n474), .B2(new_n476), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n479), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n472), .A3(new_n477), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n469), .A2(new_n470), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n466), .B(new_n467), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n457), .B(KEYINPUT8), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n441), .A2(KEYINPUT5), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n440), .A2(new_n487), .A3(G113), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n463), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n243), .B1(new_n443), .B2(new_n451), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n474), .A2(new_n476), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT7), .A3(new_n473), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n473), .A2(KEYINPUT7), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n474), .A2(new_n476), .A3(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(G902), .B1(new_n485), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT84), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n484), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n498), .B1(new_n484), .B2(new_n497), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n484), .A2(new_n497), .A3(new_n501), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n436), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n187), .B1(new_n435), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n318), .A2(new_n262), .A3(G210), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT27), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT26), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT27), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n506), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT26), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n198), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n512), .A3(G101), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n514), .A2(KEYINPUT69), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT69), .B1(new_n514), .B2(new_n515), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n226), .A2(G134), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n232), .B1(new_n519), .B2(new_n229), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n252), .B2(new_n257), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n289), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n453), .A2(new_n454), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(new_n523), .C1(new_n239), .C2(new_n221), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT28), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT70), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(KEYINPUT70), .A3(new_n525), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT68), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n272), .A2(new_n222), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n521), .A2(new_n289), .A3(KEYINPUT68), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n531), .A2(new_n523), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n523), .ZN(new_n535));
  INV_X1    g349(.A(new_n522), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n221), .B1(new_n289), .B2(new_n269), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n525), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n518), .B1(new_n529), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n521), .A2(new_n289), .A3(KEYINPUT68), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n537), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n543), .B2(new_n531), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n522), .B(new_n541), .C1(new_n239), .C2(new_n221), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n535), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n515), .ZN(new_n548));
  AOI21_X1  g362(.A(G101), .B1(new_n508), .B2(new_n512), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n534), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT31), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n532), .A2(new_n533), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT68), .B1(new_n521), .B2(new_n289), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT30), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n523), .B1(new_n556), .B2(new_n545), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT31), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n557), .A2(new_n558), .A3(new_n551), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n540), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(G472), .A2(G902), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(KEYINPUT32), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n558), .B1(new_n557), .B2(new_n551), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n546), .B1(KEYINPUT30), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n552), .B(KEYINPUT31), .C1(new_n566), .C2(new_n523), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n524), .A2(KEYINPUT70), .A3(new_n525), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(new_n526), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n534), .A2(new_n538), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT28), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n564), .A2(new_n567), .B1(new_n572), .B2(new_n518), .ZN(new_n573));
  INV_X1    g387(.A(new_n561), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n563), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n523), .B1(new_n543), .B2(new_n531), .ZN(new_n576));
  INV_X1    g390(.A(new_n534), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT28), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n569), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n539), .A2(new_n568), .A3(new_n526), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n518), .A2(KEYINPUT29), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n579), .A2(KEYINPUT29), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n550), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n547), .A2(new_n534), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(KEYINPUT29), .ZN(new_n585));
  AOI21_X1  g399(.A(G902), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G472), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n562), .B(new_n575), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n412), .B1(G234), .B2(new_n306), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n335), .A2(new_n337), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT24), .B(G110), .Z(new_n592));
  XNOR2_X1  g406(.A(G119), .B(G128), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT71), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n595), .B(KEYINPUT23), .C1(new_n244), .C2(G119), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n439), .A2(G128), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n596), .B(new_n597), .C1(new_n595), .C2(KEYINPUT23), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n599), .A3(G110), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n591), .A2(new_n594), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n363), .A2(new_n364), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n329), .A2(new_n205), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT72), .B(G110), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n598), .B2(new_n599), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n592), .A2(new_n593), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n601), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT22), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G137), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n601), .B(new_n611), .C1(new_n602), .C2(new_n607), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n306), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT25), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT74), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n613), .A2(new_n306), .A3(new_n617), .A4(new_n614), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n590), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n613), .A2(new_n614), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n589), .A2(G902), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n588), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n355), .B1(new_n370), .B2(new_n373), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT89), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n434), .A2(new_n374), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n436), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n484), .A2(new_n497), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT84), .ZN(new_n631));
  INV_X1    g445(.A(new_n501), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n484), .A2(new_n497), .A3(new_n498), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n484), .A2(new_n497), .A3(new_n501), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n629), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n628), .A2(new_n636), .A3(KEYINPUT93), .A4(new_n314), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n505), .A2(new_n625), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G101), .ZN(G3));
  NOR2_X1   g453(.A1(new_n417), .A2(G902), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(G478), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT33), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n415), .B2(new_n416), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT94), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT94), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n422), .A2(new_n645), .A3(new_n642), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n421), .A2(KEYINPUT33), .A3(new_n414), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT95), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT95), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n421), .A2(new_n649), .A3(KEYINPUT33), .A4(new_n414), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n644), .A2(new_n646), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n383), .A2(G902), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n641), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n627), .B2(new_n374), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n501), .B1(new_n484), .B2(new_n497), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n629), .B1(new_n657), .B2(new_n635), .ZN(new_n658));
  INV_X1    g472(.A(new_n433), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n573), .B2(G902), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n560), .A2(new_n561), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n624), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n311), .A2(new_n313), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT34), .B(G104), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G6));
  NAND3_X1  g484(.A1(new_n368), .A2(new_n369), .A3(new_n356), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n379), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n672), .A2(new_n355), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n426), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n660), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT35), .B(G107), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT96), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n676), .B(new_n678), .ZN(G9));
  INV_X1    g493(.A(KEYINPUT97), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n619), .A2(new_n620), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n589), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n612), .A2(KEYINPUT36), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n608), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n623), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n680), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n682), .A2(new_n680), .A3(new_n685), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n664), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n505), .A2(new_n637), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  NOR2_X1   g505(.A1(new_n687), .A2(new_n686), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n436), .B1(new_n503), .B2(new_n656), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n666), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(G900), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n430), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n429), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n674), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n588), .A2(new_n692), .A3(new_n694), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G128), .ZN(G30));
  XOR2_X1   g514(.A(new_n697), .B(KEYINPUT100), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT39), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n666), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT40), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n516), .A2(new_n517), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n565), .A2(new_n535), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n705), .B1(new_n534), .B2(new_n706), .ZN(new_n707));
  OAI22_X1  g521(.A1(new_n707), .A2(KEYINPUT99), .B1(new_n557), .B2(new_n551), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n707), .A2(KEYINPUT99), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n306), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G472), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n711), .A2(new_n575), .A3(new_n562), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n426), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n627), .B2(new_n374), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n682), .A2(new_n685), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n629), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n704), .A2(new_n713), .A3(new_n715), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n634), .A2(new_n635), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n203), .ZN(G45));
  AOI211_X1 g537(.A(new_n653), .B(new_n697), .C1(new_n627), .C2(new_n374), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n588), .A2(new_n724), .A3(new_n692), .A4(new_n694), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G146), .ZN(G48));
  NAND2_X1  g540(.A1(new_n297), .A2(new_n302), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n308), .B1(new_n727), .B2(new_n268), .ZN(new_n728));
  OAI21_X1  g542(.A(G469), .B1(new_n728), .B2(G902), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n313), .A3(new_n309), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT101), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(KEYINPUT101), .A3(new_n313), .A4(new_n309), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n625), .A2(new_n661), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NAND3_X1  g551(.A1(new_n625), .A2(new_n675), .A3(new_n734), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  NAND3_X1  g553(.A1(new_n732), .A2(new_n658), .A3(new_n733), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT102), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n732), .A2(KEYINPUT102), .A3(new_n658), .A4(new_n733), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n588), .A2(new_n628), .A3(new_n692), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G119), .ZN(G21));
  NAND2_X1  g561(.A1(new_n564), .A2(new_n567), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n579), .A2(new_n518), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n561), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n662), .A2(new_n751), .A3(new_n624), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT103), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n715), .A2(new_n658), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n732), .A2(new_n659), .A3(new_n733), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  AOI21_X1  g572(.A(new_n574), .B1(new_n748), .B2(new_n749), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n560), .A2(new_n306), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n759), .B1(new_n760), .B2(G472), .ZN(new_n761));
  INV_X1    g575(.A(new_n697), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n654), .A3(new_n716), .A4(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n742), .B2(new_n743), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n331), .ZN(G27));
  NAND2_X1  g579(.A1(new_n588), .A2(new_n624), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n503), .A2(new_n629), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n634), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT104), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n634), .A2(new_n769), .A3(KEYINPUT104), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n772), .A2(new_n314), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(KEYINPUT42), .A3(new_n724), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n314), .A3(new_n773), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n654), .A2(new_n762), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n776), .A2(new_n766), .A3(new_n777), .ZN(new_n778));
  OAI22_X1  g592(.A1(new_n768), .A2(new_n775), .B1(new_n778), .B2(KEYINPUT42), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G131), .ZN(G33));
  INV_X1    g594(.A(new_n698), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n776), .A2(new_n766), .A3(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT106), .B(G134), .Z(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G36));
  AOI22_X1  g598(.A1(new_n662), .A2(new_n663), .B1(new_n682), .B2(new_n685), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT108), .ZN(new_n786));
  INV_X1    g600(.A(new_n653), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n382), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT43), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT44), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n786), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT107), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n286), .B1(new_n303), .B2(new_n266), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT45), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n305), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n798), .B2(new_n797), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n310), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n796), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n800), .A2(KEYINPUT107), .A3(KEYINPUT46), .A4(new_n310), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n309), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n313), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n772), .A2(new_n773), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n807), .A2(new_n702), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n795), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G137), .ZN(G39));
  NAND2_X1  g625(.A1(new_n807), .A2(KEYINPUT47), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n806), .A2(new_n813), .A3(new_n313), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n808), .A2(new_n588), .A3(new_n624), .A4(new_n777), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  INV_X1    g631(.A(new_n429), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n790), .A2(new_n818), .A3(new_n753), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n744), .ZN(new_n820));
  INV_X1    g634(.A(G952), .ZN(new_n821));
  INV_X1    g635(.A(new_n734), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n808), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n624), .A2(new_n823), .A3(new_n818), .A4(new_n712), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n821), .B(G953), .C1(new_n824), .C2(new_n654), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n790), .A2(new_n818), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(new_n823), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT48), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n766), .B(KEYINPUT105), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n827), .B2(new_n829), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n820), .B(new_n825), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n812), .A2(new_n814), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n729), .A2(new_n309), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n833), .B1(new_n313), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n819), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n808), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n837), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n824), .A2(new_n382), .A3(new_n653), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n826), .A2(new_n716), .A3(new_n761), .A4(new_n823), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT50), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n822), .B2(new_n436), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n734), .A2(KEYINPUT112), .A3(new_n629), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n721), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n847), .B1(new_n839), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n851), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(KEYINPUT50), .A3(new_n819), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n846), .A2(KEYINPUT51), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n832), .B1(new_n842), .B2(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n839), .A2(new_n847), .A3(new_n851), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT50), .B1(new_n853), .B2(new_n819), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT113), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n852), .A2(new_n861), .A3(new_n854), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n860), .A2(new_n846), .A3(KEYINPUT114), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n836), .A2(new_n840), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n845), .B1(new_n855), .B2(KEYINPUT113), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT114), .B1(new_n866), .B2(new_n862), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n857), .B1(new_n868), .B2(KEYINPUT51), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT42), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n776), .A2(new_n870), .A3(new_n777), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n774), .A2(new_n625), .A3(new_n724), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n829), .A2(new_n871), .B1(new_n872), .B2(new_n870), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT110), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n436), .B(new_n659), .C1(new_n502), .C2(new_n503), .ZN(new_n875));
  INV_X1    g689(.A(new_n418), .ZN(new_n876));
  INV_X1    g690(.A(new_n423), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n375), .A2(new_n381), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n874), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n636), .A2(KEYINPUT110), .A3(new_n879), .A4(new_n659), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n667), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n746), .A2(new_n757), .A3(new_n883), .A4(new_n738), .ZN(new_n884));
  INV_X1    g698(.A(new_n875), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n654), .A2(KEYINPUT109), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n654), .A2(KEYINPUT109), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n667), .A2(new_n885), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n638), .A2(new_n689), .A3(new_n735), .A4(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n876), .A2(new_n877), .A3(new_n697), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n588), .A2(new_n673), .A3(new_n692), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n763), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n774), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n774), .A2(new_n625), .A3(new_n698), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR4_X1   g709(.A1(new_n873), .A2(new_n884), .A3(new_n889), .A4(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n763), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n744), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n725), .A2(new_n699), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n716), .A2(new_n697), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n715), .A2(new_n314), .A3(new_n658), .A4(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n712), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n898), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT52), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n725), .A2(new_n699), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n764), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(KEYINPUT52), .A3(new_n903), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n896), .A2(KEYINPUT53), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n884), .A2(new_n889), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n872), .A2(new_n870), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n829), .A2(new_n871), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n895), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n910), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT53), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n911), .A2(new_n918), .ZN(new_n919));
  AND4_X1   g733(.A1(new_n738), .A2(new_n746), .A3(new_n757), .A4(new_n883), .ZN(new_n920));
  AND4_X1   g734(.A1(new_n638), .A2(new_n689), .A3(new_n735), .A4(new_n888), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n776), .B1(new_n763), .B2(new_n891), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n922), .A2(new_n782), .A3(new_n917), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n920), .A2(new_n921), .A3(new_n779), .A4(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT52), .B1(new_n908), .B2(new_n903), .ZN(new_n925));
  NOR4_X1   g739(.A1(new_n764), .A2(new_n907), .A3(new_n905), .A4(new_n902), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT111), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT53), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n873), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT111), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n910), .A2(new_n930), .A3(new_n931), .A4(new_n912), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT54), .B1(new_n916), .B2(new_n917), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n919), .A2(KEYINPUT54), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI22_X1  g750(.A1(new_n869), .A2(new_n936), .B1(G952), .B2(G953), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n835), .A2(KEYINPUT49), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n624), .A2(new_n436), .A3(new_n313), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n835), .A2(KEYINPUT49), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n788), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(new_n721), .A3(new_n712), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n937), .A2(new_n943), .ZN(G75));
  NAND2_X1  g758(.A1(new_n821), .A2(G953), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT116), .Z(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT56), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n933), .A2(new_n918), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(G902), .ZN(new_n950));
  INV_X1    g764(.A(G210), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n469), .A2(new_n470), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(new_n483), .Z(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT55), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n955), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n948), .B(new_n957), .C1(new_n950), .C2(new_n951), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n947), .B1(new_n956), .B2(new_n958), .ZN(G51));
  INV_X1    g773(.A(new_n728), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT117), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n933), .A2(new_n961), .A3(new_n934), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(new_n933), .B2(new_n934), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT54), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n933), .B2(new_n918), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n310), .B(KEYINPUT57), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n960), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n950), .A2(new_n800), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n947), .B1(new_n968), .B2(new_n969), .ZN(G54));
  AND4_X1   g784(.A1(KEYINPUT58), .A2(new_n949), .A3(G475), .A4(G902), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n971), .A2(new_n371), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n371), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n947), .B1(new_n972), .B2(new_n973), .ZN(G60));
  INV_X1    g788(.A(new_n651), .ZN(new_n975));
  NAND2_X1  g789(.A1(G478), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT59), .Z(new_n977));
  OR2_X1    g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n946), .B1(new_n966), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT118), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT53), .B1(new_n896), .B2(new_n910), .ZN(new_n981));
  AND4_X1   g795(.A1(KEYINPUT53), .A2(new_n910), .A3(new_n912), .A4(new_n915), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT54), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n933), .A2(new_n934), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n977), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n980), .B1(new_n985), .B2(new_n651), .ZN(new_n986));
  OAI211_X1 g800(.A(KEYINPUT118), .B(new_n975), .C1(new_n935), .C2(new_n977), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n979), .A2(new_n988), .ZN(G63));
  XNOR2_X1  g803(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n412), .A2(new_n306), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n949), .A2(new_n684), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n622), .ZN(new_n994));
  AOI22_X1  g808(.A1(new_n928), .A2(new_n932), .B1(new_n917), .B2(new_n916), .ZN(new_n995));
  INV_X1    g809(.A(new_n992), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n993), .A2(new_n997), .A3(new_n946), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n998), .A2(KEYINPUT119), .A3(KEYINPUT61), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT61), .B1(new_n998), .B2(KEYINPUT119), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(G66));
  NOR3_X1   g815(.A1(new_n431), .A2(new_n471), .A3(new_n262), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n912), .B2(new_n262), .ZN(new_n1003));
  INV_X1    g817(.A(G898), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n953), .B1(new_n1004), .B2(G953), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1003), .B(new_n1005), .Z(G69));
  NAND2_X1  g820(.A1(new_n886), .A2(new_n887), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n702), .B1(new_n1007), .B2(new_n880), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n776), .A2(new_n766), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(KEYINPUT123), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT123), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1008), .A2(new_n1012), .A3(new_n1009), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n810), .A2(new_n816), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n908), .A2(KEYINPUT122), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT122), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n764), .B2(new_n907), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n722), .ZN(new_n1020));
  AOI21_X1  g834(.A(KEYINPUT62), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n1019), .A2(KEYINPUT62), .A3(new_n1020), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1015), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n262), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n360), .A2(new_n361), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1025), .B(KEYINPUT121), .Z(new_n1026));
  XNOR2_X1  g840(.A(new_n566), .B(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1027), .B1(G900), .B2(G953), .ZN(new_n1029));
  AND2_X1   g843(.A1(new_n810), .A2(new_n816), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n807), .A2(new_n702), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n768), .A2(new_n754), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n782), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n1033), .A2(new_n779), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1030), .A2(new_n1034), .A3(new_n1019), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1029), .B1(new_n1035), .B2(G953), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1038), .B1(new_n1036), .B2(KEYINPUT124), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1037), .B(new_n1039), .Z(G72));
  OAI211_X1 g854(.A(new_n1015), .B(new_n912), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1041));
  NAND2_X1  g855(.A1(G472), .A2(G902), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT63), .Z(new_n1043));
  AND3_X1   g857(.A1(new_n1041), .A2(KEYINPUT125), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g858(.A(KEYINPUT125), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1045));
  INV_X1    g859(.A(new_n584), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1046), .A2(new_n583), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  NOR3_X1   g862(.A1(new_n1044), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  NAND4_X1  g863(.A1(new_n1030), .A2(new_n1034), .A3(new_n912), .A4(new_n1019), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1050), .A2(new_n1043), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1046), .A2(new_n583), .ZN(new_n1052));
  XNOR2_X1  g866(.A(new_n1052), .B(KEYINPUT126), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g868(.A(new_n919), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1048), .A2(new_n1043), .A3(new_n1052), .ZN(new_n1056));
  OAI211_X1 g870(.A(new_n1054), .B(new_n946), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g871(.A(KEYINPUT127), .B1(new_n1049), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1045), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n1041), .A2(KEYINPUT125), .A3(new_n1043), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1059), .A2(new_n1060), .A3(new_n1047), .ZN(new_n1061));
  INV_X1    g875(.A(KEYINPUT127), .ZN(new_n1062));
  OR2_X1    g876(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1063));
  AOI21_X1  g877(.A(new_n947), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1064));
  NAND4_X1  g878(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1058), .A2(new_n1065), .ZN(G57));
endmodule


