

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U552 ( .A1(G8), .A2(n686), .ZN(n730) );
  OR2_X1 U553 ( .A1(KEYINPUT33), .A2(n713), .ZN(n721) );
  OR2_X1 U554 ( .A1(n730), .A2(n729), .ZN(n518) );
  AND2_X1 U555 ( .A1(n731), .A2(n518), .ZN(n519) );
  INV_X1 U556 ( .A(KEYINPUT30), .ZN(n625) );
  INV_X1 U557 ( .A(KEYINPUT96), .ZN(n628) );
  NOR2_X1 U558 ( .A1(n730), .A2(G1966), .ZN(n623) );
  AND2_X1 U559 ( .A1(n732), .A2(n519), .ZN(n733) );
  NOR2_X1 U560 ( .A1(G651), .A2(G543), .ZN(n779) );
  NOR2_X1 U561 ( .A1(G651), .A2(n543), .ZN(n785) );
  INV_X1 U562 ( .A(G651), .ZN(n525) );
  NOR2_X1 U563 ( .A1(G543), .A2(n525), .ZN(n521) );
  XNOR2_X1 U564 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n520) );
  XNOR2_X1 U565 ( .A(n521), .B(n520), .ZN(n783) );
  NAND2_X1 U566 ( .A1(G60), .A2(n783), .ZN(n523) );
  XOR2_X1 U567 ( .A(KEYINPUT0), .B(G543), .Z(n543) );
  NAND2_X1 U568 ( .A1(G47), .A2(n785), .ZN(n522) );
  NAND2_X1 U569 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U570 ( .A(KEYINPUT66), .B(n524), .Z(n529) );
  NAND2_X1 U571 ( .A1(G85), .A2(n779), .ZN(n527) );
  NOR2_X1 U572 ( .A1(n543), .A2(n525), .ZN(n780) );
  NAND2_X1 U573 ( .A1(G72), .A2(n780), .ZN(n526) );
  AND2_X1 U574 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U575 ( .A1(n529), .A2(n528), .ZN(G290) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  XOR2_X2 U577 ( .A(KEYINPUT17), .B(n530), .Z(n869) );
  NAND2_X1 U578 ( .A1(G138), .A2(n869), .ZN(n532) );
  INV_X1 U579 ( .A(G2105), .ZN(n533) );
  AND2_X1 U580 ( .A1(n533), .A2(G2104), .ZN(n871) );
  NAND2_X1 U581 ( .A1(G102), .A2(n871), .ZN(n531) );
  NAND2_X1 U582 ( .A1(n532), .A2(n531), .ZN(n537) );
  AND2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n864) );
  NAND2_X1 U584 ( .A1(G114), .A2(n864), .ZN(n535) );
  NOR2_X1 U585 ( .A1(G2104), .A2(n533), .ZN(n865) );
  NAND2_X1 U586 ( .A1(G126), .A2(n865), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U588 ( .A1(n537), .A2(n536), .ZN(G164) );
  NAND2_X1 U589 ( .A1(G651), .A2(G74), .ZN(n538) );
  XOR2_X1 U590 ( .A(KEYINPUT75), .B(n538), .Z(n540) );
  NAND2_X1 U591 ( .A1(n785), .A2(G49), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U593 ( .A(KEYINPUT76), .B(n541), .ZN(n542) );
  NOR2_X1 U594 ( .A1(n783), .A2(n542), .ZN(n545) );
  NAND2_X1 U595 ( .A1(n543), .A2(G87), .ZN(n544) );
  NAND2_X1 U596 ( .A1(n545), .A2(n544), .ZN(G288) );
  NAND2_X1 U597 ( .A1(G88), .A2(n779), .ZN(n547) );
  NAND2_X1 U598 ( .A1(G75), .A2(n780), .ZN(n546) );
  NAND2_X1 U599 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U600 ( .A1(G62), .A2(n783), .ZN(n549) );
  NAND2_X1 U601 ( .A1(G50), .A2(n785), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U603 ( .A1(n551), .A2(n550), .ZN(G166) );
  INV_X1 U604 ( .A(G166), .ZN(G303) );
  NAND2_X1 U605 ( .A1(n780), .A2(G76), .ZN(n552) );
  XNOR2_X1 U606 ( .A(KEYINPUT72), .B(n552), .ZN(n555) );
  NAND2_X1 U607 ( .A1(n779), .A2(G89), .ZN(n553) );
  XNOR2_X1 U608 ( .A(KEYINPUT4), .B(n553), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U610 ( .A(n556), .B(KEYINPUT5), .ZN(n561) );
  NAND2_X1 U611 ( .A1(G63), .A2(n783), .ZN(n558) );
  NAND2_X1 U612 ( .A1(G51), .A2(n785), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U614 ( .A(KEYINPUT6), .B(n559), .Z(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U616 ( .A(n562), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U617 ( .A1(n785), .A2(G52), .ZN(n564) );
  NAND2_X1 U618 ( .A1(n783), .A2(G64), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n564), .A2(n563), .ZN(n569) );
  NAND2_X1 U620 ( .A1(G90), .A2(n779), .ZN(n566) );
  NAND2_X1 U621 ( .A1(G77), .A2(n780), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U623 ( .A(KEYINPUT9), .B(n567), .Z(n568) );
  NOR2_X1 U624 ( .A1(n569), .A2(n568), .ZN(G171) );
  INV_X1 U625 ( .A(G171), .ZN(G301) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G86), .A2(n779), .ZN(n571) );
  NAND2_X1 U628 ( .A1(G61), .A2(n783), .ZN(n570) );
  NAND2_X1 U629 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U630 ( .A(KEYINPUT77), .B(n572), .Z(n575) );
  NAND2_X1 U631 ( .A1(n780), .A2(G73), .ZN(n573) );
  XOR2_X1 U632 ( .A(KEYINPUT2), .B(n573), .Z(n574) );
  NOR2_X1 U633 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U634 ( .A(n576), .B(KEYINPUT78), .ZN(n578) );
  NAND2_X1 U635 ( .A1(G48), .A2(n785), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n578), .A2(n577), .ZN(G305) );
  XNOR2_X1 U637 ( .A(G1986), .B(G290), .ZN(n938) );
  NOR2_X1 U638 ( .A1(G164), .A2(G1384), .ZN(n621) );
  NAND2_X1 U639 ( .A1(G101), .A2(n871), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT23), .B(n579), .Z(n752) );
  AND2_X1 U641 ( .A1(G40), .A2(n752), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n864), .A2(G113), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n869), .A2(G137), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U645 ( .A(KEYINPUT64), .B(n582), .Z(n584) );
  NAND2_X1 U646 ( .A1(n865), .A2(G125), .ZN(n583) );
  AND2_X1 U647 ( .A1(n584), .A2(n583), .ZN(n753) );
  AND2_X1 U648 ( .A1(n585), .A2(n753), .ZN(n622) );
  INV_X1 U649 ( .A(n622), .ZN(n586) );
  NOR2_X1 U650 ( .A1(n621), .A2(n586), .ZN(n747) );
  NAND2_X1 U651 ( .A1(n938), .A2(n747), .ZN(n736) );
  NAND2_X1 U652 ( .A1(n869), .A2(G141), .ZN(n594) );
  NAND2_X1 U653 ( .A1(G117), .A2(n864), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G129), .A2(n865), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U656 ( .A(KEYINPUT88), .B(n589), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n871), .A2(G105), .ZN(n590) );
  XOR2_X1 U658 ( .A(KEYINPUT38), .B(n590), .Z(n591) );
  NOR2_X1 U659 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U661 ( .A(KEYINPUT89), .B(n595), .Z(n881) );
  NAND2_X1 U662 ( .A1(G1996), .A2(n881), .ZN(n604) );
  NAND2_X1 U663 ( .A1(G107), .A2(n864), .ZN(n597) );
  NAND2_X1 U664 ( .A1(G119), .A2(n865), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U666 ( .A1(G131), .A2(n869), .ZN(n598) );
  XNOR2_X1 U667 ( .A(KEYINPUT87), .B(n598), .ZN(n599) );
  NOR2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n871), .A2(G95), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n602), .A2(n601), .ZN(n877) );
  NAND2_X1 U671 ( .A1(G1991), .A2(n877), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U673 ( .A(KEYINPUT90), .B(n605), .Z(n973) );
  XNOR2_X1 U674 ( .A(n747), .B(KEYINPUT91), .ZN(n606) );
  NOR2_X1 U675 ( .A1(n973), .A2(n606), .ZN(n739) );
  INV_X1 U676 ( .A(n739), .ZN(n619) );
  NAND2_X1 U677 ( .A1(G140), .A2(n869), .ZN(n608) );
  NAND2_X1 U678 ( .A1(G104), .A2(n871), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U680 ( .A(KEYINPUT34), .B(n609), .ZN(n617) );
  XNOR2_X1 U681 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n615) );
  NAND2_X1 U682 ( .A1(n864), .A2(G116), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n610), .B(KEYINPUT84), .ZN(n612) );
  NAND2_X1 U684 ( .A1(G128), .A2(n865), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n613), .B(KEYINPUT35), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n615), .B(n614), .ZN(n616) );
  NOR2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(KEYINPUT36), .ZN(n889) );
  XNOR2_X1 U690 ( .A(G2067), .B(KEYINPUT37), .ZN(n744) );
  NOR2_X1 U691 ( .A1(n889), .A2(n744), .ZN(n967) );
  NAND2_X1 U692 ( .A1(n747), .A2(n967), .ZN(n742) );
  NAND2_X1 U693 ( .A1(n619), .A2(n742), .ZN(n734) );
  NOR2_X1 U694 ( .A1(G1976), .A2(G288), .ZN(n714) );
  NOR2_X1 U695 ( .A1(G1971), .A2(G303), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n714), .A2(n620), .ZN(n941) );
  XOR2_X1 U697 ( .A(n941), .B(KEYINPUT97), .Z(n708) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n686) );
  XNOR2_X1 U699 ( .A(n623), .B(KEYINPUT93), .ZN(n702) );
  NAND2_X1 U700 ( .A1(G8), .A2(n702), .ZN(n624) );
  NOR2_X1 U701 ( .A1(G2084), .A2(n686), .ZN(n699) );
  NOR2_X1 U702 ( .A1(n624), .A2(n699), .ZN(n626) );
  XNOR2_X1 U703 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X1 U704 ( .A1(G168), .A2(n627), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n629), .B(n628), .ZN(n633) );
  XOR2_X1 U706 ( .A(G2078), .B(KEYINPUT25), .Z(n923) );
  NOR2_X1 U707 ( .A1(n923), .A2(n686), .ZN(n631) );
  INV_X1 U708 ( .A(n686), .ZN(n657) );
  NOR2_X1 U709 ( .A1(n657), .A2(G1961), .ZN(n630) );
  NOR2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n635), .A2(G301), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U713 ( .A(KEYINPUT31), .B(n634), .ZN(n700) );
  OR2_X1 U714 ( .A1(n635), .A2(G301), .ZN(n685) );
  NAND2_X1 U715 ( .A1(G65), .A2(n783), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G53), .A2(n785), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G91), .A2(n779), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G78), .A2(n780), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U721 ( .A1(n641), .A2(n640), .ZN(n947) );
  NAND2_X1 U722 ( .A1(G2072), .A2(n657), .ZN(n644) );
  XOR2_X1 U723 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n642) );
  XNOR2_X1 U724 ( .A(KEYINPUT27), .B(n642), .ZN(n643) );
  XNOR2_X1 U725 ( .A(n644), .B(n643), .ZN(n646) );
  AND2_X1 U726 ( .A1(n686), .A2(G1956), .ZN(n645) );
  NOR2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n648) );
  NOR2_X1 U728 ( .A1(n947), .A2(n648), .ZN(n647) );
  XOR2_X1 U729 ( .A(n647), .B(KEYINPUT28), .Z(n682) );
  NAND2_X1 U730 ( .A1(n947), .A2(n648), .ZN(n680) );
  NAND2_X1 U731 ( .A1(n785), .A2(G54), .ZN(n655) );
  NAND2_X1 U732 ( .A1(G92), .A2(n779), .ZN(n650) );
  NAND2_X1 U733 ( .A1(G79), .A2(n780), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U735 ( .A1(G66), .A2(n783), .ZN(n651) );
  XNOR2_X1 U736 ( .A(KEYINPUT71), .B(n651), .ZN(n652) );
  NOR2_X1 U737 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U738 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U739 ( .A(KEYINPUT15), .B(n656), .Z(n950) );
  NAND2_X1 U740 ( .A1(G1348), .A2(n686), .ZN(n659) );
  NAND2_X1 U741 ( .A1(n657), .A2(G2067), .ZN(n658) );
  NAND2_X1 U742 ( .A1(n659), .A2(n658), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n950), .A2(n674), .ZN(n678) );
  XOR2_X1 U744 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n661) );
  NAND2_X1 U745 ( .A1(G56), .A2(n783), .ZN(n660) );
  XNOR2_X1 U746 ( .A(n661), .B(n660), .ZN(n667) );
  NAND2_X1 U747 ( .A1(n779), .A2(G81), .ZN(n662) );
  XNOR2_X1 U748 ( .A(n662), .B(KEYINPUT12), .ZN(n664) );
  NAND2_X1 U749 ( .A1(G68), .A2(n780), .ZN(n663) );
  NAND2_X1 U750 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U751 ( .A(KEYINPUT13), .B(n665), .Z(n666) );
  NOR2_X1 U752 ( .A1(n667), .A2(n666), .ZN(n669) );
  NAND2_X1 U753 ( .A1(n785), .A2(G43), .ZN(n668) );
  NAND2_X1 U754 ( .A1(n669), .A2(n668), .ZN(n937) );
  INV_X1 U755 ( .A(G1996), .ZN(n916) );
  NOR2_X1 U756 ( .A1(n686), .A2(n916), .ZN(n670) );
  XOR2_X1 U757 ( .A(n670), .B(KEYINPUT26), .Z(n672) );
  NAND2_X1 U758 ( .A1(n686), .A2(G1341), .ZN(n671) );
  NAND2_X1 U759 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U760 ( .A1(n937), .A2(n673), .ZN(n676) );
  NOR2_X1 U761 ( .A1(n950), .A2(n674), .ZN(n675) );
  OR2_X1 U762 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U763 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U765 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U766 ( .A(KEYINPUT29), .B(n683), .Z(n684) );
  NAND2_X1 U767 ( .A1(n685), .A2(n684), .ZN(n701) );
  INV_X1 U768 ( .A(G8), .ZN(n691) );
  NOR2_X1 U769 ( .A1(G1971), .A2(n730), .ZN(n688) );
  NOR2_X1 U770 ( .A1(G2090), .A2(n686), .ZN(n687) );
  NOR2_X1 U771 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U772 ( .A1(n689), .A2(G303), .ZN(n690) );
  OR2_X1 U773 ( .A1(n691), .A2(n690), .ZN(n693) );
  AND2_X1 U774 ( .A1(n701), .A2(n693), .ZN(n692) );
  NAND2_X1 U775 ( .A1(n700), .A2(n692), .ZN(n697) );
  INV_X1 U776 ( .A(n693), .ZN(n695) );
  AND2_X1 U777 ( .A1(G286), .A2(G8), .ZN(n694) );
  OR2_X1 U778 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U779 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U780 ( .A(n698), .B(KEYINPUT32), .ZN(n707) );
  NAND2_X1 U781 ( .A1(G8), .A2(n699), .ZN(n705) );
  NAND2_X1 U782 ( .A1(n701), .A2(n700), .ZN(n703) );
  AND2_X1 U783 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U784 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U785 ( .A1(n707), .A2(n706), .ZN(n724) );
  NAND2_X1 U786 ( .A1(n708), .A2(n724), .ZN(n709) );
  XNOR2_X1 U787 ( .A(n709), .B(KEYINPUT98), .ZN(n712) );
  NAND2_X1 U788 ( .A1(G1976), .A2(G288), .ZN(n940) );
  INV_X1 U789 ( .A(n940), .ZN(n710) );
  NOR2_X1 U790 ( .A1(n730), .A2(n710), .ZN(n711) );
  AND2_X1 U791 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U792 ( .A1(KEYINPUT33), .A2(n714), .ZN(n715) );
  XOR2_X1 U793 ( .A(KEYINPUT99), .B(n715), .Z(n716) );
  NOR2_X1 U794 ( .A1(n730), .A2(n716), .ZN(n717) );
  XNOR2_X1 U795 ( .A(n717), .B(KEYINPUT100), .ZN(n719) );
  XOR2_X1 U796 ( .A(G1981), .B(G305), .Z(n953) );
  INV_X1 U797 ( .A(n953), .ZN(n718) );
  NOR2_X1 U798 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U799 ( .A1(n721), .A2(n720), .ZN(n732) );
  NOR2_X1 U800 ( .A1(G2090), .A2(G303), .ZN(n722) );
  NAND2_X1 U801 ( .A1(G8), .A2(n722), .ZN(n723) );
  NAND2_X1 U802 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U803 ( .A(KEYINPUT101), .B(n725), .Z(n726) );
  NAND2_X1 U804 ( .A1(n726), .A2(n730), .ZN(n731) );
  NOR2_X1 U805 ( .A1(G1981), .A2(G305), .ZN(n727) );
  XOR2_X1 U806 ( .A(n727), .B(KEYINPUT24), .Z(n728) );
  XNOR2_X1 U807 ( .A(KEYINPUT92), .B(n728), .ZN(n729) );
  NOR2_X1 U808 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U809 ( .A1(n736), .A2(n735), .ZN(n750) );
  NOR2_X1 U810 ( .A1(G1996), .A2(n881), .ZN(n985) );
  NOR2_X1 U811 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U812 ( .A1(G1991), .A2(n877), .ZN(n969) );
  NOR2_X1 U813 ( .A1(n737), .A2(n969), .ZN(n738) );
  NOR2_X1 U814 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U815 ( .A1(n985), .A2(n740), .ZN(n741) );
  XNOR2_X1 U816 ( .A(n741), .B(KEYINPUT39), .ZN(n743) );
  NAND2_X1 U817 ( .A1(n743), .A2(n742), .ZN(n745) );
  NAND2_X1 U818 ( .A1(n889), .A2(n744), .ZN(n965) );
  NAND2_X1 U819 ( .A1(n745), .A2(n965), .ZN(n746) );
  NAND2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U821 ( .A(KEYINPUT102), .B(n748), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U823 ( .A(n751), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U824 ( .A1(n753), .A2(n752), .ZN(G160) );
  AND2_X1 U825 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U826 ( .A1(G7), .A2(G661), .ZN(n754) );
  XNOR2_X1 U827 ( .A(n754), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U828 ( .A(G223), .B(KEYINPUT68), .Z(n819) );
  NAND2_X1 U829 ( .A1(n819), .A2(G567), .ZN(n755) );
  XNOR2_X1 U830 ( .A(n755), .B(KEYINPUT11), .ZN(n756) );
  XNOR2_X1 U831 ( .A(KEYINPUT69), .B(n756), .ZN(G234) );
  INV_X1 U832 ( .A(G860), .ZN(n762) );
  OR2_X1 U833 ( .A1(n937), .A2(n762), .ZN(G153) );
  NAND2_X1 U834 ( .A1(G868), .A2(G301), .ZN(n758) );
  INV_X1 U835 ( .A(G868), .ZN(n759) );
  NAND2_X1 U836 ( .A1(n950), .A2(n759), .ZN(n757) );
  NAND2_X1 U837 ( .A1(n758), .A2(n757), .ZN(G284) );
  INV_X1 U838 ( .A(n947), .ZN(G299) );
  NOR2_X1 U839 ( .A1(G286), .A2(n759), .ZN(n761) );
  NOR2_X1 U840 ( .A1(G868), .A2(G299), .ZN(n760) );
  NOR2_X1 U841 ( .A1(n761), .A2(n760), .ZN(G297) );
  NAND2_X1 U842 ( .A1(n762), .A2(G559), .ZN(n763) );
  INV_X1 U843 ( .A(n950), .ZN(n893) );
  NAND2_X1 U844 ( .A1(n763), .A2(n893), .ZN(n764) );
  XNOR2_X1 U845 ( .A(n764), .B(KEYINPUT73), .ZN(n765) );
  XOR2_X1 U846 ( .A(KEYINPUT16), .B(n765), .Z(G148) );
  NOR2_X1 U847 ( .A1(G868), .A2(n937), .ZN(n768) );
  NAND2_X1 U848 ( .A1(G868), .A2(n893), .ZN(n766) );
  NOR2_X1 U849 ( .A1(G559), .A2(n766), .ZN(n767) );
  NOR2_X1 U850 ( .A1(n768), .A2(n767), .ZN(G282) );
  NAND2_X1 U851 ( .A1(G123), .A2(n865), .ZN(n769) );
  XNOR2_X1 U852 ( .A(n769), .B(KEYINPUT18), .ZN(n771) );
  NAND2_X1 U853 ( .A1(n864), .A2(G111), .ZN(n770) );
  NAND2_X1 U854 ( .A1(n771), .A2(n770), .ZN(n775) );
  NAND2_X1 U855 ( .A1(G135), .A2(n869), .ZN(n773) );
  NAND2_X1 U856 ( .A1(G99), .A2(n871), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U858 ( .A1(n775), .A2(n774), .ZN(n970) );
  XNOR2_X1 U859 ( .A(G2096), .B(n970), .ZN(n777) );
  INV_X1 U860 ( .A(G2100), .ZN(n776) );
  NAND2_X1 U861 ( .A1(n777), .A2(n776), .ZN(G156) );
  NAND2_X1 U862 ( .A1(n893), .A2(G559), .ZN(n799) );
  XNOR2_X1 U863 ( .A(n937), .B(n799), .ZN(n778) );
  NOR2_X1 U864 ( .A1(n778), .A2(G860), .ZN(n790) );
  NAND2_X1 U865 ( .A1(G93), .A2(n779), .ZN(n782) );
  NAND2_X1 U866 ( .A1(G80), .A2(n780), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n789) );
  NAND2_X1 U868 ( .A1(n783), .A2(G67), .ZN(n784) );
  XNOR2_X1 U869 ( .A(n784), .B(KEYINPUT74), .ZN(n787) );
  NAND2_X1 U870 ( .A1(G55), .A2(n785), .ZN(n786) );
  NAND2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U872 ( .A1(n789), .A2(n788), .ZN(n802) );
  XNOR2_X1 U873 ( .A(n790), .B(n802), .ZN(G145) );
  XNOR2_X1 U874 ( .A(KEYINPUT19), .B(KEYINPUT79), .ZN(n792) );
  XNOR2_X1 U875 ( .A(G290), .B(KEYINPUT80), .ZN(n791) );
  XNOR2_X1 U876 ( .A(n792), .B(n791), .ZN(n793) );
  XNOR2_X1 U877 ( .A(n947), .B(n793), .ZN(n798) );
  XNOR2_X1 U878 ( .A(G166), .B(n802), .ZN(n796) );
  XOR2_X1 U879 ( .A(n937), .B(G305), .Z(n794) );
  XNOR2_X1 U880 ( .A(G288), .B(n794), .ZN(n795) );
  XNOR2_X1 U881 ( .A(n796), .B(n795), .ZN(n797) );
  XNOR2_X1 U882 ( .A(n798), .B(n797), .ZN(n892) );
  XNOR2_X1 U883 ( .A(n892), .B(n799), .ZN(n800) );
  NAND2_X1 U884 ( .A1(n800), .A2(G868), .ZN(n801) );
  XOR2_X1 U885 ( .A(KEYINPUT81), .B(n801), .Z(n804) );
  OR2_X1 U886 ( .A1(n802), .A2(G868), .ZN(n803) );
  NAND2_X1 U887 ( .A1(n804), .A2(n803), .ZN(G295) );
  NAND2_X1 U888 ( .A1(G2078), .A2(G2084), .ZN(n805) );
  XOR2_X1 U889 ( .A(KEYINPUT20), .B(n805), .Z(n806) );
  NAND2_X1 U890 ( .A1(G2090), .A2(n806), .ZN(n807) );
  XNOR2_X1 U891 ( .A(KEYINPUT21), .B(n807), .ZN(n808) );
  NAND2_X1 U892 ( .A1(n808), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U893 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U894 ( .A(KEYINPUT67), .B(G57), .ZN(G237) );
  NAND2_X1 U895 ( .A1(G132), .A2(G82), .ZN(n809) );
  XNOR2_X1 U896 ( .A(n809), .B(KEYINPUT22), .ZN(n810) );
  XNOR2_X1 U897 ( .A(n810), .B(KEYINPUT82), .ZN(n811) );
  NOR2_X1 U898 ( .A1(G218), .A2(n811), .ZN(n812) );
  NAND2_X1 U899 ( .A1(G96), .A2(n812), .ZN(n824) );
  NAND2_X1 U900 ( .A1(n824), .A2(G2106), .ZN(n816) );
  NAND2_X1 U901 ( .A1(G108), .A2(G120), .ZN(n813) );
  NOR2_X1 U902 ( .A1(G237), .A2(n813), .ZN(n814) );
  NAND2_X1 U903 ( .A1(G69), .A2(n814), .ZN(n823) );
  NAND2_X1 U904 ( .A1(G567), .A2(n823), .ZN(n815) );
  NAND2_X1 U905 ( .A1(n816), .A2(n815), .ZN(n847) );
  NAND2_X1 U906 ( .A1(G483), .A2(G661), .ZN(n817) );
  NOR2_X1 U907 ( .A1(n847), .A2(n817), .ZN(n822) );
  NAND2_X1 U908 ( .A1(n822), .A2(G36), .ZN(n818) );
  XOR2_X1 U909 ( .A(KEYINPUT83), .B(n818), .Z(G176) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n819), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n820) );
  NAND2_X1 U912 ( .A1(G661), .A2(n820), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n822), .A2(n821), .ZN(G188) );
  INV_X1 U916 ( .A(G132), .ZN(G219) );
  INV_X1 U917 ( .A(G120), .ZN(G236) );
  INV_X1 U918 ( .A(G108), .ZN(G238) );
  INV_X1 U919 ( .A(G82), .ZN(G220) );
  INV_X1 U920 ( .A(G69), .ZN(G235) );
  NOR2_X1 U921 ( .A1(n824), .A2(n823), .ZN(G325) );
  INV_X1 U922 ( .A(G325), .ZN(G261) );
  XOR2_X1 U923 ( .A(G2096), .B(KEYINPUT43), .Z(n826) );
  XNOR2_X1 U924 ( .A(G2072), .B(G2678), .ZN(n825) );
  XNOR2_X1 U925 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U926 ( .A(n827), .B(KEYINPUT42), .Z(n829) );
  XNOR2_X1 U927 ( .A(G2067), .B(G2090), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U929 ( .A(KEYINPUT104), .B(G2100), .Z(n831) );
  XNOR2_X1 U930 ( .A(G2078), .B(G2084), .ZN(n830) );
  XNOR2_X1 U931 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(G227) );
  XOR2_X1 U933 ( .A(G2474), .B(KEYINPUT106), .Z(n835) );
  XNOR2_X1 U934 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U936 ( .A(n836), .B(KEYINPUT105), .Z(n838) );
  XNOR2_X1 U937 ( .A(G1996), .B(G1991), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n846) );
  XOR2_X1 U939 ( .A(G1981), .B(G1971), .Z(n840) );
  XNOR2_X1 U940 ( .A(G1966), .B(G1956), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U942 ( .A(KEYINPUT107), .B(G1986), .Z(n842) );
  XNOR2_X1 U943 ( .A(G1961), .B(G1976), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U945 ( .A(n844), .B(n843), .Z(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(G229) );
  INV_X1 U947 ( .A(n847), .ZN(G319) );
  NAND2_X1 U948 ( .A1(G124), .A2(n865), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U950 ( .A1(n864), .A2(G112), .ZN(n849) );
  NAND2_X1 U951 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U952 ( .A1(G136), .A2(n869), .ZN(n852) );
  NAND2_X1 U953 ( .A1(G100), .A2(n871), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U955 ( .A1(n854), .A2(n853), .ZN(G162) );
  NAND2_X1 U956 ( .A1(G118), .A2(n864), .ZN(n856) );
  NAND2_X1 U957 ( .A1(G130), .A2(n865), .ZN(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n863) );
  XNOR2_X1 U959 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G142), .A2(n869), .ZN(n858) );
  NAND2_X1 U961 ( .A1(G106), .A2(n871), .ZN(n857) );
  NAND2_X1 U962 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n859), .B(KEYINPUT45), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n861), .B(n860), .ZN(n862) );
  NOR2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n888) );
  NAND2_X1 U966 ( .A1(G115), .A2(n864), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G127), .A2(n865), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U969 ( .A(KEYINPUT47), .B(n868), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G139), .A2(n869), .ZN(n870) );
  XOR2_X1 U971 ( .A(KEYINPUT112), .B(n870), .Z(n874) );
  NAND2_X1 U972 ( .A1(G103), .A2(n871), .ZN(n872) );
  XNOR2_X1 U973 ( .A(KEYINPUT111), .B(n872), .ZN(n873) );
  NOR2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n978) );
  XNOR2_X1 U976 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n877), .B(KEYINPUT46), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(n883) );
  XOR2_X1 U979 ( .A(G162), .B(n970), .Z(n880) );
  XNOR2_X1 U980 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U981 ( .A(n883), .B(n882), .Z(n885) );
  XNOR2_X1 U982 ( .A(G160), .B(G164), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U984 ( .A(n978), .B(n886), .Z(n887) );
  XNOR2_X1 U985 ( .A(n888), .B(n887), .ZN(n890) );
  XOR2_X1 U986 ( .A(n890), .B(n889), .Z(n891) );
  NOR2_X1 U987 ( .A1(G37), .A2(n891), .ZN(G395) );
  XOR2_X1 U988 ( .A(n892), .B(G286), .Z(n895) );
  XNOR2_X1 U989 ( .A(G171), .B(n893), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U991 ( .A1(G37), .A2(n896), .ZN(G397) );
  NOR2_X1 U992 ( .A1(G227), .A2(G229), .ZN(n898) );
  XNOR2_X1 U993 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n910) );
  XOR2_X1 U995 ( .A(KEYINPUT103), .B(G2427), .Z(n900) );
  XNOR2_X1 U996 ( .A(G2435), .B(G2438), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n907) );
  XOR2_X1 U998 ( .A(G2443), .B(G2430), .Z(n902) );
  XNOR2_X1 U999 ( .A(G2454), .B(G2446), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1001 ( .A(n903), .B(G2451), .Z(n905) );
  XNOR2_X1 U1002 ( .A(G1348), .B(G1341), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(n908), .A2(G14), .ZN(n913) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n913), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G96), .ZN(G221) );
  INV_X1 U1012 ( .A(n913), .ZN(G401) );
  INV_X1 U1013 ( .A(KEYINPUT55), .ZN(n992) );
  XNOR2_X1 U1014 ( .A(G2090), .B(G35), .ZN(n928) );
  XNOR2_X1 U1015 ( .A(G2067), .B(G26), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(G1991), .B(G25), .ZN(n914) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(G32), .B(n916), .ZN(n917) );
  NAND2_X1 U1019 ( .A1(n917), .A2(G28), .ZN(n920) );
  XOR2_X1 U1020 ( .A(KEYINPUT119), .B(G2072), .Z(n918) );
  XNOR2_X1 U1021 ( .A(G33), .B(n918), .ZN(n919) );
  NOR2_X1 U1022 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(G27), .B(n923), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(KEYINPUT53), .B(n926), .ZN(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n931) );
  XOR2_X1 U1028 ( .A(G2084), .B(G34), .Z(n929) );
  XNOR2_X1 U1029 ( .A(KEYINPUT54), .B(n929), .ZN(n930) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n992), .B(n932), .ZN(n934) );
  INV_X1 U1032 ( .A(G29), .ZN(n933) );
  NAND2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(G11), .A2(n935), .ZN(n964) );
  XOR2_X1 U1035 ( .A(G16), .B(KEYINPUT56), .Z(n961) );
  XOR2_X1 U1036 ( .A(G1341), .B(KEYINPUT121), .Z(n936) );
  XNOR2_X1 U1037 ( .A(n937), .B(n936), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n946) );
  AND2_X1 U1039 ( .A1(G303), .A2(G1971), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(n944), .B(KEYINPUT120), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n959) );
  XNOR2_X1 U1044 ( .A(n947), .B(G1956), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(G171), .B(G1961), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G1348), .B(n950), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G168), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(n955), .B(KEYINPUT57), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n962), .B(KEYINPUT122), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n996) );
  INV_X1 U1057 ( .A(n965), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n977) );
  XNOR2_X1 U1059 ( .A(G160), .B(G2084), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n968), .B(KEYINPUT115), .ZN(n975) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(n971), .B(KEYINPUT116), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1065 ( .A1(n977), .A2(n976), .ZN(n990) );
  XNOR2_X1 U1066 ( .A(KEYINPUT117), .B(n978), .ZN(n979) );
  XOR2_X1 U1067 ( .A(G2072), .B(n979), .Z(n981) );
  XOR2_X1 U1068 ( .A(G164), .B(G2078), .Z(n980) );
  NOR2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(n982), .B(KEYINPUT118), .ZN(n983) );
  XNOR2_X1 U1071 ( .A(n983), .B(KEYINPUT50), .ZN(n988) );
  XOR2_X1 U1072 ( .A(G2090), .B(G162), .Z(n984) );
  NOR2_X1 U1073 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1074 ( .A(KEYINPUT51), .B(n986), .Z(n987) );
  NAND2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1076 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1077 ( .A(KEYINPUT52), .B(n991), .ZN(n993) );
  NAND2_X1 U1078 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1079 ( .A1(n994), .A2(G29), .ZN(n995) );
  NAND2_X1 U1080 ( .A1(n996), .A2(n995), .ZN(n1024) );
  XOR2_X1 U1081 ( .A(G1961), .B(G5), .Z(n1012) );
  XOR2_X1 U1082 ( .A(G1966), .B(G21), .Z(n997) );
  XNOR2_X1 U1083 ( .A(KEYINPUT125), .B(n997), .ZN(n1009) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(KEYINPUT123), .B(n1000), .Z(n1004) );
  XNOR2_X1 U1088 ( .A(KEYINPUT59), .B(G4), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(n1001), .B(KEYINPUT124), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G1348), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G20), .B(G1956), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1007), .Z(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(KEYINPUT126), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1020) );
  XOR2_X1 U1098 ( .A(G1976), .B(G23), .Z(n1016) );
  XNOR2_X1 U1099 ( .A(G1971), .B(G22), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G24), .B(G1986), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1017), .Z(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT127), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1021), .Z(n1022) );
  NOR2_X1 U1107 ( .A1(G16), .A2(n1022), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(n1025), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

