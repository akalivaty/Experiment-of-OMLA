//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n210), .A2(G20), .A3(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n214), .B1(new_n202), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n205), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n208), .B(new_n213), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n221), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XOR2_X1   g0036(.A(G50), .B(G58), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NAND2_X1  g0042(.A1(G58), .A2(G68), .ZN(new_n243));
  OR2_X1    g0043(.A1(new_n243), .A2(KEYINPUT73), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(KEYINPUT73), .ZN(new_n245));
  OAI211_X1 g0045(.A(new_n244), .B(new_n245), .C1(G58), .C2(G68), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n246), .A2(G20), .B1(G159), .B2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G20), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT7), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT71), .B(G33), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n252), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT7), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n255), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n248), .B1(new_n260), .B2(new_n222), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT16), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT74), .ZN(new_n264));
  INV_X1    g0064(.A(new_n250), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n251), .A2(KEYINPUT71), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT71), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT72), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT72), .A4(KEYINPUT3), .ZN(new_n272));
  AOI21_X1  g0072(.A(G20), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(G68), .B1(new_n273), .B2(new_n258), .ZN(new_n274));
  AOI211_X1 g0074(.A(KEYINPUT7), .B(G20), .C1(new_n271), .C2(new_n272), .ZN(new_n275));
  OAI211_X1 g0075(.A(KEYINPUT16), .B(new_n248), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n211), .B1(new_n205), .B2(new_n251), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT64), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n277), .A2(new_n278), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT74), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n261), .A2(new_n282), .A3(new_n262), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n264), .A2(new_n276), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G1), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n285), .A2(G20), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n287), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT75), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n292), .A2(KEYINPUT75), .A3(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n269), .A2(new_n270), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(new_n272), .A3(new_n250), .ZN(new_n300));
  INV_X1    g0100(.A(G226), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G1698), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(G223), .B2(G1698), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n300), .A2(new_n303), .B1(new_n251), .B2(new_n216), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G41), .ZN(new_n307));
  INV_X1    g0107(.A(G45), .ZN(new_n308));
  AOI21_X1  g0108(.A(G1), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G274), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n310), .A2(new_n305), .A3(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n305), .A2(new_n309), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n312), .B1(G232), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n306), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G200), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n306), .A2(G190), .A3(new_n314), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n284), .A2(new_n298), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT17), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n284), .A2(new_n298), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n315), .A2(G169), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n315), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT18), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT18), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n321), .A2(new_n327), .A3(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n288), .A2(G50), .A3(new_n291), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n251), .A2(G20), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT65), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(new_n289), .ZN(new_n334));
  INV_X1    g0134(.A(G150), .ZN(new_n335));
  INV_X1    g0135(.A(new_n247), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n335), .A2(new_n336), .B1(new_n201), .B2(new_n254), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n281), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n331), .B(new_n338), .C1(G50), .C2(new_n286), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT9), .ZN(new_n340));
  INV_X1    g0140(.A(new_n253), .ZN(new_n341));
  INV_X1    g0141(.A(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G222), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G223), .A2(G1698), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n305), .C1(G77), .C2(new_n341), .ZN(new_n346));
  INV_X1    g0146(.A(new_n312), .ZN(new_n347));
  INV_X1    g0147(.A(new_n313), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n346), .B(new_n347), .C1(new_n301), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G200), .ZN(new_n350));
  INV_X1    g0150(.A(G190), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n340), .B(new_n350), .C1(new_n351), .C2(new_n349), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n352), .B(KEYINPUT10), .ZN(new_n353));
  INV_X1    g0153(.A(G169), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n339), .B(new_n355), .C1(G179), .C2(new_n349), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n288), .A2(G68), .A3(new_n291), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT69), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n247), .A2(G50), .B1(G20), .B2(new_n222), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n333), .B2(new_n202), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n361), .A2(new_n281), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n362), .A2(KEYINPUT11), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(KEYINPUT11), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n287), .A2(new_n222), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT12), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n359), .A2(new_n363), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n312), .B1(G238), .B2(new_n313), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n221), .A2(G1698), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n341), .B(new_n369), .C1(G226), .C2(G1698), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G97), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT68), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n305), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n368), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n354), .A2(KEYINPUT70), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n380), .A2(KEYINPUT14), .B1(new_n323), .B2(new_n378), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n367), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n378), .A2(G200), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n378), .A2(new_n351), .ZN(new_n385));
  OR3_X1    g0185(.A1(new_n384), .A2(new_n385), .A3(new_n367), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n288), .A2(G77), .A3(new_n291), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(G77), .B2(new_n286), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT15), .B(G87), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT66), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n333), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n393), .A2(KEYINPUT67), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n289), .A2(new_n336), .B1(new_n254), .B2(new_n202), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n395), .B1(new_n393), .B2(KEYINPUT67), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n389), .B1(new_n281), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G238), .A2(G1698), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n341), .B(new_n399), .C1(new_n221), .C2(G1698), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n400), .B(new_n305), .C1(G107), .C2(new_n341), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n312), .B1(G244), .B2(new_n313), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n354), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(G179), .B2(new_n403), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n403), .A2(new_n351), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(G200), .B2(new_n403), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n398), .B2(new_n408), .ZN(new_n409));
  AND4_X1   g0209(.A1(new_n330), .A2(new_n357), .A3(new_n387), .A4(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n285), .A2(G45), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT5), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(G41), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT77), .B1(new_n413), .B2(G41), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT77), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n416), .A2(new_n307), .A3(KEYINPUT5), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n374), .A2(new_n414), .A3(G274), .A4(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n305), .B1(new_n414), .B2(new_n418), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(KEYINPUT78), .A3(G257), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT78), .B1(new_n420), .B2(G257), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n419), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n271), .A2(G244), .A3(new_n272), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT4), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G283), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n342), .A2(KEYINPUT4), .A3(G244), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(new_n253), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT4), .B1(new_n253), .B2(new_n217), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(G1698), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n374), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(G200), .B1(new_n424), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G107), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(KEYINPUT6), .A3(G97), .ZN(new_n436));
  INV_X1    g0236(.A(G97), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(new_n435), .ZN(new_n438));
  NOR2_X1   g0238(.A1(G97), .A2(G107), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n436), .B1(new_n440), .B2(KEYINPUT6), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n441), .A2(G20), .B1(G77), .B2(new_n247), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n257), .A2(new_n259), .ZN(new_n443));
  INV_X1    g0243(.A(new_n255), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n435), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n260), .A2(KEYINPUT76), .A3(new_n435), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n281), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n286), .A2(G97), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n285), .A2(G33), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n286), .B(new_n451), .C1(new_n279), .C2(new_n280), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n450), .B1(new_n453), .B2(G97), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n434), .A2(new_n449), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT79), .B1(new_n424), .B2(new_n433), .ZN(new_n456));
  INV_X1    g0256(.A(new_n419), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n414), .A2(new_n418), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(G257), .A3(new_n374), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT78), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(new_n461), .B2(new_n421), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT79), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n431), .A2(G1698), .ZN(new_n464));
  INV_X1    g0264(.A(new_n430), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n426), .B2(new_n425), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n462), .B(new_n463), .C1(new_n467), .C2(new_n374), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n456), .A2(new_n468), .A3(G190), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n455), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n424), .A2(new_n433), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n323), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n449), .A2(new_n454), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(G169), .B1(new_n456), .B2(new_n468), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n287), .A2(KEYINPUT25), .A3(new_n435), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT82), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT25), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n286), .B2(G107), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT83), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n435), .B2(new_n452), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n216), .A2(G20), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT22), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n300), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n256), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT81), .B(G116), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n489), .A3(new_n254), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n254), .A2(G107), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT23), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT22), .ZN(new_n493));
  INV_X1    g0293(.A(new_n484), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n253), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n490), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT24), .B1(new_n486), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n271), .A2(KEYINPUT22), .A3(new_n272), .A4(new_n484), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n492), .A2(new_n495), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT24), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n490), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n483), .B1(new_n502), .B2(new_n281), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n217), .A2(new_n342), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(G257), .B2(new_n342), .ZN(new_n505));
  INV_X1    g0305(.A(G294), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n300), .A2(new_n505), .B1(new_n506), .B2(new_n256), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(new_n305), .B1(G264), .B2(new_n420), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(G190), .A3(new_n419), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n305), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n420), .A2(G264), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n419), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G200), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n503), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n470), .A2(new_n476), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n392), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n286), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT19), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n254), .B1(new_n372), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n216), .A2(new_n437), .A3(new_n435), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n520), .B1(new_n333), .B2(new_n437), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n254), .A2(G68), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(new_n300), .C2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n519), .B1(new_n526), .B2(new_n281), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n453), .A2(G87), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n305), .B1(new_n217), .B2(new_n412), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(G274), .B2(new_n412), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n223), .A2(G1698), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n300), .A2(new_n533), .B1(new_n256), .B2(new_n488), .ZN(new_n534));
  INV_X1    g0334(.A(new_n300), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n535), .A2(KEYINPUT80), .A3(G244), .A4(G1698), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT80), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n425), .B2(new_n342), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n534), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(G190), .B(new_n531), .C1(new_n539), .C2(new_n374), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n529), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n531), .B1(new_n539), .B2(new_n374), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G200), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n536), .A2(new_n538), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n305), .B1(new_n545), .B2(new_n534), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(new_n323), .A3(new_n531), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n542), .A2(new_n354), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n527), .B1(new_n392), .B2(new_n452), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  MUX2_X1   g0351(.A(G257), .B(G264), .S(G1698), .Z(new_n552));
  NAND3_X1  g0352(.A1(new_n271), .A2(new_n272), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n253), .A2(G303), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n374), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n420), .A2(G270), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n419), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n488), .A2(new_n287), .ZN(new_n559));
  INV_X1    g0359(.A(G116), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n428), .B(new_n254), .C1(G33), .C2(new_n437), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n561), .A2(new_n277), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n488), .A2(G20), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT20), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n277), .A3(new_n561), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT20), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI221_X1 g0367(.A(new_n559), .B1(new_n452), .B2(new_n560), .C1(new_n564), .C2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n558), .A2(new_n568), .A3(KEYINPUT21), .A4(G169), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n555), .A2(new_n557), .A3(new_n323), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n568), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n568), .B1(new_n558), .B2(G200), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n351), .B2(new_n558), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n512), .A2(new_n354), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n508), .A2(new_n323), .A3(new_n419), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n279), .A2(new_n280), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n497), .B2(new_n501), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n575), .B(new_n576), .C1(new_n578), .C2(new_n483), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n559), .B1(new_n567), .B2(new_n564), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n452), .A2(new_n560), .ZN(new_n582));
  OAI21_X1  g0382(.A(G169), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n555), .A2(new_n557), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n572), .A2(new_n574), .A3(new_n579), .A4(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n551), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n411), .A2(new_n517), .A3(new_n588), .ZN(G372));
  INV_X1    g0389(.A(KEYINPUT85), .ZN(new_n590));
  INV_X1    g0390(.A(new_n328), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n327), .B1(new_n321), .B2(new_n324), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n326), .A2(KEYINPUT85), .A3(new_n328), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT86), .B1(new_n398), .B2(new_n405), .ZN(new_n597));
  OR3_X1    g0397(.A1(new_n398), .A2(KEYINPUT86), .A3(new_n405), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n386), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n320), .B1(new_n599), .B2(new_n383), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n353), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n601), .A2(new_n356), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n456), .A2(new_n468), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n354), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n323), .A2(new_n471), .B1(new_n449), .B2(new_n454), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n323), .A2(new_n510), .A3(new_n419), .A4(new_n511), .ZN(new_n607));
  AOI21_X1  g0407(.A(G169), .B1(new_n508), .B2(new_n419), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n503), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n585), .A2(new_n569), .A3(new_n571), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n514), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n606), .B1(new_n611), .B2(new_n470), .ZN(new_n612));
  OR3_X1    g0412(.A1(new_n539), .A2(KEYINPUT84), .A3(new_n374), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT84), .B1(new_n539), .B2(new_n374), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n531), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G200), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT26), .B1(new_n616), .B2(new_n541), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n547), .A2(new_n549), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n354), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n612), .A2(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n544), .A2(new_n476), .A3(new_n550), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT26), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n602), .B1(new_n411), .B2(new_n624), .ZN(G369));
  NAND3_X1  g0425(.A1(new_n285), .A2(new_n254), .A3(G13), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(G213), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n630), .A2(KEYINPUT87), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(KEYINPUT87), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(G343), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n503), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n579), .B1(new_n515), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n609), .A2(new_n636), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n610), .A2(new_n636), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n609), .B2(new_n636), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n635), .A2(new_n568), .ZN(new_n644));
  XOR2_X1   g0444(.A(new_n610), .B(new_n644), .Z(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n574), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G330), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n643), .B1(new_n648), .B2(new_n640), .ZN(G399));
  INV_X1    g0449(.A(new_n206), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(G41), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n522), .A2(G116), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G1), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n209), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT29), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n619), .A2(new_n618), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n604), .A2(new_n605), .B1(new_n455), .B2(new_n469), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT89), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n609), .B2(new_n610), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n572), .A2(new_n579), .A3(KEYINPUT89), .A4(new_n585), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n659), .A2(new_n661), .A3(new_n514), .A4(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n616), .A2(new_n541), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n658), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n616), .A2(new_n541), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n606), .A2(new_n666), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n666), .A2(new_n621), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n657), .B1(new_n670), .B2(new_n636), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n623), .A2(new_n636), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(KEYINPUT29), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n512), .A2(new_n558), .A3(new_n323), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n471), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n615), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT30), .ZN(new_n678));
  INV_X1    g0478(.A(new_n603), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n570), .A2(new_n508), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n542), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NOR4_X1   g0482(.A1(new_n603), .A2(new_n542), .A3(KEYINPUT30), .A4(new_n680), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n677), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT88), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT31), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n570), .A2(new_n508), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n546), .A2(new_n688), .A3(new_n531), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT30), .B1(new_n689), .B2(new_n603), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n679), .A2(new_n681), .A3(new_n678), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(KEYINPUT88), .A3(new_n677), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n686), .A2(new_n687), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n635), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n687), .B1(new_n587), .B2(new_n516), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n684), .A2(KEYINPUT31), .A3(new_n635), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n674), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n656), .B1(new_n703), .B2(G1), .ZN(G364));
  INV_X1    g0504(.A(G13), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G20), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G45), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n652), .A2(G1), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n648), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n646), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G13), .A2(G33), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n646), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n708), .B(KEYINPUT90), .Z(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n211), .B1(G20), .B2(new_n354), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n351), .A2(G200), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n254), .B1(new_n720), .B2(new_n323), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n254), .A2(new_n323), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n351), .A3(G200), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI22_X1  g0525(.A1(G97), .A2(new_n722), .B1(new_n725), .B2(G68), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n254), .A2(new_n323), .A3(KEYINPUT92), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n720), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n726), .B1(new_n733), .B2(new_n220), .ZN(new_n734));
  INV_X1    g0534(.A(new_n730), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G190), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n734), .B1(G77), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n254), .A2(G179), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(G190), .A3(G200), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n341), .B1(new_n741), .B2(new_n216), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(KEYINPUT94), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n740), .A2(new_n351), .A3(G200), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G107), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n740), .A2(new_n736), .ZN(new_n747));
  INV_X1    g0547(.A(G159), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT32), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n747), .A2(KEYINPUT32), .A3(new_n748), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n743), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n723), .A2(G190), .A3(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT93), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n753), .A2(KEYINPUT93), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n758), .A2(G50), .B1(KEYINPUT94), .B2(new_n742), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n739), .A2(new_n752), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n747), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n341), .B1(new_n761), .B2(G329), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n763), .B2(new_n744), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(G322), .B2(new_n732), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n758), .A2(G326), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n738), .A2(G311), .ZN(new_n767));
  INV_X1    g0567(.A(G303), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n721), .A2(new_n506), .B1(new_n741), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(KEYINPUT33), .B(G317), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(new_n725), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n765), .A2(new_n766), .A3(new_n767), .A4(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n719), .B1(new_n760), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n714), .A2(new_n718), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n238), .A2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT91), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n775), .A2(new_n776), .B1(new_n308), .B2(new_n210), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n535), .A2(new_n650), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n777), .B(new_n778), .C1(new_n776), .C2(new_n775), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n650), .A2(new_n253), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n780), .A2(G355), .B1(new_n560), .B2(new_n650), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n717), .B(new_n773), .C1(new_n774), .C2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n711), .B1(new_n715), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(G396));
  INV_X1    g0585(.A(new_n708), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n398), .A2(new_n636), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n598), .A2(new_n597), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(KEYINPUT98), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n409), .B1(new_n398), .B2(new_n636), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT98), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n598), .A2(new_n791), .A3(new_n597), .A4(new_n787), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n672), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n635), .B1(new_n620), .B2(new_n622), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n793), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n786), .B1(new_n701), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n701), .B2(new_n798), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n719), .A2(new_n713), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n716), .B1(G77), .B2(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n732), .A2(G294), .B1(G97), .B2(new_n722), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT95), .Z(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n253), .B1(new_n747), .B2(new_n805), .C1(new_n724), .C2(new_n763), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n745), .A2(G87), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n435), .B2(new_n741), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n806), .B(new_n808), .C1(new_n738), .C2(new_n489), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n804), .B(new_n809), .C1(new_n768), .C2(new_n757), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n757), .A2(new_n811), .B1(new_n335), .B2(new_n724), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT96), .ZN(new_n813));
  INV_X1    g0613(.A(G143), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n814), .B2(new_n733), .C1(new_n748), .C2(new_n737), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT34), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT97), .ZN(new_n818));
  INV_X1    g0618(.A(new_n741), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n819), .A2(G50), .B1(new_n761), .B2(G132), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n744), .A2(new_n222), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(G58), .B2(new_n722), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n818), .A2(new_n535), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n817), .A2(KEYINPUT97), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n810), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n802), .B1(new_n825), .B2(new_n718), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n713), .B2(new_n793), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n800), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G384));
  NOR2_X1   g0629(.A1(new_n706), .A2(new_n285), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT105), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n367), .A2(new_n635), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n383), .A2(new_n386), .A3(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n367), .B(new_n635), .C1(new_n381), .C2(new_n382), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n835), .A2(new_n793), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n696), .B1(new_n694), .B2(new_n635), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n686), .A2(new_n693), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n635), .A2(KEYINPUT31), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n836), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n276), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n248), .B1(new_n274), .B2(new_n275), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n577), .B1(new_n843), .B2(new_n262), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n842), .B1(new_n844), .B2(KEYINPUT102), .ZN(new_n845));
  INV_X1    g0645(.A(new_n248), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n300), .A2(new_n254), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n222), .B1(new_n847), .B2(KEYINPUT7), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n273), .A2(new_n258), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n281), .B1(new_n850), .B2(KEYINPUT16), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT102), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n294), .B1(new_n845), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(new_n633), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n320), .B2(new_n329), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  INV_X1    g0657(.A(new_n318), .ZN(new_n858));
  INV_X1    g0658(.A(new_n294), .ZN(new_n859));
  OAI211_X1 g0659(.A(KEYINPUT102), .B(new_n281), .C1(new_n850), .C2(KEYINPUT16), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n276), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n844), .A2(KEYINPUT102), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n858), .B1(new_n863), .B2(new_n324), .ZN(new_n864));
  INV_X1    g0664(.A(new_n633), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n857), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n321), .A2(new_n865), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n325), .A2(new_n868), .A3(new_n318), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n856), .B(KEYINPUT38), .C1(new_n867), .C2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n324), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n318), .B1(new_n854), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n874), .B2(new_n855), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n325), .A2(new_n868), .A3(new_n318), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n857), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n878), .B2(new_n856), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT103), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n863), .A2(new_n324), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n866), .A2(new_n882), .A3(new_n318), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n870), .B1(new_n883), .B2(KEYINPUT37), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n591), .A2(new_n592), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n318), .B(KEYINPUT17), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n866), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n881), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT103), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n871), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n841), .B1(new_n880), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n831), .B1(new_n891), .B2(KEYINPUT40), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n835), .A2(new_n793), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n838), .A2(new_n839), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n894), .B2(new_n698), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n888), .A2(new_n889), .A3(new_n871), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n889), .B1(new_n888), .B2(new_n871), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(KEYINPUT105), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT104), .B1(new_n869), .B2(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n877), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n876), .A2(KEYINPUT104), .A3(new_n857), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n593), .A2(new_n594), .A3(new_n886), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n321), .A3(new_n865), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT40), .B1(new_n907), .B2(new_n872), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n892), .A2(new_n900), .B1(new_n895), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n837), .A2(new_n840), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n411), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n710), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n910), .B2(new_n912), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n796), .A2(new_n793), .B1(new_n406), .B2(new_n636), .ZN(new_n915));
  INV_X1    g0715(.A(new_n835), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n915), .B(new_n916), .C1(new_n880), .C2(new_n890), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n383), .A2(new_n635), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n868), .B1(new_n595), .B2(new_n886), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n902), .A2(new_n903), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n881), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n922), .A3(new_n871), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT39), .B1(new_n872), .B2(new_n879), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n595), .A2(new_n865), .ZN(new_n926));
  NOR3_X1   g0726(.A1(new_n917), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n410), .B1(new_n671), .B2(new_n673), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n602), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n927), .B(new_n929), .Z(new_n930));
  AOI21_X1  g0730(.A(new_n830), .B1(new_n914), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n930), .B2(new_n914), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n441), .A2(KEYINPUT35), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n441), .A2(KEYINPUT35), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n211), .A2(new_n254), .A3(new_n560), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT99), .Z(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(KEYINPUT36), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(KEYINPUT36), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n244), .A2(G77), .A3(new_n210), .A4(new_n245), .ZN(new_n941));
  INV_X1    g0741(.A(G50), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n941), .A2(KEYINPUT100), .B1(new_n942), .B2(G68), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(KEYINPUT100), .B2(new_n941), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(G1), .A3(new_n705), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT101), .Z(new_n946));
  NAND4_X1  g0746(.A1(new_n932), .A2(new_n939), .A3(new_n940), .A4(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT106), .ZN(G367));
  NAND2_X1  g0748(.A1(new_n658), .A2(new_n667), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n529), .A2(new_n636), .ZN(new_n950));
  MUX2_X1   g0750(.A(new_n949), .B(new_n658), .S(new_n950), .Z(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n714), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT46), .B1(new_n819), .B2(new_n489), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n722), .A2(G107), .B1(new_n761), .B2(G317), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n737), .B2(new_n763), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n953), .B(new_n955), .C1(G303), .C2(new_n732), .ZN(new_n956));
  AOI22_X1  g0756(.A1(G294), .A2(new_n725), .B1(new_n745), .B2(G97), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n819), .A2(KEYINPUT46), .A3(G116), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n957), .A2(new_n300), .A3(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n956), .B(new_n959), .C1(new_n805), .C2(new_n757), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n732), .A2(G150), .B1(G68), .B2(new_n722), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n814), .B2(new_n757), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(KEYINPUT109), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(KEYINPUT109), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n341), .B1(new_n747), .B2(new_n811), .C1(new_n202), .C2(new_n744), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n724), .A2(new_n748), .B1(new_n741), .B2(new_n220), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n965), .B(new_n966), .C1(new_n738), .C2(G50), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n963), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n960), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n718), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n778), .A2(new_n234), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n972), .B(new_n774), .C1(new_n206), .C2(new_n392), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n952), .A2(new_n716), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n707), .A2(G1), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n473), .A2(new_n635), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n659), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n606), .B2(new_n636), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n643), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT108), .Z(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n979), .B(KEYINPUT108), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n643), .A2(new_n978), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT45), .Z(new_n986));
  NAND3_X1  g0786(.A1(new_n982), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n648), .A2(new_n640), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n640), .B(new_n641), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n648), .B(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n703), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n651), .B(KEYINPUT41), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n975), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT43), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n951), .A2(new_n996), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n642), .A2(new_n978), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT107), .Z(new_n1001));
  OAI21_X1  g0801(.A(new_n606), .B1(new_n977), .B2(new_n579), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n999), .A2(KEYINPUT42), .B1(new_n636), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n997), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n951), .A2(new_n996), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n988), .A2(new_n978), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n974), .B1(new_n995), .B2(new_n1008), .ZN(G387));
  NAND2_X1  g0809(.A1(new_n231), .A2(G45), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT110), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n653), .B(new_n308), .C1(new_n222), .C2(new_n202), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1012), .A2(KEYINPUT111), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(KEYINPUT111), .ZN(new_n1014));
  OR3_X1    g0814(.A1(new_n289), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1015));
  OAI21_X1  g0815(.A(KEYINPUT50), .B1(new_n289), .B2(G50), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AND3_X1   g0817(.A1(new_n1011), .A2(new_n778), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n780), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1019), .A2(new_n653), .B1(G107), .B2(new_n206), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n774), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n721), .A2(new_n763), .B1(new_n741), .B2(new_n506), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n732), .A2(G317), .B1(G311), .B2(new_n725), .ZN(new_n1023));
  INV_X1    g0823(.A(G322), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1023), .B1(new_n768), .B2(new_n737), .C1(new_n1024), .C2(new_n757), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1022), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n1026), .B2(new_n1025), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT49), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n744), .A2(new_n488), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1031), .B(new_n535), .C1(G326), .C2(new_n761), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n392), .A2(new_n721), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n738), .B2(G68), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n942), .B2(new_n733), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n724), .A2(new_n289), .B1(new_n741), .B2(new_n202), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n744), .A2(new_n437), .B1(new_n747), .B2(new_n335), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n300), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n748), .B2(new_n757), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1030), .A2(new_n1033), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n718), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1021), .A2(new_n716), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n640), .B2(new_n714), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n991), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1044), .B1(new_n1045), .B2(new_n975), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n703), .A2(new_n1045), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n702), .A2(KEYINPUT112), .A3(new_n991), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n651), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT112), .B1(new_n702), .B2(new_n991), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(G393));
  NAND2_X1  g0851(.A1(new_n778), .A2(new_n241), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n774), .C1(new_n437), .C2(new_n206), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n716), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT113), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n758), .A2(G317), .B1(G311), .B2(new_n732), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT52), .Z(new_n1057));
  AOI22_X1  g0857(.A1(new_n489), .A2(new_n722), .B1(new_n725), .B2(G303), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1058), .A2(new_n253), .A3(new_n746), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G294), .B2(new_n738), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n741), .A2(new_n763), .B1(new_n747), .B2(new_n1024), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT114), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n733), .A2(new_n748), .B1(new_n757), .B2(new_n335), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT51), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n807), .B1(new_n814), .B2(new_n747), .C1(new_n737), .C2(new_n289), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n721), .A2(new_n202), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n724), .A2(new_n942), .B1(new_n741), .B2(new_n222), .ZN(new_n1068));
  NOR4_X1   g0868(.A1(new_n1066), .A2(new_n300), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1057), .A2(new_n1063), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n714), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1055), .B1(new_n719), .B2(new_n1070), .C1(new_n978), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n975), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n989), .A2(new_n1047), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n651), .B1(new_n989), .B2(new_n1047), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1072), .B1(new_n1073), .B2(new_n989), .C1(new_n1074), .C2(new_n1075), .ZN(G390));
  NAND2_X1  g0876(.A1(new_n894), .A2(new_n698), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(G330), .A3(new_n793), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n916), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n700), .A2(G330), .A3(new_n793), .A4(new_n835), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n636), .B(new_n793), .C1(new_n665), .C2(new_n669), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n406), .A2(new_n636), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT115), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT115), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1081), .A2(new_n1085), .A3(new_n1082), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1079), .A2(new_n1080), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1077), .A2(G330), .A3(new_n836), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n700), .A2(G330), .A3(new_n793), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n916), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1088), .B1(new_n915), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1077), .A2(G330), .A3(new_n410), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n928), .A2(new_n602), .A3(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT116), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1084), .A2(new_n835), .A3(new_n1086), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n918), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n921), .B2(new_n871), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n918), .B1(new_n915), .B2(new_n916), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n923), .A3(new_n924), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1101), .A2(new_n1103), .A3(new_n1080), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1089), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n652), .B1(new_n1097), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1106), .A2(new_n975), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n716), .B1(new_n290), .B2(new_n801), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n758), .A2(G128), .B1(G132), .B2(new_n732), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT119), .Z(new_n1114));
  NAND2_X1  g0914(.A1(new_n761), .A2(G125), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n341), .B1(new_n744), .B2(new_n942), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT117), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1117), .B2(new_n1116), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT118), .Z(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n741), .B2(new_n335), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n811), .B2(new_n724), .C1(new_n748), .C2(new_n721), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n819), .A2(new_n1121), .A3(G150), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT54), .B(G143), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1125), .B1(new_n737), .B2(new_n1126), .ZN(new_n1127));
  NOR4_X1   g0927(.A1(new_n1114), .A2(new_n1120), .A3(new_n1124), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1129), .A2(KEYINPUT121), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n758), .A2(G283), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n738), .A2(G97), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n253), .B1(new_n747), .B2(new_n506), .C1(new_n216), .C2(new_n741), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G116), .B2(new_n732), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n821), .B(new_n1067), .C1(G107), .C2(new_n725), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1129), .A2(KEYINPUT121), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1130), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1112), .B1(new_n1138), .B2(new_n718), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT122), .Z(new_n1140));
  AND2_X1   g0940(.A1(new_n923), .A2(new_n924), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1140), .B1(new_n1142), .B2(new_n713), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1111), .A2(KEYINPUT123), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT123), .B1(new_n1111), .B2(new_n1143), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1110), .B1(new_n1144), .B2(new_n1145), .ZN(G378));
  INV_X1    g0946(.A(KEYINPUT116), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1095), .B(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n1106), .B2(new_n1093), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n927), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n357), .B(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n339), .A2(new_n865), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n892), .A2(new_n900), .ZN(new_n1156));
  OAI21_X1  g0956(.A(G330), .B1(new_n908), .B2(new_n841), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1155), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1154), .B(new_n1157), .C1(new_n892), .C2(new_n900), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1150), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n891), .A2(new_n831), .A3(KEYINPUT40), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT105), .B1(new_n898), .B2(new_n899), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1158), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1154), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1156), .A2(new_n1158), .A3(new_n1155), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n1166), .A3(new_n927), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1149), .B1(new_n1161), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n651), .B1(new_n1168), .B2(KEYINPUT57), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1170), .B(new_n1149), .C1(new_n1161), .C2(new_n1167), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1073), .B1(new_n1161), .B2(new_n1167), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1154), .A2(new_n712), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n786), .B1(G50), .B2(new_n801), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n535), .A2(G41), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G50), .B(new_n1176), .C1(new_n251), .C2(new_n307), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G97), .A2(new_n725), .B1(new_n819), .B2(G77), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n220), .B2(new_n744), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G116), .B2(new_n758), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n721), .A2(new_n222), .B1(new_n747), .B2(new_n763), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n738), .B2(new_n518), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n732), .A2(G107), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1182), .A3(new_n1176), .A4(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT58), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1177), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G150), .A2(new_n722), .B1(new_n725), .B2(G132), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n737), .B2(new_n811), .ZN(new_n1189));
  INV_X1    g0989(.A(G128), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n733), .A2(new_n1190), .B1(new_n741), .B2(new_n1126), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT124), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1189), .B(new_n1192), .C1(G125), .C2(new_n758), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT59), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1187), .B1(new_n748), .B2(new_n744), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1186), .B1(new_n1185), .B2(new_n1184), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1175), .B1(new_n1197), .B2(new_n718), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1174), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT125), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1173), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1172), .A2(new_n1201), .ZN(G375));
  AOI22_X1  g1002(.A1(new_n738), .A2(G107), .B1(new_n489), .B2(new_n725), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n506), .B2(new_n757), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n1204), .B(KEYINPUT126), .Z(new_n1205));
  NOR2_X1   g1005(.A1(new_n741), .A2(new_n437), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n253), .B1(new_n747), .B2(new_n768), .C1(new_n202), .C2(new_n744), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n733), .A2(new_n763), .B1(new_n392), .B2(new_n721), .ZN(new_n1208));
  NOR4_X1   g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n722), .A2(G50), .B1(new_n819), .B2(G159), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n535), .B(new_n1210), .C1(new_n724), .C2(new_n1126), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n744), .A2(new_n220), .B1(new_n747), .B2(new_n1190), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n738), .B2(G150), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n811), .B2(new_n733), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1211), .B(new_n1214), .C1(G132), .C2(new_n758), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n718), .B1(new_n1209), .B2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1216), .B(new_n716), .C1(G68), .C2(new_n801), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n916), .B2(new_n712), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1093), .B2(new_n975), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1097), .A2(new_n994), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1220), .B2(new_n1221), .ZN(G381));
  OR2_X1    g1022(.A1(G387), .A2(G390), .ZN(new_n1223));
  OR2_X1    g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1223), .A2(G384), .A3(G381), .A4(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(G378), .ZN(new_n1226));
  INV_X1    g1026(.A(G375), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(G407));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1226), .ZN(new_n1229));
  OAI211_X1 g1029(.A(G407), .B(G213), .C1(G343), .C2(new_n1229), .ZN(G409));
  NAND2_X1  g1030(.A1(new_n634), .A2(G213), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1221), .A2(KEYINPUT60), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(new_n651), .A3(new_n1097), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1221), .A2(KEYINPUT60), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1219), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n828), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G384), .B(new_n1219), .C1(new_n1233), .C2(new_n1234), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n993), .B(new_n1149), .C1(new_n1161), .C2(new_n1167), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1159), .A2(new_n1160), .A3(new_n1150), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n927), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n975), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1199), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1240), .B1(new_n1244), .B2(KEYINPUT127), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT127), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1246), .A3(new_n1199), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G378), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G378), .B(new_n1201), .C1(new_n1169), .C2(new_n1171), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1231), .B(new_n1239), .C1(new_n1248), .C2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT62), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1231), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n634), .A2(G213), .A3(G2897), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1236), .A2(new_n1237), .A3(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1254), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1253), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1199), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT127), .B1(new_n1173), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1168), .A2(new_n994), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1247), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1226), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1249), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT62), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1231), .A4(new_n1239), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1252), .A2(new_n1258), .A3(new_n1259), .A4(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(new_n784), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G387), .A2(G390), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1223), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1270), .B1(new_n1223), .B2(new_n1271), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1268), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1257), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1251), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1265), .A2(KEYINPUT63), .A3(new_n1231), .A4(new_n1239), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1277), .A2(new_n1274), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1276), .A2(new_n1281), .ZN(G405));
  NAND2_X1  g1082(.A1(G375), .A2(new_n1226), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1249), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1239), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1238), .A3(new_n1249), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1275), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1285), .A2(new_n1274), .A3(new_n1286), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(G402));
endmodule


