//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n188));
  OR3_X1    g002(.A1(new_n188), .A2(KEYINPUT2), .A3(G113), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(KEYINPUT2), .B2(G113), .ZN(new_n190));
  AOI22_X1  g004(.A1(new_n189), .A2(new_n190), .B1(KEYINPUT2), .B2(G113), .ZN(new_n191));
  XNOR2_X1  g005(.A(G116), .B(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G116), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT68), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n192), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n193), .B1(new_n202), .B2(new_n191), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n204), .A2(new_n205), .A3(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(KEYINPUT64), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT64), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G134), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n209), .A3(G137), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n206), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT66), .A4(G137), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT64), .B(G134), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n204), .B1(new_n214), .B2(G137), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT65), .B(G131), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n213), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(G137), .B1(new_n207), .B2(new_n209), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n205), .A2(G137), .ZN(new_n219));
  OAI21_X1  g033(.A(G131), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT1), .B1(new_n223), .B2(G146), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(G146), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(G143), .ZN(new_n227));
  OAI211_X1 g041(.A(G128), .B(new_n224), .C1(new_n225), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n223), .A2(G146), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n229), .B(new_n230), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n228), .A2(KEYINPUT70), .A3(new_n232), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n203), .B1(new_n222), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n210), .A2(new_n211), .ZN(new_n239));
  INV_X1    g053(.A(new_n206), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n213), .B1(new_n218), .B2(KEYINPUT11), .ZN(new_n242));
  OAI21_X1  g056(.A(G131), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n217), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT0), .A4(G128), .ZN(new_n245));
  XNOR2_X1  g059(.A(G143), .B(G146), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n238), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n222), .A2(new_n237), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n248), .B1(new_n243), .B2(new_n217), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT69), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT69), .B1(new_n244), .B2(new_n249), .ZN(new_n260));
  AOI211_X1 g074(.A(new_n254), .B(new_n248), .C1(new_n243), .C2(new_n217), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n259), .A2(new_n203), .B1(new_n262), .B2(new_n238), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n253), .B1(new_n263), .B2(new_n252), .ZN(new_n264));
  INV_X1    g078(.A(G210), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n265), .A2(G237), .A3(G953), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n266), .B(KEYINPUT27), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT26), .B(G101), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n267), .B(new_n268), .Z(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT29), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n187), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT76), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n255), .A2(new_n238), .A3(new_n258), .ZN(new_n273));
  INV_X1    g087(.A(new_n233), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n217), .A2(new_n274), .A3(new_n220), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n203), .B1(new_n257), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n252), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n253), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI211_X1 g093(.A(KEYINPUT72), .B(new_n252), .C1(new_n273), .C2(new_n276), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n269), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n228), .A2(KEYINPUT70), .A3(new_n232), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT70), .B1(new_n228), .B2(new_n232), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT30), .B1(new_n221), .B2(new_n284), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n260), .A2(new_n261), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n257), .B2(new_n275), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n203), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n238), .B2(new_n262), .ZN(new_n291));
  INV_X1    g105(.A(new_n269), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT29), .B1(new_n281), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G472), .B1(new_n272), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n292), .B1(new_n279), .B2(new_n280), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n269), .B(new_n273), .C1(new_n286), .C2(new_n289), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT71), .B1(new_n297), .B2(KEYINPUT31), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(KEYINPUT31), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(KEYINPUT71), .A3(KEYINPUT31), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n296), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(G472), .A2(G902), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(KEYINPUT32), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n295), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n303), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n302), .A2(KEYINPUT73), .A3(new_n303), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT74), .B(KEYINPUT32), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT75), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n308), .A2(new_n313), .A3(new_n309), .A4(new_n310), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n305), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G125), .B(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT16), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n226), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n317), .A2(G146), .A3(new_n320), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n194), .B2(G128), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n231), .A2(KEYINPUT23), .A3(G119), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(new_n327), .C1(G119), .C2(new_n231), .ZN(new_n328));
  XNOR2_X1  g142(.A(G119), .B(G128), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT24), .B(G110), .Z(new_n330));
  AOI22_X1  g144(.A1(new_n328), .A2(G110), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n324), .A2(new_n331), .ZN(new_n332));
  OAI22_X1  g146(.A1(new_n328), .A2(G110), .B1(new_n329), .B2(new_n330), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n316), .A2(new_n226), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n323), .A3(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT22), .B(G137), .ZN(new_n337));
  INV_X1    g151(.A(G953), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(G221), .A3(G234), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n337), .B(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(new_n340), .B(KEYINPUT77), .Z(new_n342));
  OAI21_X1  g156(.A(new_n341), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(G902), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT25), .ZN(new_n345));
  INV_X1    g159(.A(G217), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(G234), .B2(new_n187), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n343), .A2(G902), .A3(new_n347), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n315), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G469), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n338), .A2(G227), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n354), .B(KEYINPUT78), .ZN(new_n355));
  XNOR2_X1  g169(.A(G110), .B(G140), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G107), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT79), .A3(G104), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT3), .ZN(new_n360));
  INV_X1    g174(.A(G101), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n362), .A2(new_n358), .A3(KEYINPUT79), .A4(G104), .ZN(new_n363));
  INV_X1    g177(.A(G104), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G107), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n360), .A2(new_n361), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n364), .A2(G107), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n358), .A2(G104), .ZN(new_n368));
  OAI21_X1  g182(.A(G101), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT10), .B1(new_n371), .B2(new_n274), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n360), .A2(new_n363), .A3(new_n365), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G101), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n366), .A2(KEYINPUT4), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n368), .B1(KEYINPUT3), .B2(new_n359), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n361), .B1(new_n377), .B2(new_n363), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n249), .B(new_n375), .C1(new_n376), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT80), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n373), .A2(G101), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(KEYINPUT4), .A3(new_n366), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n249), .A4(new_n375), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n372), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n366), .A2(KEYINPUT10), .A3(new_n369), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT81), .B1(new_n284), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n237), .A2(new_n388), .A3(KEYINPUT10), .A4(new_n371), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT84), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n244), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n244), .A2(KEYINPUT82), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n243), .B2(new_n217), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n390), .A3(new_n385), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n357), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n357), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n370), .B(new_n233), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n403), .B(new_n244), .C1(KEYINPUT83), .C2(KEYINPUT12), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT12), .B1(new_n244), .B2(KEYINPUT83), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n244), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n402), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n353), .B(new_n187), .C1(new_n401), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n404), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n400), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n357), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n385), .A2(new_n390), .A3(new_n393), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n393), .B1(new_n385), .B2(new_n390), .ZN(new_n415));
  INV_X1    g229(.A(new_n244), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n413), .B(G469), .C1(new_n417), .C2(new_n402), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n353), .A2(new_n187), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n409), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT9), .B(G234), .ZN(new_n422));
  OAI21_X1  g236(.A(G221), .B1(new_n422), .B2(G902), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G214), .B1(G237), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G122), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT5), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n199), .B2(new_n201), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n432));
  OAI21_X1  g246(.A(G113), .B1(new_n195), .B2(KEYINPUT5), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT86), .B1(new_n430), .B2(new_n433), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n435), .A2(new_n436), .A3(new_n193), .A4(new_n371), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n203), .A2(new_n382), .A3(new_n375), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(KEYINPUT85), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(KEYINPUT85), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n428), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n438), .A2(KEYINPUT85), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n443), .A2(new_n427), .A3(new_n440), .A4(new_n437), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(KEYINPUT6), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n446), .B(new_n428), .C1(new_n439), .C2(new_n441), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n248), .A2(G125), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n274), .B2(G125), .ZN(new_n449));
  MUX2_X1   g263(.A(new_n448), .B(new_n449), .S(KEYINPUT87), .Z(new_n450));
  INV_X1    g264(.A(G224), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(G953), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n450), .B(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n445), .A2(new_n447), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT7), .B1(new_n451), .B2(G953), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n450), .B2(new_n455), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n435), .A2(new_n436), .A3(new_n193), .A4(new_n370), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n427), .B(KEYINPUT8), .Z(new_n459));
  OAI21_X1  g273(.A(new_n434), .B1(new_n429), .B2(new_n198), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n193), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n459), .B1(new_n461), .B2(new_n371), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(G902), .B1(new_n464), .B2(new_n444), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n454), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G210), .B1(G237), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n454), .A2(new_n467), .A3(new_n465), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n426), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n424), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G237), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n338), .A3(G214), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(new_n223), .ZN(new_n475));
  INV_X1    g289(.A(new_n216), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n475), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n216), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT17), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(KEYINPUT88), .A3(new_n476), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n479), .A2(new_n481), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n324), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n479), .A2(new_n483), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n484), .B(new_n485), .C1(new_n486), .C2(new_n482), .ZN(new_n487));
  XNOR2_X1  g301(.A(G113), .B(G122), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(new_n364), .ZN(new_n489));
  NAND2_X1  g303(.A1(KEYINPUT18), .A2(G131), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n480), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n475), .A2(KEYINPUT18), .A3(G131), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n316), .B(new_n226), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n487), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n489), .B1(new_n487), .B2(new_n494), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n187), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G475), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n479), .A2(new_n483), .A3(new_n481), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n316), .A2(KEYINPUT89), .ZN(new_n501));
  XOR2_X1   g315(.A(new_n501), .B(KEYINPUT19), .Z(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n226), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n503), .A3(new_n323), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n504), .A2(new_n494), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n495), .B1(new_n505), .B2(new_n489), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n507));
  NOR2_X1   g321(.A1(G475), .A2(G902), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT90), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n506), .B2(new_n509), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n499), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G128), .B(G143), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT92), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n214), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT93), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n196), .A2(G122), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT91), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n196), .A2(G122), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n358), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(G107), .A3(new_n523), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(KEYINPUT14), .A3(G107), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n522), .A2(KEYINPUT14), .A3(G107), .A4(new_n523), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT93), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n517), .A2(new_n518), .A3(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n520), .A2(new_n528), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n513), .A2(KEYINPUT13), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n223), .A2(G128), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n533), .B(G134), .C1(KEYINPUT13), .C2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n517), .A2(new_n525), .A3(new_n526), .A4(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n422), .A2(new_n346), .A3(G953), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n532), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n532), .B2(new_n536), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n187), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G478), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n542), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n187), .B(new_n544), .C1(new_n538), .C2(new_n539), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n512), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G952), .ZN(new_n548));
  AOI211_X1 g362(.A(G953), .B(new_n548), .C1(G234), .C2(G237), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT21), .B(G898), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(KEYINPUT94), .ZN(new_n552));
  AOI211_X1 g366(.A(new_n187), .B(new_n338), .C1(G234), .C2(G237), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n550), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n547), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n472), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n352), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(new_n361), .ZN(G3));
  NAND2_X1  g373(.A1(new_n302), .A2(new_n187), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G472), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n308), .A2(new_n561), .A3(new_n309), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n471), .A2(new_n555), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n538), .A2(new_n539), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT33), .B1(new_n538), .B2(new_n539), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G478), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n541), .A2(new_n187), .ZN(new_n571));
  INV_X1    g385(.A(new_n540), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(new_n541), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n512), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n563), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n562), .A2(new_n350), .A3(new_n424), .A4(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G104), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G6));
  INV_X1    g393(.A(new_n512), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n546), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n563), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n562), .A2(new_n350), .A3(new_n424), .A4(new_n582), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G107), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G9));
  INV_X1    g399(.A(new_n336), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n342), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n586), .B(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n589), .A2(G902), .A3(new_n347), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n348), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n556), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n562), .A2(new_n472), .A3(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT37), .B(G110), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G12));
  NAND2_X1  g409(.A1(new_n312), .A2(new_n314), .ZN(new_n596));
  INV_X1    g410(.A(new_n305), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n424), .A2(new_n591), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n554), .A2(G900), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n550), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n581), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n471), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n598), .A2(KEYINPUT96), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n315), .B2(new_n604), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G128), .ZN(G30));
  XNOR2_X1  g424(.A(new_n601), .B(KEYINPUT39), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n424), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT40), .Z(new_n613));
  NAND2_X1  g427(.A1(new_n263), .A2(new_n292), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n291), .B2(new_n292), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n615), .B2(KEYINPUT97), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(KEYINPUT97), .B2(new_n615), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(G472), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n304), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n302), .A2(KEYINPUT73), .A3(new_n303), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT73), .B1(new_n302), .B2(new_n303), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n313), .B1(new_n623), .B2(new_n310), .ZN(new_n624));
  INV_X1    g438(.A(new_n314), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n620), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n469), .A2(new_n470), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT38), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n512), .A2(new_n546), .ZN(new_n630));
  NOR4_X1   g444(.A1(new_n629), .A2(new_n426), .A3(new_n591), .A4(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n613), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT98), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G143), .ZN(G45));
  NOR2_X1   g448(.A1(new_n574), .A2(new_n602), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n599), .A2(new_n471), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n315), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(new_n226), .ZN(G48));
  NOR2_X1   g452(.A1(new_n401), .A2(new_n408), .ZN(new_n639));
  OAI21_X1  g453(.A(G469), .B1(new_n639), .B2(G902), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(new_n423), .A3(new_n409), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT99), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n598), .A2(new_n350), .A3(new_n575), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT41), .B(G113), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G15));
  NAND4_X1  g463(.A1(new_n598), .A2(new_n350), .A3(new_n582), .A4(new_n646), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G116), .ZN(G18));
  INV_X1    g465(.A(new_n592), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n596), .B2(new_n597), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n471), .A2(new_n640), .A3(new_n423), .A4(new_n409), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT100), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G119), .ZN(G21));
  INV_X1    g472(.A(new_n563), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n630), .B(KEYINPUT102), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n643), .A2(new_n659), .A3(new_n645), .A4(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n264), .A2(new_n292), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n297), .B(KEYINPUT31), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n303), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n561), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT101), .B1(new_n560), .B2(G472), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n350), .B(new_n664), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n669), .B(G122), .Z(G24));
  OAI211_X1 g484(.A(new_n591), .B(new_n664), .C1(new_n666), .C2(new_n667), .ZN(new_n671));
  INV_X1    g485(.A(new_n635), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n655), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(G125), .Z(G27));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n418), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n402), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n395), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n678), .A2(KEYINPUT103), .A3(G469), .A4(new_n413), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n409), .A2(new_n676), .A3(new_n420), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(KEYINPUT104), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n680), .A2(KEYINPUT104), .ZN(new_n683));
  OAI211_X1 g497(.A(KEYINPUT105), .B(new_n423), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n627), .A2(new_n426), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n423), .ZN(new_n687));
  INV_X1    g501(.A(new_n400), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n412), .B1(new_n417), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n677), .A2(new_n410), .ZN(new_n690));
  AOI21_X1  g504(.A(G902), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n419), .B1(new_n691), .B2(new_n353), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n676), .A2(new_n679), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n687), .B1(new_n695), .B2(new_n681), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(KEYINPUT105), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n686), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  INV_X1    g513(.A(new_n304), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT32), .B1(new_n302), .B2(new_n303), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT32), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n306), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(KEYINPUT106), .A3(new_n304), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n705), .A3(new_n295), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n706), .A2(new_n707), .A3(new_n350), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n707), .B1(new_n706), .B2(new_n350), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n698), .B(new_n635), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n696), .A2(KEYINPUT105), .ZN(new_n711));
  INV_X1    g525(.A(new_n685), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n712), .B1(new_n696), .B2(KEYINPUT105), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n714), .A2(new_n315), .A3(new_n351), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n672), .A2(KEYINPUT42), .ZN(new_n716));
  AOI22_X1  g530(.A1(KEYINPUT42), .A2(new_n710), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G131), .ZN(G33));
  NAND3_X1  g532(.A1(new_n352), .A2(new_n603), .A3(new_n698), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G134), .ZN(G36));
  OAI21_X1  g534(.A(new_n413), .B1(new_n417), .B2(new_n402), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n353), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n722), .B2(new_n721), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n724), .A2(new_n420), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT46), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n726), .B(KEYINPUT108), .Z(new_n727));
  NOR2_X1   g541(.A1(new_n725), .A2(KEYINPUT46), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n353), .B2(new_n691), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n730), .A2(new_n423), .A3(new_n611), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n512), .B(KEYINPUT109), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n573), .B1(new_n568), .B2(new_n541), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n734), .A3(KEYINPUT43), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n735), .A2(KEYINPUT110), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(KEYINPUT110), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n733), .A2(new_n512), .ZN(new_n738));
  OAI22_X1  g552(.A1(new_n736), .A2(new_n737), .B1(KEYINPUT43), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n562), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n591), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n712), .B1(new_n741), .B2(new_n742), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n731), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G137), .ZN(G39));
  NOR4_X1   g560(.A1(new_n598), .A2(new_n350), .A3(new_n672), .A4(new_n712), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT47), .B1(new_n730), .B2(new_n423), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n749));
  AOI211_X1 g563(.A(new_n749), .B(new_n687), .C1(new_n727), .C2(new_n729), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n747), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G140), .ZN(G42));
  NOR3_X1   g566(.A1(new_n351), .A2(new_n687), .A3(new_n426), .ZN(new_n753));
  AND4_X1   g567(.A1(new_n734), .A2(new_n753), .A3(new_n629), .A4(new_n732), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n619), .B1(new_n312), .B2(new_n314), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n640), .A2(new_n409), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n754), .A2(new_n755), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n673), .B1(new_n606), .B2(new_n608), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n695), .A2(new_n681), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n348), .A2(new_n687), .A3(new_n590), .A4(new_n602), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n764), .A2(new_n660), .A3(new_n471), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n626), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT113), .B1(new_n755), .B2(new_n766), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n637), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n762), .A2(new_n770), .A3(KEYINPUT114), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT114), .B1(new_n762), .B2(new_n770), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n761), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT96), .B1(new_n598), .B2(new_n605), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n315), .A2(new_n607), .A3(new_n604), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n561), .B(new_n665), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n591), .A3(new_n635), .A4(new_n664), .ZN(new_n778));
  OAI22_X1  g592(.A1(new_n775), .A2(new_n776), .B1(new_n655), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n637), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n763), .B1(new_n626), .B2(new_n767), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n755), .A2(KEYINPUT113), .A3(new_n766), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n774), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n762), .A2(new_n770), .A3(KEYINPUT114), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(KEYINPUT52), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n710), .A2(KEYINPUT42), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n715), .A2(new_n716), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n576), .A2(new_n583), .A3(new_n593), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n352), .B2(new_n557), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n669), .B1(new_n653), .B2(new_n656), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n792), .A3(new_n647), .A4(new_n650), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n580), .A2(new_n543), .A3(new_n545), .A4(new_n601), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT111), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n547), .A2(new_n796), .A3(new_n601), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n797), .A3(new_n685), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n795), .A2(new_n797), .A3(KEYINPUT112), .A4(new_n685), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n599), .A3(new_n801), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(new_n315), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n719), .B(new_n803), .C1(new_n778), .C2(new_n714), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n789), .A2(new_n793), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n773), .A2(new_n786), .A3(new_n805), .A4(KEYINPUT53), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n761), .B1(new_n762), .B2(new_n770), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n784), .A2(new_n785), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(new_n761), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n805), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n806), .A2(new_n807), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n808), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT54), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n773), .A2(new_n786), .A3(new_n805), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n813), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n792), .A2(new_n647), .A3(new_n650), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n791), .A2(KEYINPUT53), .ZN(new_n823));
  OAI22_X1  g637(.A1(new_n714), .A2(new_n778), .B1(new_n802), .B2(new_n315), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n603), .B2(new_n715), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n717), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n811), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n819), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n817), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n739), .A2(new_n549), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n668), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n426), .A3(new_n629), .A4(new_n642), .ZN(new_n834));
  XOR2_X1   g648(.A(new_n834), .B(KEYINPUT50), .Z(new_n835));
  NOR2_X1   g649(.A1(new_n712), .A2(new_n641), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n626), .A2(new_n837), .A3(new_n351), .A4(new_n550), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n580), .A3(new_n733), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n832), .A2(new_n837), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n835), .B(new_n839), .C1(new_n671), .C2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n833), .A2(new_n685), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n748), .A2(new_n750), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n756), .A2(new_n687), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n842), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n843), .B1(new_n842), .B2(new_n847), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n708), .A2(new_n709), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n840), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT48), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(KEYINPUT117), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n833), .A2(new_n656), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n838), .A2(new_n512), .A3(new_n734), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n854), .A2(new_n855), .A3(G952), .A4(new_n338), .ZN(new_n856));
  INV_X1    g670(.A(new_n851), .ZN(new_n857));
  XNOR2_X1  g671(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n848), .A2(new_n849), .A3(new_n853), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n831), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(G952), .A2(G953), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n760), .B1(new_n861), .B2(new_n862), .ZN(G75));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n187), .B1(new_n819), .B2(new_n828), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n864), .B1(new_n866), .B2(new_n265), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n445), .A2(new_n447), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT118), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n453), .B(KEYINPUT55), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n869), .B(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n867), .A2(new_n871), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n338), .A2(G952), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G51));
  AND3_X1   g689(.A1(new_n792), .A2(new_n647), .A3(new_n650), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n717), .A2(new_n876), .A3(new_n825), .A4(new_n791), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n810), .B2(new_n761), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT53), .B1(new_n878), .B2(new_n786), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT52), .B1(new_n784), .B2(new_n785), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n880), .A2(new_n822), .A3(new_n809), .A4(new_n826), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT54), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n830), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n419), .B(KEYINPUT57), .Z(new_n885));
  OAI22_X1  g699(.A1(new_n884), .A2(new_n885), .B1(new_n401), .B2(new_n408), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n724), .B(KEYINPUT119), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n865), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n874), .B1(new_n886), .B2(new_n888), .ZN(G54));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n890));
  INV_X1    g704(.A(new_n874), .ZN(new_n891));
  AND2_X1   g705(.A1(KEYINPUT58), .A2(G475), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n865), .A2(new_n506), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n506), .B1(new_n865), .B2(new_n892), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n891), .B(new_n893), .C1(new_n894), .C2(KEYINPUT120), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n819), .A2(new_n828), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n896), .A2(G902), .A3(new_n892), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT120), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n506), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n890), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n898), .B1(new_n897), .B2(new_n506), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n874), .B1(new_n897), .B2(new_n506), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n894), .A2(KEYINPUT120), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT121), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n900), .A2(new_n904), .ZN(G60));
  XNOR2_X1  g719(.A(new_n571), .B(KEYINPUT59), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n569), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT122), .B1(new_n883), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n909));
  INV_X1    g723(.A(new_n907), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n909), .B(new_n910), .C1(new_n882), .C2(new_n830), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n891), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n906), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n568), .B1(new_n831), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(G63));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n813), .A2(new_n818), .B1(new_n811), .B2(new_n827), .ZN(new_n917));
  XNOR2_X1  g731(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n346), .A2(new_n187), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT124), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n896), .A2(new_n923), .A3(new_n920), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n924), .A3(new_n343), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n891), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n589), .B1(new_n922), .B2(new_n924), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n916), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n922), .A2(new_n924), .ZN(new_n929));
  INV_X1    g743(.A(new_n589), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n931), .A2(KEYINPUT61), .A3(new_n891), .A4(new_n925), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n932), .ZN(G66));
  INV_X1    g747(.A(new_n552), .ZN(new_n934));
  OAI21_X1  g748(.A(G953), .B1(new_n934), .B2(new_n451), .ZN(new_n935));
  INV_X1    g749(.A(new_n793), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(G953), .ZN(new_n937));
  INV_X1    g751(.A(new_n869), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(G898), .B2(new_n338), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n937), .B(new_n939), .ZN(G69));
  AOI21_X1  g754(.A(new_n338), .B1(G227), .B2(G900), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n731), .A2(new_n471), .A3(new_n660), .A4(new_n850), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(new_n751), .A3(new_n745), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n762), .A2(new_n780), .A3(new_n719), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n943), .A2(new_n789), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(G953), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n338), .A2(G900), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n946), .A2(KEYINPUT126), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n262), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n288), .B1(new_n950), .B2(new_n285), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(new_n502), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT126), .B1(new_n946), .B2(new_n947), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n949), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI211_X1 g769(.A(new_n712), .B(new_n612), .C1(new_n574), .C2(new_n581), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n352), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n745), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT125), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n633), .A2(new_n780), .A3(new_n762), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n959), .A2(new_n751), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n338), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n952), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n941), .B1(new_n955), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n954), .A2(new_n953), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n965), .B(new_n941), .C1(new_n967), .C2(new_n948), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n966), .A2(new_n969), .ZN(G72));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n963), .B2(new_n793), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n291), .A2(new_n292), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n972), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n945), .B2(new_n936), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n975), .B(new_n891), .C1(new_n293), .C2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n293), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n979), .A2(new_n974), .A3(new_n976), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n978), .B1(new_n816), .B2(new_n980), .ZN(G57));
endmodule


