//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203));
  AND2_X1   g002(.A1(G113gat), .A2(G120gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G113gat), .A2(G120gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G113gat), .A2(G120gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(KEYINPUT70), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212));
  XNOR2_X1  g011(.A(G127gat), .B(G134gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n206), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT69), .B1(new_n204), .B2(new_n205), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT69), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n209), .A2(new_n216), .A3(new_n210), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n215), .A2(new_n217), .A3(new_n212), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(KEYINPUT68), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n220));
  INV_X1    g019(.A(G127gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G134gat), .ZN(new_n222));
  INV_X1    g021(.A(G134gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G127gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n220), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n214), .B1(new_n218), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT24), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n231), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G169gat), .ZN(new_n239));
  INV_X1    g038(.A(G176gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(KEYINPUT65), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244));
  NOR2_X1   g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(KEYINPUT23), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n241), .B2(new_n242), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n238), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n246), .B2(new_n243), .ZN(new_n253));
  INV_X1    g052(.A(new_n235), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n233), .B2(new_n254), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n251), .A2(new_n252), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT26), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n257), .A3(new_n248), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n245), .A2(KEYINPUT26), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n259), .A3(new_n229), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT27), .B(G183gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(G190gat), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT67), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT27), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G183gat), .ZN(new_n266));
  INV_X1    g065(.A(G183gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT27), .ZN(new_n268));
  AND4_X1   g067(.A1(KEYINPUT67), .A2(new_n263), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G183gat), .ZN(new_n272));
  AOI21_X1  g071(.A(G190gat), .B1(new_n272), .B2(KEYINPUT27), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n265), .A3(G183gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n262), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n260), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n228), .B1(new_n256), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n260), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n266), .A3(new_n268), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n261), .A2(KEYINPUT67), .A3(new_n263), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT28), .B1(new_n273), .B2(new_n274), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n279), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT25), .B1(new_n253), .B2(new_n238), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n255), .A2(new_n247), .A3(new_n250), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n286), .B(new_n227), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n278), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G227gat), .A2(G233gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n202), .B1(new_n292), .B2(KEYINPUT34), .ZN(new_n293));
  INV_X1    g092(.A(new_n291), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n294), .B1(new_n278), .B2(new_n289), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT34), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(KEYINPUT72), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n292), .A2(new_n299), .A3(KEYINPUT34), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT71), .B1(new_n295), .B2(new_n296), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n278), .A2(new_n294), .A3(new_n289), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT32), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT33), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G15gat), .B(G43gat), .Z(new_n307));
  XNOR2_X1  g106(.A(G71gat), .B(G99gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n309), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n303), .B(KEYINPUT32), .C1(new_n305), .C2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n298), .A2(new_n302), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n299), .B1(new_n292), .B2(KEYINPUT34), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n295), .A2(KEYINPUT71), .A3(new_n296), .ZN(new_n315));
  AND4_X1   g114(.A1(KEYINPUT72), .A2(new_n290), .A3(new_n296), .A4(new_n291), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT72), .B1(new_n295), .B2(new_n296), .ZN(new_n317));
  OAI22_X1  g116(.A1(new_n314), .A2(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n310), .A2(new_n312), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G141gat), .ZN(new_n321));
  INV_X1    g120(.A(G148gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324));
  AND2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(KEYINPUT75), .A3(new_n324), .ZN(new_n328));
  NOR2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT2), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G155gat), .B(G162gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n334), .B(new_n337), .C1(new_n338), .C2(KEYINPUT75), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(G211gat), .A2(G218gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(G211gat), .A2(G218gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(G197gat), .A2(G204gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G211gat), .B(G218gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G197gat), .B(G204gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n347), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT29), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n340), .B1(new_n353), .B2(KEYINPUT3), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT78), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n356), .B(new_n340), .C1(new_n353), .C2(KEYINPUT3), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n331), .A2(new_n358), .A3(new_n339), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n348), .A2(new_n352), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n355), .A2(new_n357), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n358), .B1(new_n353), .B2(KEYINPUT79), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n369));
  AOI211_X1 g168(.A(new_n369), .B(KEYINPUT29), .C1(new_n348), .C2(new_n352), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n340), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n366), .B1(new_n361), .B2(new_n363), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n371), .B2(new_n373), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n367), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G22gat), .ZN(new_n377));
  INV_X1    g176(.A(G22gat), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n378), .B(new_n367), .C1(new_n374), .C2(new_n375), .ZN(new_n379));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT31), .B(G50gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n377), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n382), .B1(new_n377), .B2(new_n379), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n313), .B(new_n320), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G226gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(new_n360), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n251), .A2(new_n252), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n253), .A2(new_n255), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n386), .B1(new_n392), .B2(new_n286), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n363), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n387), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n392), .B2(new_n286), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n362), .B(new_n395), .C1(new_n396), .C2(new_n387), .ZN(new_n397));
  XOR2_X1   g196(.A(G8gat), .B(G36gat), .Z(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(KEYINPUT74), .ZN(new_n399));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n394), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n394), .A2(new_n397), .A3(KEYINPUT30), .A4(new_n401), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n394), .A2(new_n397), .ZN(new_n406));
  INV_X1    g205(.A(new_n401), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n385), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT87), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT35), .ZN(new_n412));
  XOR2_X1   g211(.A(G1gat), .B(G29gat), .Z(new_n413));
  XNOR2_X1  g212(.A(G57gat), .B(G85gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n331), .A2(new_n339), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n215), .A2(new_n217), .A3(new_n212), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n225), .A3(new_n219), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n214), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n227), .A2(new_n340), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G225gat), .A2(G233gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n418), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(new_n227), .B2(new_n340), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n340), .A2(KEYINPUT3), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n227), .A3(new_n359), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n419), .A2(KEYINPUT4), .A3(new_n214), .A4(new_n421), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n429), .A2(new_n431), .A3(new_n425), .A4(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n417), .B1(new_n427), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT77), .ZN(new_n435));
  AND4_X1   g234(.A1(new_n425), .A2(new_n429), .A3(new_n431), .A4(new_n432), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(new_n418), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n433), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n417), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(new_n435), .A3(new_n418), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT77), .B1(new_n433), .B2(KEYINPUT5), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n433), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT83), .B1(new_n441), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(KEYINPUT6), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n446), .B1(new_n437), .B2(new_n438), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n417), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT6), .B1(new_n445), .B2(new_n434), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n448), .A2(new_n449), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n410), .A2(new_n411), .A3(new_n412), .A4(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n318), .A2(new_n319), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n298), .A2(new_n302), .B1(new_n310), .B2(new_n312), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n382), .ZN(new_n460));
  INV_X1    g259(.A(new_n375), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n378), .B1(new_n463), .B2(new_n367), .ZN(new_n464));
  INV_X1    g263(.A(new_n379), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n377), .A2(new_n379), .A3(new_n382), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n409), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n459), .A2(new_n412), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n448), .A2(new_n449), .A3(new_n454), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT87), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n451), .A2(new_n453), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n449), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n469), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n385), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n459), .A2(KEYINPUT88), .A3(new_n468), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n456), .B(new_n472), .C1(new_n479), .C2(new_n412), .ZN(new_n480));
  INV_X1    g279(.A(new_n468), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n426), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n483), .A2(KEYINPUT39), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT39), .B1(new_n424), .B2(new_n426), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n485), .A2(KEYINPUT81), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n483), .B1(new_n485), .B2(KEYINPUT81), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n484), .B(new_n442), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT82), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(KEYINPUT40), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n487), .A2(new_n486), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n489), .A2(KEYINPUT40), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n491), .A2(new_n484), .A3(new_n442), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n447), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n481), .B1(new_n494), .B2(new_n409), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT84), .B(KEYINPUT37), .Z(new_n497));
  NAND3_X1  g296(.A1(new_n394), .A2(new_n397), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT85), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n394), .A2(new_n397), .A3(new_n500), .A4(new_n497), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n401), .B1(new_n406), .B2(KEYINPUT37), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n496), .B1(new_n504), .B2(KEYINPUT38), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(KEYINPUT38), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT38), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n502), .A2(KEYINPUT86), .A3(new_n507), .A4(new_n503), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n505), .A2(new_n506), .A3(new_n508), .A4(new_n402), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n495), .B1(new_n509), .B2(new_n455), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n511), .A2(KEYINPUT73), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(KEYINPUT73), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n459), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n320), .A2(new_n313), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(KEYINPUT73), .B2(new_n511), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n514), .A2(new_n516), .B1(new_n475), .B2(new_n481), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n480), .A2(KEYINPUT89), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT89), .B1(new_n480), .B2(new_n518), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G43gat), .B(G50gat), .Z(new_n522));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n522), .A2(new_n523), .B1(G29gat), .B2(G36gat), .ZN(new_n524));
  OR3_X1    g323(.A1(KEYINPUT92), .A2(G29gat), .A3(G36gat), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT92), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(KEYINPUT14), .A3(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n526), .A2(KEYINPUT14), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n522), .A2(new_n523), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n530), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(new_n524), .A3(new_n527), .A4(new_n528), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OR3_X1    g337(.A1(new_n534), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT17), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G85gat), .A2(G92gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544));
  INV_X1    g343(.A(G85gat), .ZN(new_n545));
  INV_X1    g344(.A(G92gat), .ZN(new_n546));
  AOI22_X1  g345(.A1(KEYINPUT8), .A2(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G99gat), .B(G106gat), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n548), .B(new_n549), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n541), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT100), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT101), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT99), .Z(new_n558));
  INV_X1    g357(.A(KEYINPUT41), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n548), .B(new_n549), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n560), .B1(new_n534), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n553), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n556), .B1(new_n553), .B2(new_n562), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n558), .A2(new_n559), .ZN(new_n565));
  XNOR2_X1  g364(.A(G134gat), .B(G162gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  OR3_X1    g367(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n563), .B2(new_n564), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT104), .ZN(new_n573));
  XOR2_X1   g372(.A(G176gat), .B(G204gat), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G57gat), .B(G64gat), .Z(new_n578));
  INV_X1    g377(.A(KEYINPUT9), .ZN(new_n579));
  INV_X1    g378(.A(G71gat), .ZN(new_n580));
  INV_X1    g379(.A(G78gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(KEYINPUT97), .A3(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G71gat), .B(G78gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n550), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n583), .B(new_n584), .Z(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n561), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT10), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n561), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n577), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n576), .B1(new_n586), .B2(new_n588), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n575), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT105), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT106), .ZN(new_n597));
  INV_X1    g396(.A(new_n593), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n598), .A2(KEYINPUT103), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(KEYINPUT103), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n599), .A2(new_n600), .A3(new_n575), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n590), .A2(new_n591), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n577), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n590), .A2(KEYINPUT102), .A3(new_n591), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n596), .A2(new_n597), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n597), .B1(new_n596), .B2(new_n607), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT21), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n585), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G127gat), .ZN(new_n616));
  INV_X1    g415(.A(G8gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G15gat), .B(G22gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT16), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n618), .B1(new_n619), .B2(G1gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT93), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(G1gat), .B2(new_n618), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n612), .B2(new_n585), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n616), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G183gat), .B(G211gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT98), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n335), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n631), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n629), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n571), .A2(new_n611), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G113gat), .B(G141gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G169gat), .B(G197gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT12), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n626), .A2(new_n534), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n541), .B2(new_n627), .ZN(new_n648));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n648), .B(new_n649), .C1(KEYINPUT95), .C2(KEYINPUT18), .ZN(new_n650));
  INV_X1    g449(.A(new_n540), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n534), .A2(new_n536), .A3(new_n538), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n627), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(new_n649), .A3(new_n646), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT95), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT18), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OR3_X1    g456(.A1(new_n626), .A2(new_n534), .A3(KEYINPUT96), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT96), .B1(new_n626), .B2(new_n534), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n658), .A2(new_n646), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n649), .B(KEYINPUT13), .Z(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n650), .A2(new_n657), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT91), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n645), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n645), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n664), .A2(KEYINPUT91), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n639), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n521), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n474), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n409), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G8gat), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  NAND4_X1  g480(.A1(new_n673), .A2(KEYINPUT42), .A3(new_n409), .A4(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n681), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n680), .B(new_n682), .C1(new_n684), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g484(.A(new_n673), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n514), .A2(new_n516), .ZN(new_n687));
  OAI21_X1  g486(.A(G15gat), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n515), .A2(G15gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n686), .B2(new_n689), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n481), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT108), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT43), .B(G22gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(new_n638), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n611), .A2(new_n695), .A3(new_n670), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n571), .B(new_n696), .C1(new_n519), .C2(new_n520), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n697), .A2(G29gat), .A3(new_n474), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT45), .Z(new_n699));
  INV_X1    g498(.A(new_n696), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n571), .B1(new_n519), .B2(new_n520), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT44), .ZN(new_n702));
  INV_X1    g501(.A(new_n571), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n703), .B1(new_n480), .B2(new_n518), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n700), .B1(new_n702), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n474), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n699), .A2(new_n709), .ZN(G1328gat));
  OAI21_X1  g509(.A(G36gat), .B1(new_n708), .B2(new_n469), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n697), .A2(G36gat), .A3(new_n469), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT46), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(G1329gat));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n708), .A2(new_n687), .ZN(new_n716));
  INV_X1    g515(.A(G43gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OR3_X1    g517(.A1(new_n697), .A2(G43gat), .A3(new_n515), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n716), .B2(new_n717), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  OAI221_X1 g521(.A(new_n719), .B1(new_n715), .B2(KEYINPUT47), .C1(new_n716), .C2(new_n717), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1330gat));
  INV_X1    g523(.A(G50gat), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n707), .B2(new_n481), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n521), .A2(KEYINPUT111), .A3(new_n571), .A4(new_n696), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n697), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n468), .A2(G50gat), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT112), .B1(new_n726), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT48), .B1(new_n733), .B2(KEYINPUT110), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735));
  INV_X1    g534(.A(new_n706), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n701), .B2(KEYINPUT44), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(new_n468), .A3(new_n700), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n735), .B(new_n733), .C1(new_n738), .C2(new_n725), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n732), .A2(new_n734), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n734), .B1(new_n732), .B2(new_n739), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(G1331gat));
  NAND4_X1  g541(.A1(new_n703), .A2(new_n670), .A3(new_n695), .A4(new_n611), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(new_n518), .B2(new_n480), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n674), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n409), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT49), .B(G64gat), .Z(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1333gat));
  INV_X1    g549(.A(new_n687), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n580), .B1(new_n744), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n515), .A2(G71gat), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n744), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n744), .A2(new_n481), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT113), .B(G78gat), .Z(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1335gat));
  NOR2_X1   g557(.A1(new_n671), .A2(new_n695), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n611), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n737), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G85gat), .B1(new_n762), .B2(new_n474), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n704), .A2(new_n759), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT51), .Z(new_n765));
  NAND4_X1  g564(.A1(new_n765), .A2(new_n545), .A3(new_n674), .A4(new_n611), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(G1336gat));
  OAI21_X1  g566(.A(G92gat), .B1(new_n762), .B2(new_n469), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n611), .A2(new_n546), .A3(new_n409), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT114), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT52), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n768), .A2(new_n774), .A3(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1337gat));
  OAI21_X1  g575(.A(G99gat), .B1(new_n762), .B2(new_n687), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n610), .A2(G99gat), .A3(new_n515), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT115), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n765), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(G1338gat));
  INV_X1    g580(.A(G106gat), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n765), .A2(new_n782), .A3(new_n481), .A4(new_n611), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n737), .A2(new_n468), .A3(new_n760), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n782), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n784), .B2(new_n782), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(KEYINPUT53), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789));
  OAI221_X1 g588(.A(new_n783), .B1(new_n786), .B2(new_n789), .C1(new_n784), .C2(new_n782), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1339gat));
  OAI21_X1  g590(.A(KEYINPUT117), .B1(new_n648), .B2(new_n649), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n660), .A2(new_n662), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n648), .A2(KEYINPUT117), .A3(new_n649), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n644), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n665), .A2(new_n668), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n796), .B(new_n797), .C1(new_n608), .C2(new_n609), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT54), .B1(new_n602), .B2(new_n576), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n605), .B2(new_n604), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n602), .A2(new_n576), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n575), .B1(new_n801), .B2(KEYINPUT54), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n803), .A2(KEYINPUT55), .B1(new_n606), .B2(new_n601), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n800), .B2(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n798), .A2(KEYINPUT118), .B1(new_n670), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n798), .A2(KEYINPUT118), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n703), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n797), .A2(new_n796), .ZN(new_n811));
  INV_X1    g610(.A(new_n807), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n571), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n695), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  NOR4_X1   g613(.A1(new_n571), .A2(new_n671), .A3(new_n611), .A4(new_n638), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n674), .A3(new_n410), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT119), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n816), .A2(new_n819), .A3(new_n674), .A4(new_n410), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n821), .A2(new_n207), .A3(new_n670), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n816), .A2(new_n674), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n477), .A2(new_n478), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n409), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n671), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n822), .A2(new_n828), .ZN(G1340gat));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n208), .A3(new_n611), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n818), .A2(new_n611), .A3(new_n820), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n831), .A2(KEYINPUT120), .A3(G120gat), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT120), .B1(new_n831), .B2(G120gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(G1341gat));
  OAI21_X1  g633(.A(G127gat), .B1(new_n821), .B2(new_n638), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n827), .A2(new_n221), .A3(new_n695), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1342gat));
  NAND4_X1  g636(.A1(new_n823), .A2(new_n223), .A3(new_n571), .A4(new_n825), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n838), .A2(KEYINPUT56), .ZN(new_n839));
  OAI21_X1  g638(.A(G134gat), .B1(new_n821), .B2(new_n703), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(KEYINPUT56), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(G1343gat));
  NAND2_X1  g641(.A1(new_n687), .A2(new_n481), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n409), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n823), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n321), .B1(new_n845), .B2(new_n670), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n751), .A2(new_n474), .A3(new_n409), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n804), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n806), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n806), .A2(new_n850), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n671), .A2(new_n853), .B1(new_n611), .B2(new_n811), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n813), .B1(new_n854), .B2(new_n571), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n815), .B1(new_n855), .B2(new_n638), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n856), .A2(new_n857), .A3(new_n468), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n848), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n670), .A2(new_n321), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n816), .B2(new_n481), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n855), .A2(new_n638), .ZN(new_n863));
  INV_X1    g662(.A(new_n815), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(KEYINPUT57), .A3(new_n481), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT122), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n860), .B(new_n861), .C1(new_n862), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n846), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n846), .A2(KEYINPUT58), .A3(new_n868), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1344gat));
  INV_X1    g672(.A(new_n845), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n322), .A3(new_n611), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G148gat), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n867), .A2(new_n862), .ZN(new_n878));
  INV_X1    g677(.A(new_n860), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n877), .B1(new_n880), .B2(new_n611), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n857), .B1(new_n856), .B2(new_n468), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT57), .B(new_n481), .C1(new_n814), .C2(new_n815), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n611), .A3(new_n847), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n876), .B1(new_n885), .B2(G148gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n875), .B1(new_n881), .B2(new_n886), .ZN(G1345gat));
  AOI21_X1  g686(.A(G155gat), .B1(new_n874), .B2(new_n695), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n638), .A2(new_n335), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT123), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n888), .B1(new_n880), .B2(new_n890), .ZN(G1346gat));
  AOI21_X1  g690(.A(G162gat), .B1(new_n874), .B2(new_n571), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n703), .A2(new_n336), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n880), .B2(new_n893), .ZN(G1347gat));
  AND2_X1   g693(.A1(new_n816), .A2(new_n474), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n824), .A2(new_n469), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n239), .B1(new_n897), .B2(new_n670), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n385), .A2(new_n469), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n895), .A2(G169gat), .A3(new_n671), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n898), .A2(KEYINPUT124), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1348gat));
  NAND3_X1  g704(.A1(new_n895), .A2(new_n611), .A3(new_n899), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G176gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n611), .A2(new_n240), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n897), .B2(new_n908), .ZN(G1349gat));
  NAND4_X1  g708(.A1(new_n816), .A2(new_n474), .A3(new_n695), .A4(new_n899), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G183gat), .ZN(new_n911));
  NAND2_X1  g710(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n695), .A2(new_n261), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n911), .B(new_n912), .C1(new_n897), .C2(new_n913), .ZN(new_n914));
  OR2_X1    g713(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n895), .A2(new_n571), .A3(new_n899), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G190gat), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(KEYINPUT61), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(KEYINPUT61), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n703), .A2(G190gat), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n919), .A2(new_n920), .B1(new_n897), .B2(new_n921), .ZN(G1351gat));
  NOR2_X1   g721(.A1(new_n843), .A2(new_n469), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n895), .A2(new_n923), .ZN(new_n924));
  OR3_X1    g723(.A1(new_n924), .A2(G197gat), .A3(new_n670), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n751), .A2(new_n674), .A3(new_n469), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n927), .B1(new_n882), .B2(new_n883), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n929), .A2(new_n670), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(KEYINPUT126), .ZN(new_n931));
  OAI21_X1  g730(.A(G197gat), .B1(new_n930), .B2(KEYINPUT126), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n925), .B1(new_n931), .B2(new_n932), .ZN(G1352gat));
  OR2_X1    g732(.A1(new_n610), .A2(G204gat), .ZN(new_n934));
  OR3_X1    g733(.A1(new_n924), .A2(KEYINPUT62), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G204gat), .B1(new_n929), .B2(new_n610), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT62), .B1(new_n924), .B2(new_n934), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(G1353gat));
  INV_X1    g737(.A(G211gat), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n895), .A2(new_n939), .A3(new_n695), .A4(new_n923), .ZN(new_n940));
  AOI211_X1 g739(.A(new_n638), .B(new_n927), .C1(new_n882), .C2(new_n883), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n928), .B2(new_n695), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT63), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n884), .A2(new_n942), .A3(new_n695), .A4(new_n926), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G211gat), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n948), .A2(new_n944), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n940), .B1(new_n946), .B2(new_n950), .ZN(G1354gat));
  OAI21_X1  g750(.A(G218gat), .B1(new_n929), .B2(new_n703), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n703), .A2(G218gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n924), .B2(new_n953), .ZN(G1355gat));
endmodule


