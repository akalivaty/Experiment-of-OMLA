//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G219), .A2(G218), .A3(G221), .A4(G220), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND3_X1  g030(.A1(new_n455), .A2(KEYINPUT68), .A3(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  AOI21_X1  g033(.A(KEYINPUT68), .B1(new_n455), .B2(G2106), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n473), .A2(G137), .A3(new_n474), .A4(new_n463), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n470), .B2(new_n472), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n469), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n473), .A2(new_n463), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n474), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n474), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n482), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT70), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(new_n474), .A3(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n466), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n474), .A2(G138), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n473), .A2(new_n463), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n491), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n473), .A2(G126), .A3(G2105), .A4(new_n463), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT71), .B(G114), .ZN(new_n497));
  OAI211_X1 g072(.A(G2104), .B(new_n496), .C1(new_n497), .C2(new_n474), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT72), .B1(new_n502), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n502), .A2(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n507), .A2(G88), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(G50), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n510), .A2(KEYINPUT73), .A3(new_n511), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n504), .B1(KEYINPUT5), .B2(new_n505), .ZN(new_n516));
  NOR3_X1   g091(.A1(new_n502), .A2(KEYINPUT72), .A3(G543), .ZN(new_n517));
  OAI211_X1 g092(.A(G62), .B(new_n508), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n507), .A2(KEYINPUT74), .A3(G62), .A4(new_n508), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n514), .A2(new_n515), .B1(new_n523), .B2(G651), .ZN(G166));
  AND2_X1   g099(.A1(new_n507), .A2(new_n508), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n509), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(new_n509), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n526), .B(new_n529), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT75), .ZN(new_n534));
  XOR2_X1   g109(.A(new_n534), .B(KEYINPUT7), .Z(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n528), .A2(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n530), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n538), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  XOR2_X1   g121(.A(KEYINPUT76), .B(G43), .Z(new_n547));
  OAI22_X1  g122(.A1(new_n530), .A2(new_n546), .B1(new_n527), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT77), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n551), .B1(new_n545), .B2(new_n548), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT78), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(KEYINPUT79), .B2(KEYINPUT9), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n528), .B(new_n561), .C1(KEYINPUT79), .C2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n563), .B(new_n564), .C1(new_n527), .C2(new_n560), .ZN(new_n565));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n562), .B(new_n565), .C1(new_n530), .C2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n525), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n538), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  NAND2_X1  g148(.A1(new_n514), .A2(new_n515), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n523), .A2(G651), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G303));
  AND2_X1   g151(.A1(new_n525), .A2(new_n509), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G87), .B1(G49), .B2(new_n528), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G288));
  NAND3_X1  g155(.A1(new_n525), .A2(G86), .A3(new_n509), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n528), .A2(G48), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g158(.A1(new_n507), .A2(G61), .A3(new_n508), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n538), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n528), .A2(G47), .ZN(new_n591));
  XNOR2_X1  g166(.A(KEYINPUT80), .B(G85), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n530), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n577), .A2(new_n597), .A3(G92), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT81), .B1(new_n530), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n598), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT10), .B1(new_n598), .B2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n528), .A2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n525), .A2(G66), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n603), .B1(new_n606), .B2(new_n538), .ZN(new_n607));
  NOR3_X1   g182(.A1(new_n601), .A2(new_n602), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n596), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n596), .B1(new_n608), .B2(G868), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n570), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(new_n570), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n608), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n608), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g194(.A1(new_n463), .A2(new_n465), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n476), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT83), .B(G2100), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT84), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n481), .A2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n483), .A2(G123), .ZN(new_n630));
  OR2_X1    g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n631), .B(G2104), .C1(G111), .C2(new_n474), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n624), .A2(new_n626), .ZN(new_n636));
  NAND4_X1  g211(.A1(new_n628), .A2(new_n634), .A3(new_n635), .A4(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT85), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT86), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n655), .A2(new_n656), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n663), .B(new_n667), .Z(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n673), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  AOI211_X1 g252(.A(new_n675), .B(new_n677), .C1(new_n670), .C2(new_n674), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G229));
  NAND3_X1  g259(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT25), .Z(new_n686));
  AOI22_X1  g261(.A1(new_n620), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n474), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G139), .B2(new_n481), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n690), .B2(G33), .ZN(new_n692));
  INV_X1    g267(.A(G2072), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT87), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G34), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(new_n690), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n478), .B2(new_n690), .ZN(new_n699));
  INV_X1    g274(.A(G2084), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n481), .A2(G141), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n483), .A2(G129), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT26), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  AOI22_X1  g282(.A1(G105), .A2(new_n476), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n702), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G29), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT89), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n710), .B(new_n711), .C1(G29), .C2(G32), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(new_n710), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT27), .B(G1996), .Z(new_n714));
  OAI221_X1 g289(.A(new_n701), .B1(new_n693), .B2(new_n692), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  OR3_X1    g290(.A1(new_n695), .A2(KEYINPUT90), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT90), .B1(new_n695), .B2(new_n715), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G19), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n553), .B2(new_n718), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1341), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G168), .B2(new_n718), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n718), .A2(G5), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G171), .B2(new_n718), .ZN(new_n725));
  AOI22_X1  g300(.A1(G1966), .A2(new_n723), .B1(new_n725), .B2(G1961), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G1961), .B2(new_n725), .ZN(new_n727));
  NOR2_X1   g302(.A1(G27), .A2(G29), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G164), .B2(G29), .ZN(new_n729));
  INV_X1    g304(.A(G2078), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G28), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(KEYINPUT30), .ZN(new_n733));
  AOI21_X1  g308(.A(G29), .B1(new_n732), .B2(KEYINPUT30), .ZN(new_n734));
  OR2_X1    g309(.A1(KEYINPUT31), .A2(G11), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n733), .A2(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n633), .B2(new_n690), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n700), .B2(new_n699), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n731), .B(new_n739), .C1(G1966), .C2(new_n723), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n721), .A2(new_n727), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n716), .A2(new_n717), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G4), .A2(G16), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n608), .B2(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G1348), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n718), .A2(G20), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT92), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT23), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n570), .B2(new_n718), .ZN(new_n749));
  INV_X1    g324(.A(G1956), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n713), .A2(new_n714), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n481), .A2(G140), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n483), .A2(G128), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n474), .A2(G116), .ZN(new_n755));
  OAI21_X1  g330(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n753), .B(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G29), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n690), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2067), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AND4_X1   g338(.A1(new_n745), .A2(new_n751), .A3(new_n752), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n690), .A2(G35), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT91), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n690), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT29), .B(G2090), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n764), .B(new_n769), .C1(G1348), .C2(new_n744), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n742), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n718), .A2(G23), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n578), .A2(new_n579), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n718), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT33), .B(G1976), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n774), .B(new_n775), .Z(new_n776));
  NAND2_X1  g351(.A1(G166), .A2(G16), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G16), .B2(G22), .ZN(new_n778));
  INV_X1    g353(.A(G1971), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n776), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G6), .A2(G16), .ZN(new_n783));
  INV_X1    g358(.A(new_n587), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n581), .A2(new_n582), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n783), .B1(new_n786), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT32), .ZN(new_n788));
  INV_X1    g363(.A(G1981), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n782), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(KEYINPUT34), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT34), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n782), .A2(new_n793), .A3(new_n790), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n481), .A2(G131), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n483), .A2(G119), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n474), .A2(G107), .ZN(new_n797));
  OAI21_X1  g372(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n795), .B(new_n796), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G25), .B(new_n799), .S(G29), .Z(new_n800));
  XOR2_X1   g375(.A(KEYINPUT35), .B(G1991), .Z(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n800), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n718), .A2(G24), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n594), .B2(new_n718), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1986), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n792), .A2(new_n794), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT36), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT36), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n771), .B1(new_n809), .B2(new_n810), .ZN(G311));
  INV_X1    g386(.A(KEYINPUT93), .ZN(new_n812));
  XNOR2_X1  g387(.A(G311), .B(new_n812), .ZN(G150));
  AOI22_X1  g388(.A1(new_n577), .A2(G93), .B1(G55), .B2(new_n528), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT94), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(new_n538), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n550), .A2(new_n552), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n815), .A2(new_n549), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT38), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n608), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n826));
  AOI21_X1  g401(.A(G860), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n826), .B2(new_n825), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n818), .A2(G860), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT37), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(G145));
  NAND2_X1  g406(.A1(new_n481), .A2(G142), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT97), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n474), .A2(G118), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n483), .A2(G130), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n623), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n799), .B(KEYINPUT98), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT99), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n757), .B(new_n500), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n709), .ZN(new_n844));
  INV_X1    g419(.A(new_n689), .ZN(new_n845));
  OR3_X1    g420(.A1(new_n844), .A2(KEYINPUT96), .A3(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n689), .B(KEYINPUT96), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n842), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n478), .B(KEYINPUT95), .ZN(new_n851));
  XNOR2_X1  g426(.A(G162), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n633), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n842), .A2(new_n849), .ZN(new_n855));
  INV_X1    g430(.A(new_n849), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n853), .B1(new_n856), .B2(new_n841), .ZN(new_n857));
  AOI21_X1  g432(.A(G37), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g435(.A(KEYINPUT103), .ZN(new_n861));
  INV_X1    g436(.A(new_n818), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(G868), .ZN(new_n863));
  INV_X1    g438(.A(G868), .ZN(new_n864));
  XNOR2_X1  g439(.A(G166), .B(KEYINPUT100), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n786), .ZN(new_n866));
  XNOR2_X1  g441(.A(G288), .B(new_n594), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  OR3_X1    g443(.A1(new_n866), .A2(KEYINPUT102), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT102), .B1(new_n866), .B2(new_n868), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n865), .B(G305), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(new_n867), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n866), .A2(KEYINPUT101), .A3(new_n868), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n869), .A2(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(KEYINPUT42), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(KEYINPUT42), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n822), .B(new_n616), .Z(new_n880));
  NOR2_X1   g455(.A1(new_n608), .A2(new_n570), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n608), .A2(new_n570), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(KEYINPUT41), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n884), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(new_n880), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n864), .B1(new_n879), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n877), .A3(new_n878), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n863), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n878), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n891), .B1(new_n896), .B2(new_n876), .ZN(new_n897));
  AND4_X1   g472(.A1(KEYINPUT103), .A2(new_n894), .A3(new_n897), .A4(G868), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n895), .A2(new_n898), .ZN(G295));
  NOR2_X1   g474(.A1(new_n895), .A2(new_n898), .ZN(G331));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  NOR2_X1   g477(.A1(G171), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(G171), .A2(new_n902), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(G168), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(G286), .A2(G301), .A3(KEYINPUT104), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n822), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n820), .A2(new_n821), .B1(new_n906), .B2(new_n907), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n912), .A3(new_n890), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n886), .B(new_n887), .C1(new_n909), .C2(new_n911), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n901), .B1(new_n915), .B2(new_n875), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n913), .A2(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n869), .A2(new_n870), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n873), .A2(new_n874), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n918), .A2(new_n921), .A3(KEYINPUT105), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n915), .B2(new_n875), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n917), .B(KEYINPUT43), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n918), .A2(new_n921), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n926), .B1(new_n927), .B2(new_n916), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT44), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n917), .B(new_n926), .C1(new_n922), .C2(new_n924), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT43), .B1(new_n927), .B2(new_n916), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n935), .ZN(G397));
  INV_X1    g511(.A(G1384), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(new_n494), .B2(new_n499), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n469), .A2(G40), .A3(new_n475), .A4(new_n477), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n757), .B(new_n762), .ZN(new_n944));
  INV_X1    g519(.A(G1996), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n709), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n709), .A2(new_n945), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n942), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT106), .Z(new_n950));
  NOR2_X1   g525(.A1(new_n799), .A2(new_n802), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n757), .A2(G2067), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n943), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n799), .A2(new_n802), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n942), .B1(new_n955), .B2(new_n951), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n943), .A2(G1986), .A3(G290), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(KEYINPUT48), .Z(new_n958));
  AND3_X1   g533(.A1(new_n950), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n943), .B1(new_n944), .B2(new_n709), .ZN(new_n960));
  OR3_X1    g535(.A1(new_n943), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT46), .B1(new_n943), .B2(G1996), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n954), .A2(new_n959), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G8), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n938), .A2(KEYINPUT50), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n969), .B(new_n937), .C1(new_n494), .C2(new_n499), .ZN(new_n970));
  INV_X1    g545(.A(new_n941), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G2090), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT45), .B(new_n937), .C1(new_n494), .C2(new_n499), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n940), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT108), .B(G1971), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n972), .A2(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n967), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n976), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n941), .B1(new_n938), .B2(KEYINPUT50), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n970), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G2090), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT109), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n510), .A2(KEYINPUT73), .A3(new_n511), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT73), .B1(new_n510), .B2(new_n511), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n518), .A2(new_n519), .B1(G75), .B2(G543), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n538), .B1(new_n990), .B2(new_n521), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT55), .B(G8), .C1(new_n989), .C2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(G303), .A2(KEYINPUT110), .A3(KEYINPUT55), .A4(G8), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n967), .B1(new_n574), .B2(new_n575), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(KEYINPUT55), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT111), .B(new_n1000), .C1(G166), .C2(new_n967), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n996), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n986), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT112), .B1(new_n996), .B2(new_n1002), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n994), .A2(new_n995), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n999), .A4(new_n1001), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1006), .A2(new_n985), .A3(new_n979), .A4(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n938), .A2(new_n941), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(new_n967), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n789), .B1(new_n583), .B2(new_n587), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n784), .A2(new_n785), .A3(G1981), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(KEYINPUT114), .B(new_n1014), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1013), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1015), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n786), .A2(new_n789), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(KEYINPUT49), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT115), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1022), .A2(new_n1023), .A3(new_n1026), .A4(KEYINPUT49), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1012), .B(new_n1029), .C1(new_n1030), .C2(G288), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1012), .A2(new_n1030), .A3(G288), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT113), .B1(new_n773), .B2(G1976), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n773), .A2(G1976), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1035), .B(new_n1012), .C1(new_n1036), .C2(KEYINPUT52), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1021), .A2(new_n1028), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n940), .A2(new_n971), .A3(new_n974), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n1039), .A2(G1966), .B1(new_n983), .B2(G2084), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G8), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(G286), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT63), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1005), .A2(new_n1010), .A3(new_n1038), .A4(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n968), .A2(new_n1047), .A3(new_n971), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n970), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n982), .A2(new_n1047), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT118), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n968), .A2(new_n971), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT117), .ZN(new_n1053));
  INV_X1    g628(.A(new_n970), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n982), .B2(new_n1047), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1051), .A2(new_n973), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n967), .B1(new_n1058), .B2(new_n980), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1010), .B(new_n1038), .C1(new_n1059), .C2(new_n1004), .ZN(new_n1060));
  OAI211_X1 g635(.A(KEYINPUT119), .B(new_n1044), .C1(new_n1060), .C2(new_n1043), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1063));
  AOI21_X1  g638(.A(G2090), .B1(new_n1063), .B2(KEYINPUT118), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n981), .B1(new_n1064), .B2(new_n1057), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1003), .B1(new_n1065), .B2(new_n967), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1066), .A2(new_n1010), .A3(new_n1038), .A4(new_n1042), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT119), .B1(new_n1067), .B2(new_n1044), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1046), .B1(new_n1062), .B2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1012), .B(KEYINPUT116), .ZN(new_n1070));
  AOI211_X1 g645(.A(G1976), .B(G288), .C1(new_n1021), .C2(new_n1028), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n1016), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1038), .A2(new_n986), .A3(new_n1006), .A4(new_n1009), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G286), .A2(G8), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1041), .B(new_n1075), .C1(new_n1076), .C2(KEYINPUT51), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT51), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(G8), .C1(new_n1040), .C2(G286), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1040), .A2(G8), .A3(G286), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1081), .A2(KEYINPUT62), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(KEYINPUT62), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1039), .A2(new_n730), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n975), .A2(G2078), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1088), .A2(KEYINPUT126), .A3(KEYINPUT53), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1085), .A2(new_n1086), .B1(G1961), .B2(new_n972), .ZN(new_n1091));
  OAI21_X1  g666(.A(G171), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1082), .A2(new_n1083), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1060), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1074), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1069), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1091), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1097), .B(G301), .C1(new_n1087), .C2(new_n1089), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1092), .A2(KEYINPUT54), .A3(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1099), .A2(new_n1081), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1092), .A2(new_n1098), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1100), .B(new_n1094), .C1(KEYINPUT54), .C2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT56), .B(G2072), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1039), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1063), .B2(new_n750), .ZN(new_n1106));
  AOI211_X1 g681(.A(KEYINPUT120), .B(G1956), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n570), .B(KEYINPUT57), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n608), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n500), .A2(new_n971), .A3(new_n937), .A4(new_n762), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1011), .A2(KEYINPUT121), .A3(new_n762), .ZN(new_n1116));
  INV_X1    g691(.A(G1348), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1115), .A2(new_n1116), .B1(new_n983), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1111), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1109), .B(new_n1104), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT58), .B(G1341), .ZN(new_n1122));
  OAI22_X1  g697(.A1(new_n975), .A2(G1996), .B1(new_n1011), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n553), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n1127));
  AOI211_X1 g702(.A(new_n1127), .B(new_n608), .C1(new_n1118), .C2(KEYINPUT60), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n983), .A2(new_n1117), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(KEYINPUT60), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1112), .B1(new_n1131), .B2(KEYINPUT123), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1128), .A2(new_n1132), .B1(KEYINPUT123), .B2(new_n1131), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1118), .A2(KEYINPUT60), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1126), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1111), .A2(KEYINPUT61), .A3(new_n1120), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT61), .B1(new_n1111), .B2(new_n1120), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1135), .B(new_n1136), .C1(new_n1137), .C2(KEYINPUT122), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1137), .A2(KEYINPUT122), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1121), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1102), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT124), .B(new_n1121), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1096), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n594), .B(G1986), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n950), .B(new_n956), .C1(new_n943), .C2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(KEYINPUT107), .Z(new_n1147));
  OAI21_X1  g722(.A(new_n966), .B1(new_n1144), .B2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g723(.A(G319), .ZN(new_n1150));
  NOR4_X1   g724(.A1(G229), .A2(new_n1150), .A3(G401), .A4(G227), .ZN(new_n1151));
  NAND3_X1  g725(.A1(new_n933), .A2(new_n1151), .A3(new_n859), .ZN(G225));
  INV_X1    g726(.A(G225), .ZN(G308));
endmodule


