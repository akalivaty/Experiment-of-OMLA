

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594;

  OR2_X1 U324 ( .A1(n592), .A2(n565), .ZN(n507) );
  XNOR2_X1 U325 ( .A(G36GAT), .B(G190GAT), .ZN(n333) );
  XNOR2_X1 U326 ( .A(n333), .B(G218GAT), .ZN(n372) );
  XNOR2_X1 U327 ( .A(n332), .B(n331), .ZN(n341) );
  XNOR2_X1 U328 ( .A(n341), .B(n340), .ZN(n345) );
  XNOR2_X1 U329 ( .A(KEYINPUT122), .B(KEYINPUT55), .ZN(n554) );
  XNOR2_X1 U330 ( .A(n555), .B(n554), .ZN(n570) );
  XOR2_X1 U331 ( .A(n348), .B(n347), .Z(n568) );
  NOR2_X1 U332 ( .A1(n560), .A2(n564), .ZN(n562) );
  XOR2_X1 U333 ( .A(n404), .B(n403), .Z(n556) );
  XOR2_X1 U334 ( .A(KEYINPUT28), .B(n552), .Z(n523) );
  XOR2_X1 U335 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n293) );
  XNOR2_X1 U336 ( .A(KEYINPUT67), .B(KEYINPUT69), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n310) );
  XOR2_X1 U338 ( .A(G113GAT), .B(G36GAT), .Z(n295) );
  XNOR2_X1 U339 ( .A(G169GAT), .B(G50GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U341 ( .A(KEYINPUT68), .B(KEYINPUT66), .Z(n297) );
  XNOR2_X1 U342 ( .A(G197GAT), .B(G8GAT), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U344 ( .A(n299), .B(n298), .Z(n308) );
  XOR2_X1 U345 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n301) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(G29GAT), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U348 ( .A(KEYINPUT7), .B(n302), .ZN(n346) );
  XOR2_X1 U349 ( .A(G141GAT), .B(G22GAT), .Z(n410) );
  XNOR2_X1 U350 ( .A(G15GAT), .B(G1GAT), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n303), .B(KEYINPUT71), .ZN(n354) );
  XOR2_X1 U352 ( .A(n410), .B(n354), .Z(n305) );
  NAND2_X1 U353 ( .A1(G229GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U355 ( .A(n346), .B(n306), .Z(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n581) );
  XOR2_X1 U358 ( .A(G64GAT), .B(KEYINPUT72), .Z(n312) );
  XNOR2_X1 U359 ( .A(G176GAT), .B(G92GAT), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U361 ( .A(G204GAT), .B(n313), .Z(n376) );
  XNOR2_X1 U362 ( .A(G106GAT), .B(G78GAT), .ZN(n316) );
  INV_X1 U363 ( .A(n316), .ZN(n314) );
  NAND2_X1 U364 ( .A1(n314), .A2(G148GAT), .ZN(n318) );
  INV_X1 U365 ( .A(G148GAT), .ZN(n315) );
  NAND2_X1 U366 ( .A1(n316), .A2(n315), .ZN(n317) );
  NAND2_X1 U367 ( .A1(n318), .A2(n317), .ZN(n422) );
  XOR2_X1 U368 ( .A(G99GAT), .B(G85GAT), .Z(n328) );
  XNOR2_X1 U369 ( .A(n422), .B(n328), .ZN(n320) );
  NAND2_X1 U370 ( .A1(G230GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U372 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n322) );
  XNOR2_X1 U373 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n326) );
  XOR2_X1 U376 ( .A(G120GAT), .B(G71GAT), .Z(n396) );
  XOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT13), .Z(n355) );
  XOR2_X1 U378 ( .A(n396), .B(n355), .Z(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U380 ( .A(n376), .B(n327), .Z(n584) );
  INV_X1 U381 ( .A(n584), .ZN(n508) );
  NAND2_X1 U382 ( .A1(n581), .A2(n508), .ZN(n472) );
  XOR2_X1 U383 ( .A(KEYINPUT65), .B(KEYINPUT75), .Z(n330) );
  XOR2_X1 U384 ( .A(G50GAT), .B(G162GAT), .Z(n409) );
  XNOR2_X1 U385 ( .A(n409), .B(n328), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n332) );
  XOR2_X1 U387 ( .A(G134GAT), .B(G106GAT), .Z(n331) );
  NAND2_X1 U388 ( .A1(n372), .A2(KEYINPUT74), .ZN(n337) );
  INV_X1 U389 ( .A(n372), .ZN(n335) );
  INV_X1 U390 ( .A(KEYINPUT74), .ZN(n334) );
  NAND2_X1 U391 ( .A1(n335), .A2(n334), .ZN(n336) );
  NAND2_X1 U392 ( .A1(n337), .A2(n336), .ZN(n339) );
  AND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U395 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n343) );
  XNOR2_X1 U396 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n348) );
  INV_X1 U399 ( .A(n346), .ZN(n347) );
  INV_X1 U400 ( .A(n568), .ZN(n532) );
  XOR2_X1 U401 ( .A(G211GAT), .B(G78GAT), .Z(n350) );
  XNOR2_X1 U402 ( .A(G127GAT), .B(G71GAT), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U404 ( .A(G8GAT), .B(G183GAT), .Z(n379) );
  XOR2_X1 U405 ( .A(n351), .B(n379), .Z(n353) );
  XNOR2_X1 U406 ( .A(G22GAT), .B(G155GAT), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n359) );
  XOR2_X1 U408 ( .A(n355), .B(n354), .Z(n357) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U411 ( .A(n359), .B(n358), .Z(n367) );
  XOR2_X1 U412 ( .A(KEYINPUT15), .B(KEYINPUT76), .Z(n361) );
  XNOR2_X1 U413 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U415 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n363) );
  XNOR2_X1 U416 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U419 ( .A(n367), .B(n366), .Z(n565) );
  NOR2_X1 U420 ( .A1(n532), .A2(n565), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n368), .B(KEYINPUT16), .ZN(n454) );
  XOR2_X1 U422 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n370) );
  XNOR2_X1 U423 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U425 ( .A(G169GAT), .B(n371), .Z(n403) );
  INV_X1 U426 ( .A(n403), .ZN(n385) );
  XOR2_X1 U427 ( .A(n372), .B(KEYINPUT93), .Z(n374) );
  NAND2_X1 U428 ( .A1(G226GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n383) );
  XOR2_X1 U431 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n381) );
  XOR2_X1 U432 ( .A(G211GAT), .B(KEYINPUT21), .Z(n378) );
  XNOR2_X1 U433 ( .A(G197GAT), .B(KEYINPUT87), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n418) );
  XNOR2_X1 U435 ( .A(n418), .B(n379), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U437 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U438 ( .A(n385), .B(n384), .Z(n549) );
  INV_X1 U439 ( .A(n549), .ZN(n500) );
  XOR2_X1 U440 ( .A(KEYINPUT81), .B(G190GAT), .Z(n387) );
  XNOR2_X1 U441 ( .A(G43GAT), .B(G99GAT), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U443 ( .A(G176GAT), .B(G183GAT), .Z(n389) );
  XNOR2_X1 U444 ( .A(G15GAT), .B(KEYINPUT80), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U446 ( .A(n391), .B(n390), .Z(n402) );
  XOR2_X1 U447 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n393) );
  XNOR2_X1 U448 ( .A(KEYINPUT85), .B(KEYINPUT83), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n393), .B(n392), .ZN(n400) );
  XOR2_X1 U450 ( .A(G127GAT), .B(KEYINPUT0), .Z(n395) );
  XNOR2_X1 U451 ( .A(G113GAT), .B(G134GAT), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n441) );
  XOR2_X1 U453 ( .A(n396), .B(n441), .Z(n398) );
  NAND2_X1 U454 ( .A1(G227GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n402), .B(n401), .ZN(n404) );
  NAND2_X1 U458 ( .A1(n500), .A2(n556), .ZN(n424) );
  XOR2_X1 U459 ( .A(G155GAT), .B(KEYINPUT3), .Z(n406) );
  XNOR2_X1 U460 ( .A(KEYINPUT2), .B(KEYINPUT88), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n440) );
  XOR2_X1 U462 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n408) );
  XNOR2_X1 U463 ( .A(KEYINPUT89), .B(G204GAT), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n414) );
  XOR2_X1 U465 ( .A(KEYINPUT22), .B(G218GAT), .Z(n412) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U468 ( .A(n414), .B(n413), .Z(n416) );
  NAND2_X1 U469 ( .A1(G228GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U471 ( .A(n417), .B(KEYINPUT86), .Z(n420) );
  XNOR2_X1 U472 ( .A(n418), .B(KEYINPUT23), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U474 ( .A(n440), .B(n421), .ZN(n423) );
  XNOR2_X1 U475 ( .A(n423), .B(n422), .ZN(n552) );
  NAND2_X1 U476 ( .A1(n424), .A2(n552), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n425), .B(KEYINPUT97), .ZN(n426) );
  XNOR2_X1 U478 ( .A(KEYINPUT25), .B(n426), .ZN(n429) );
  NOR2_X1 U479 ( .A1(n552), .A2(n556), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n427), .B(KEYINPUT26), .ZN(n578) );
  XNOR2_X1 U481 ( .A(KEYINPUT27), .B(n500), .ZN(n449) );
  NAND2_X1 U482 ( .A1(n578), .A2(n449), .ZN(n428) );
  NAND2_X1 U483 ( .A1(n429), .A2(n428), .ZN(n448) );
  XOR2_X1 U484 ( .A(G162GAT), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U485 ( .A(G141GAT), .B(G120GAT), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n433) );
  XOR2_X1 U487 ( .A(G29GAT), .B(G85GAT), .Z(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n445) );
  XOR2_X1 U489 ( .A(G57GAT), .B(KEYINPUT5), .Z(n435) );
  XNOR2_X1 U490 ( .A(KEYINPUT92), .B(KEYINPUT4), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U492 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n437) );
  XNOR2_X1 U493 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U495 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n447) );
  NAND2_X1 U499 ( .A1(G225GAT), .A2(G233GAT), .ZN(n446) );
  XOR2_X1 U500 ( .A(n447), .B(n446), .Z(n577) );
  NAND2_X1 U501 ( .A1(n448), .A2(n577), .ZN(n453) );
  INV_X1 U502 ( .A(n577), .ZN(n497) );
  NAND2_X1 U503 ( .A1(n449), .A2(n497), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n450), .B(KEYINPUT96), .ZN(n521) );
  NOR2_X1 U505 ( .A1(n521), .A2(n523), .ZN(n451) );
  INV_X1 U506 ( .A(n556), .ZN(n567) );
  NAND2_X1 U507 ( .A1(n451), .A2(n567), .ZN(n452) );
  NAND2_X1 U508 ( .A1(n453), .A2(n452), .ZN(n468) );
  NAND2_X1 U509 ( .A1(n454), .A2(n468), .ZN(n483) );
  NOR2_X1 U510 ( .A1(n472), .A2(n483), .ZN(n455) );
  XNOR2_X1 U511 ( .A(KEYINPUT98), .B(n455), .ZN(n465) );
  NAND2_X1 U512 ( .A1(n465), .A2(n497), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n456), .B(KEYINPUT34), .ZN(n457) );
  XNOR2_X1 U514 ( .A(G1GAT), .B(n457), .ZN(G1324GAT) );
  XOR2_X1 U515 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n459) );
  NAND2_X1 U516 ( .A1(n500), .A2(n465), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U518 ( .A(G8GAT), .B(n460), .ZN(G1325GAT) );
  XOR2_X1 U519 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n462) );
  NAND2_X1 U520 ( .A1(n556), .A2(n465), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n462), .B(n461), .ZN(n464) );
  XOR2_X1 U522 ( .A(G15GAT), .B(KEYINPUT101), .Z(n463) );
  XNOR2_X1 U523 ( .A(n464), .B(n463), .ZN(G1326GAT) );
  NAND2_X1 U524 ( .A1(n465), .A2(n523), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n466), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U526 ( .A(G29GAT), .B(KEYINPUT39), .Z(n476) );
  XOR2_X1 U527 ( .A(KEYINPUT36), .B(KEYINPUT103), .Z(n467) );
  XNOR2_X1 U528 ( .A(n568), .B(n467), .ZN(n592) );
  NAND2_X1 U529 ( .A1(n565), .A2(n468), .ZN(n469) );
  NOR2_X1 U530 ( .A1(n592), .A2(n469), .ZN(n471) );
  XNOR2_X1 U531 ( .A(KEYINPUT37), .B(KEYINPUT104), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n471), .B(n470), .ZN(n496) );
  NOR2_X1 U533 ( .A1(n496), .A2(n472), .ZN(n473) );
  XOR2_X1 U534 ( .A(KEYINPUT38), .B(n473), .Z(n474) );
  XNOR2_X1 U535 ( .A(KEYINPUT105), .B(n474), .ZN(n480) );
  NAND2_X1 U536 ( .A1(n497), .A2(n480), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(G1328GAT) );
  NAND2_X1 U538 ( .A1(n480), .A2(n500), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n477), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U540 ( .A1(n480), .A2(n556), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n478), .B(KEYINPUT40), .ZN(n479) );
  XNOR2_X1 U542 ( .A(G43GAT), .B(n479), .ZN(G1330GAT) );
  NAND2_X1 U543 ( .A1(n480), .A2(n523), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n481), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n485) );
  XOR2_X1 U546 ( .A(n508), .B(KEYINPUT41), .Z(n560) );
  INV_X1 U547 ( .A(n560), .ZN(n526) );
  INV_X1 U548 ( .A(n581), .ZN(n557) );
  NAND2_X1 U549 ( .A1(n526), .A2(n557), .ZN(n482) );
  XNOR2_X1 U550 ( .A(n482), .B(KEYINPUT106), .ZN(n495) );
  NOR2_X1 U551 ( .A1(n495), .A2(n483), .ZN(n492) );
  NAND2_X1 U552 ( .A1(n492), .A2(n497), .ZN(n484) );
  XNOR2_X1 U553 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U554 ( .A(G57GAT), .B(n486), .ZN(G1332GAT) );
  NAND2_X1 U555 ( .A1(n492), .A2(n500), .ZN(n487) );
  XNOR2_X1 U556 ( .A(n487), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U557 ( .A1(n492), .A2(n556), .ZN(n488) );
  XNOR2_X1 U558 ( .A(n488), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n490) );
  XNOR2_X1 U560 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n489) );
  XNOR2_X1 U561 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U562 ( .A(KEYINPUT108), .B(n491), .Z(n494) );
  NAND2_X1 U563 ( .A1(n492), .A2(n523), .ZN(n493) );
  XNOR2_X1 U564 ( .A(n494), .B(n493), .ZN(G1335GAT) );
  XOR2_X1 U565 ( .A(G85GAT), .B(KEYINPUT111), .Z(n499) );
  NOR2_X1 U566 ( .A1(n496), .A2(n495), .ZN(n504) );
  NAND2_X1 U567 ( .A1(n504), .A2(n497), .ZN(n498) );
  XNOR2_X1 U568 ( .A(n499), .B(n498), .ZN(G1336GAT) );
  NAND2_X1 U569 ( .A1(n504), .A2(n500), .ZN(n501) );
  XNOR2_X1 U570 ( .A(n501), .B(KEYINPUT112), .ZN(n502) );
  XNOR2_X1 U571 ( .A(G92GAT), .B(n502), .ZN(G1337GAT) );
  NAND2_X1 U572 ( .A1(n504), .A2(n556), .ZN(n503) );
  XNOR2_X1 U573 ( .A(n503), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U574 ( .A1(n523), .A2(n504), .ZN(n505) );
  XNOR2_X1 U575 ( .A(n505), .B(KEYINPUT44), .ZN(n506) );
  XNOR2_X1 U576 ( .A(G106GAT), .B(n506), .ZN(G1339GAT) );
  XOR2_X1 U577 ( .A(G113GAT), .B(KEYINPUT115), .Z(n525) );
  XNOR2_X1 U578 ( .A(n507), .B(KEYINPUT45), .ZN(n510) );
  NAND2_X1 U579 ( .A1(n508), .A2(n557), .ZN(n509) );
  NOR2_X1 U580 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U581 ( .A(n511), .B(KEYINPUT114), .ZN(n518) );
  NOR2_X1 U582 ( .A1(n557), .A2(n560), .ZN(n513) );
  XNOR2_X1 U583 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n512) );
  XNOR2_X1 U584 ( .A(n513), .B(n512), .ZN(n515) );
  INV_X1 U585 ( .A(n565), .ZN(n588) );
  NOR2_X1 U586 ( .A1(n588), .A2(n532), .ZN(n514) );
  AND2_X1 U587 ( .A1(n515), .A2(n514), .ZN(n516) );
  XOR2_X1 U588 ( .A(KEYINPUT47), .B(n516), .Z(n517) );
  NOR2_X1 U589 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U590 ( .A(n519), .B(KEYINPUT64), .ZN(n520) );
  XNOR2_X1 U591 ( .A(n520), .B(KEYINPUT48), .ZN(n550) );
  NOR2_X1 U592 ( .A1(n550), .A2(n521), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n556), .A2(n536), .ZN(n522) );
  NOR2_X1 U594 ( .A1(n523), .A2(n522), .ZN(n533) );
  NAND2_X1 U595 ( .A1(n533), .A2(n581), .ZN(n524) );
  XNOR2_X1 U596 ( .A(n525), .B(n524), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U598 ( .A1(n533), .A2(n526), .ZN(n527) );
  XNOR2_X1 U599 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n530) );
  NAND2_X1 U601 ( .A1(n533), .A2(n588), .ZN(n529) );
  XNOR2_X1 U602 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U603 ( .A(G127GAT), .B(n531), .Z(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n535) );
  NAND2_X1 U605 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U606 ( .A(n535), .B(n534), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n536), .A2(n578), .ZN(n545) );
  NOR2_X1 U608 ( .A1(n557), .A2(n545), .ZN(n537) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n537), .Z(G1344GAT) );
  NOR2_X1 U610 ( .A1(n560), .A2(n545), .ZN(n542) );
  XOR2_X1 U611 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n539) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n538) );
  XNOR2_X1 U613 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U614 ( .A(KEYINPUT117), .B(n540), .ZN(n541) );
  XNOR2_X1 U615 ( .A(n542), .B(n541), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n565), .A2(n545), .ZN(n544) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n543) );
  XNOR2_X1 U618 ( .A(n544), .B(n543), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n568), .A2(n545), .ZN(n547) );
  XNOR2_X1 U620 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n546) );
  XNOR2_X1 U621 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U622 ( .A(G162GAT), .B(n548), .ZN(G1347GAT) );
  NOR2_X1 U623 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U624 ( .A(n551), .B(KEYINPUT54), .ZN(n576) );
  AND2_X1 U625 ( .A1(n577), .A2(n552), .ZN(n553) );
  NAND2_X1 U626 ( .A1(n576), .A2(n553), .ZN(n555) );
  NAND2_X1 U627 ( .A1(n570), .A2(n556), .ZN(n564) );
  NOR2_X1 U628 ( .A1(n564), .A2(n557), .ZN(n558) );
  XNOR2_X1 U629 ( .A(n558), .B(KEYINPUT123), .ZN(n559) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  XNOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n561) );
  XNOR2_X1 U632 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(n563), .ZN(G1349GAT) );
  NOR2_X1 U634 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U635 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  NOR2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U638 ( .A(n571), .B(KEYINPUT58), .Z(n572) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(n572), .ZN(G1351GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n574) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(n575), .Z(n583) );
  AND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(KEYINPUT124), .B(n580), .ZN(n591) );
  INV_X1 U647 ( .A(n591), .ZN(n589) );
  NAND2_X1 U648 ( .A1(n589), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U651 ( .A1(n584), .A2(n589), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U653 ( .A(G204GAT), .B(n587), .Z(G1353GAT) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(KEYINPUT62), .B(n593), .Z(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

