//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1041, new_n1042;
  INV_X1    g000(.A(KEYINPUT5), .ZN(new_n202));
  OR2_X1    g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G141gat), .B(G148gat), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT75), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n203), .A2(new_n209), .A3(new_n204), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n204), .A2(KEYINPUT2), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT76), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT76), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n204), .A2(new_n213), .A3(KEYINPUT2), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n216), .B1(new_n205), .B2(KEYINPUT75), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n208), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G113gat), .ZN(new_n219));
  INV_X1    g018(.A(G120gat), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT1), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G113gat), .A2(G120gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G127gat), .B(G134gat), .Z(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G127gat), .B(G134gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(new_n222), .A3(new_n221), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n218), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G155gat), .B(G162gat), .Z(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(KEYINPUT2), .B2(new_n216), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n206), .B1(new_n231), .B2(new_n209), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n228), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n202), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n242), .B(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n243), .A3(new_n228), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n245));
  INV_X1    g044(.A(new_n227), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n226), .B1(new_n222), .B2(new_n221), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n225), .A2(KEYINPUT68), .A3(new_n227), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n218), .A2(new_n248), .A3(KEYINPUT4), .A4(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n251));
  OAI22_X1  g050(.A1(new_n235), .A2(new_n228), .B1(new_n251), .B2(new_n239), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n244), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n240), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n248), .A2(new_n249), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n251), .B1(new_n255), .B2(new_n235), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n218), .A2(KEYINPUT4), .A3(new_n229), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n256), .A2(new_n244), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G57gat), .B(G85gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(G1gat), .B(G29gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n254), .A2(new_n259), .A3(new_n265), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n260), .A2(KEYINPUT6), .A3(new_n266), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G211gat), .B(G218gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(G197gat), .B(G204gat), .Z(new_n275));
  INV_X1    g074(.A(G211gat), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n276), .A2(KEYINPUT72), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(KEYINPUT72), .ZN(new_n278));
  OAI21_X1  g077(.A(G218gat), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT22), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n275), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n274), .B1(new_n281), .B2(KEYINPUT73), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT72), .B(G211gat), .ZN(new_n283));
  INV_X1    g082(.A(G218gat), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n275), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(new_n288), .A3(new_n273), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT23), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(G169gat), .B2(G176gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n295), .A2(new_n296), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301));
  INV_X1    g100(.A(G183gat), .ZN(new_n302));
  INV_X1    g101(.A(G190gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n303), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n300), .B1(KEYINPUT64), .B2(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n307), .A2(KEYINPUT64), .ZN(new_n309));
  INV_X1    g108(.A(new_n299), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(KEYINPUT23), .B2(new_n294), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n312), .A2(new_n301), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n305), .B1(new_n312), .B2(new_n301), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n311), .B(new_n298), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n308), .A2(new_n309), .B1(new_n315), .B2(KEYINPUT25), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT27), .B(G183gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n303), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT67), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT66), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(KEYINPUT28), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT67), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(new_n322), .A3(new_n303), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n317), .B2(new_n303), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n302), .A2(KEYINPUT27), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT27), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G183gat), .ZN(new_n328));
  AND4_X1   g127(.A1(new_n322), .A2(new_n326), .A3(new_n328), .A4(new_n303), .ZN(new_n329));
  OAI22_X1  g128(.A1(new_n325), .A2(new_n329), .B1(new_n320), .B2(KEYINPUT28), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT26), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n310), .B1(new_n331), .B2(new_n294), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n332), .A2(new_n333), .B1(G183gat), .B2(G190gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n324), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n316), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n293), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n292), .B(KEYINPUT74), .Z(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n316), .B2(new_n335), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n291), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n336), .A2(new_n293), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT29), .B1(new_n316), .B2(new_n335), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n343), .B(new_n290), .C1(new_n344), .C2(new_n339), .ZN(new_n345));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(G64gat), .ZN(new_n347));
  INV_X1    g146(.A(G92gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n342), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n350), .B1(new_n342), .B2(new_n345), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI211_X1 g154(.A(new_n354), .B(new_n350), .C1(new_n342), .C2(new_n345), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n272), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(KEYINPUT69), .B2(KEYINPUT34), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n335), .A2(new_n316), .A3(new_n255), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n255), .B1(new_n335), .B2(new_n316), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT70), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n365), .B(new_n360), .C1(new_n361), .C2(new_n362), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n255), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n336), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n335), .A2(new_n316), .A3(new_n255), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n359), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT33), .ZN(new_n374));
  XOR2_X1   g173(.A(G15gat), .B(G43gat), .Z(new_n375));
  XNOR2_X1  g174(.A(G71gat), .B(G99gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n373), .B(KEYINPUT32), .C1(new_n374), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n373), .A2(KEYINPUT32), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n373), .A2(new_n374), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n377), .ZN(new_n382));
  AOI211_X1 g181(.A(KEYINPUT71), .B(new_n369), .C1(new_n379), .C2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n379), .ZN(new_n385));
  INV_X1    g184(.A(new_n369), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n382), .A2(new_n379), .A3(new_n369), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G228gat), .ZN(new_n391));
  INV_X1    g190(.A(G233gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n287), .A2(new_n273), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n285), .A2(new_n274), .A3(new_n286), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n337), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n218), .B1(new_n397), .B2(new_n242), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n282), .A2(new_n289), .B1(new_n243), .B2(new_n337), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n394), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n282), .A2(new_n289), .A3(new_n337), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n218), .B1(new_n401), .B2(new_n242), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n243), .A2(new_n337), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n290), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n393), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n400), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(G22gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n401), .A2(new_n242), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n235), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n399), .A2(new_n394), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G22gat), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(new_n400), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT78), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n406), .B2(G22gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT31), .B(G50gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n414), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n407), .A2(new_n415), .A3(new_n413), .A4(new_n419), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n390), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n358), .A2(new_n388), .A3(new_n423), .A4(KEYINPUT35), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT35), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n385), .A2(new_n386), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT29), .B1(new_n287), .B2(new_n273), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT3), .B1(new_n427), .B2(new_n396), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n404), .B1(new_n218), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n394), .A2(new_n429), .B1(new_n409), .B2(new_n410), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT78), .B1(new_n430), .B2(new_n412), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n431), .A2(new_n419), .B1(new_n413), .B2(new_n407), .ZN(new_n432));
  INV_X1    g231(.A(new_n422), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n426), .B(new_n389), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n352), .A2(KEYINPUT30), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n435), .A2(new_n356), .A3(new_n351), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n272), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n425), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n424), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n355), .A2(new_n357), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n256), .A2(new_n244), .A3(new_n257), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n441), .A2(new_n239), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT39), .B1(new_n237), .B2(new_n239), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n265), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(KEYINPUT79), .B(KEYINPUT39), .Z(new_n445));
  AND3_X1   g244(.A1(new_n441), .A2(new_n239), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT80), .B1(new_n447), .B2(KEYINPUT40), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n265), .B1(new_n254), .B2(new_n259), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n447), .B2(KEYINPUT40), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT80), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT40), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n451), .B(new_n452), .C1(new_n444), .C2(new_n446), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n440), .A2(new_n448), .A3(new_n450), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n421), .A2(new_n422), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n343), .B(new_n291), .C1(new_n344), .C2(new_n339), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n290), .B1(new_n338), .B2(new_n341), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT37), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n349), .A2(KEYINPUT38), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n342), .A2(new_n345), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT82), .B(KEYINPUT37), .Z(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AOI211_X1 g266(.A(KEYINPUT83), .B(new_n465), .C1(new_n342), .C2(new_n345), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n461), .B(new_n462), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n272), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n353), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n467), .A2(new_n468), .ZN(new_n473));
  INV_X1    g272(.A(new_n464), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n349), .B1(new_n474), .B2(KEYINPUT37), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n454), .B(new_n455), .C1(new_n471), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n426), .A2(KEYINPUT71), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n369), .B1(new_n382), .B2(new_n379), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n384), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n478), .A2(KEYINPUT36), .A3(new_n389), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n426), .A2(new_n389), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n455), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n481), .A2(new_n484), .B1(new_n437), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n439), .B1(new_n477), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G1gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT16), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n412), .A2(G15gat), .ZN(new_n490));
  INV_X1    g289(.A(G15gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G22gat), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n490), .A2(new_n492), .A3(KEYINPUT86), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT86), .B1(new_n490), .B2(new_n492), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n491), .A2(G22gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n412), .A2(G15gat), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n490), .A2(new_n492), .A3(KEYINPUT86), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n488), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n495), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n497), .A2(new_n504), .A3(G8gat), .ZN(new_n505));
  INV_X1    g304(.A(G8gat), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n495), .B(new_n503), .C1(new_n496), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G29gat), .ZN(new_n509));
  INV_X1    g308(.A(G36gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT14), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT14), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(G29gat), .B2(G36gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(G29gat), .A2(G36gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G43gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G50gat), .ZN(new_n517));
  INV_X1    g316(.A(G50gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G43gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n519), .A3(KEYINPUT15), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n515), .B(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT85), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n516), .A2(KEYINPUT85), .A3(G50gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n519), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT15), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n508), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT17), .B1(new_n521), .B2(new_n528), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n515), .A2(KEYINPUT15), .A3(new_n517), .A4(new_n519), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n520), .A2(new_n513), .A3(new_n514), .A4(new_n511), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n536), .A3(new_n527), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n505), .A2(new_n532), .A3(new_n507), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n530), .A2(new_n531), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n530), .A2(KEYINPUT18), .A3(new_n538), .A4(new_n531), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n531), .B(KEYINPUT13), .Z(new_n543));
  NOR2_X1   g342(.A1(new_n508), .A2(new_n529), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n535), .A2(new_n527), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n545), .B1(new_n505), .B2(new_n507), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n543), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n541), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n549));
  XNOR2_X1  g348(.A(G113gat), .B(G141gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT11), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(G169gat), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n550), .A2(KEYINPUT11), .ZN(new_n553));
  INV_X1    g352(.A(G169gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(KEYINPUT11), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(new_n556), .A3(G197gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(G197gat), .B1(new_n552), .B2(new_n556), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n549), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n559), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(KEYINPUT12), .A3(new_n557), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT84), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n563), .B1(new_n560), .B2(new_n562), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n560), .A2(new_n562), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n541), .A2(new_n568), .A3(new_n542), .A4(new_n547), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT88), .B1(new_n487), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n477), .A2(new_n486), .ZN(new_n573));
  AND4_X1   g372(.A1(new_n455), .A2(new_n478), .A3(new_n389), .A4(new_n480), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n437), .A2(new_n425), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n390), .A2(new_n479), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n576), .A2(new_n455), .A3(new_n272), .A4(new_n436), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n574), .A2(new_n575), .B1(new_n577), .B2(new_n425), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT88), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n570), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n572), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT95), .B(G218gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(G99gat), .ZN(new_n585));
  INV_X1    g384(.A(G106gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(KEYINPUT93), .A2(G85gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(KEYINPUT93), .A2(G85gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n592), .A2(new_n348), .B1(KEYINPUT8), .B2(new_n588), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n594));
  OAI211_X1 g393(.A(G85gat), .B(G92gat), .C1(new_n594), .C2(KEYINPUT92), .ZN(new_n595));
  NAND2_X1  g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT92), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n597), .A3(KEYINPUT7), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n589), .B1(new_n593), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n591), .ZN(new_n601));
  NAND2_X1  g400(.A1(KEYINPUT93), .A2(G85gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n348), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT8), .ZN(new_n604));
  AND4_X1   g403(.A1(new_n589), .A2(new_n599), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n529), .A2(new_n606), .B1(KEYINPUT41), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n599), .A2(new_n603), .A3(new_n604), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n588), .A3(new_n587), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n589), .A3(new_n599), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n532), .A2(new_n537), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n607), .A2(KEYINPUT41), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n608), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n616), .B1(new_n608), .B2(new_n613), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT94), .B(G190gat), .ZN(new_n620));
  NOR3_X1   g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n608), .A2(new_n613), .ZN(new_n623));
  INV_X1    g422(.A(new_n616), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n622), .B1(new_n625), .B2(new_n617), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n584), .B1(new_n621), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n620), .B1(new_n618), .B2(new_n619), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n625), .A2(new_n622), .A3(new_n617), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n629), .A3(new_n583), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G57gat), .B(G64gat), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT89), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(G71gat), .A2(G78gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(G71gat), .A2(G78gat), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n638), .B(KEYINPUT89), .C1(new_n634), .C2(new_n633), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT21), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n505), .A2(new_n507), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(new_n302), .ZN(new_n645));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(new_n642), .B2(KEYINPUT21), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT21), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n640), .A2(new_n641), .A3(new_n649), .A4(new_n646), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G127gat), .B(G155gat), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n648), .A2(new_n650), .A3(new_n652), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n654), .B2(new_n657), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n645), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT91), .B(KEYINPUT20), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G211gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n644), .B(G183gat), .ZN(new_n664));
  INV_X1    g463(.A(new_n657), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n652), .B1(new_n648), .B2(new_n650), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n655), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n667), .A3(new_n658), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n661), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n663), .ZN(new_n670));
  INV_X1    g469(.A(new_n668), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n664), .B1(new_n667), .B2(new_n658), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n632), .A2(KEYINPUT96), .A3(new_n669), .A4(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n669), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n676), .B2(new_n631), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G176gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(G204gat), .Z(new_n681));
  OAI211_X1 g480(.A(new_n640), .B(new_n641), .C1(new_n600), .C2(new_n605), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n642), .A2(new_n610), .A3(new_n611), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT10), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n642), .A2(new_n610), .A3(KEYINPUT10), .A4(new_n611), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(G230gat), .A2(G233gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n682), .B2(new_n683), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n681), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n688), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n693), .B1(new_n685), .B2(new_n686), .ZN(new_n694));
  INV_X1    g493(.A(new_n681), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n694), .A2(new_n690), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT97), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n689), .A2(new_n691), .A3(new_n681), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT97), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n695), .B1(new_n694), .B2(new_n690), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n678), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n582), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n470), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g505(.A(new_n580), .B1(new_n579), .B2(new_n570), .ZN(new_n707));
  AOI211_X1 g506(.A(KEYINPUT88), .B(new_n571), .C1(new_n573), .C2(new_n578), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n440), .B(new_n703), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT16), .B(G8gat), .Z(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT98), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n582), .A2(KEYINPUT98), .A3(new_n440), .A4(new_n703), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n716), .A3(new_n711), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n713), .B1(new_n717), .B2(new_n710), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT99), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n716), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(G8gat), .ZN(new_n721));
  AOI211_X1 g520(.A(KEYINPUT99), .B(new_n506), .C1(new_n715), .C2(new_n716), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(G1325gat));
  NAND3_X1  g522(.A1(new_n704), .A2(new_n491), .A3(new_n576), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n481), .A2(new_n484), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n704), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n727), .B2(new_n491), .ZN(G1326gat));
  NAND2_X1  g527(.A1(new_n704), .A2(new_n485), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT43), .B(G22gat), .Z(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT100), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n729), .B(new_n731), .ZN(G1327gat));
  INV_X1    g531(.A(new_n702), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n676), .A2(new_n733), .A3(new_n631), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n572), .B2(new_n581), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n272), .A2(G29gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n735), .A2(KEYINPUT45), .A3(new_n736), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n676), .B(KEYINPUT101), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n702), .B(KEYINPUT102), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n741), .A2(new_n571), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n579), .B2(new_n631), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT103), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n631), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n627), .A2(KEYINPUT103), .A3(new_n630), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI211_X1 g548(.A(KEYINPUT44), .B(new_n749), .C1(new_n573), .C2(new_n578), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n470), .B(new_n743), .C1(new_n745), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G29gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n739), .A2(new_n740), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT104), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n755), .A3(new_n740), .A4(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1328gat));
  NAND3_X1  g556(.A1(new_n735), .A2(new_n510), .A3(new_n440), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT46), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n745), .A2(new_n750), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n743), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n763), .B2(new_n436), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G36gat), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n763), .A2(new_n761), .A3(new_n436), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n760), .B1(new_n765), .B2(new_n766), .ZN(G1329gat));
  NAND3_X1  g566(.A1(new_n735), .A2(new_n516), .A3(new_n576), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n725), .B(new_n743), .C1(new_n745), .C2(new_n750), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n768), .B1(new_n770), .B2(new_n516), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1330gat));
  NOR2_X1   g572(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n455), .A2(G50gat), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n735), .B2(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n485), .B(new_n743), .C1(new_n745), .C2(new_n750), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G50gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1331gat));
  INV_X1    g580(.A(new_n742), .ZN(new_n782));
  NOR4_X1   g581(.A1(new_n487), .A2(new_n570), .A3(new_n678), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n470), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT107), .B(G57gat), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1332gat));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n440), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT49), .B(G64gat), .Z(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n787), .B2(new_n789), .ZN(G1333gat));
  NAND2_X1  g589(.A1(new_n783), .A2(new_n725), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n482), .A2(G71gat), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n791), .A2(G71gat), .B1(new_n783), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g593(.A1(new_n783), .A2(new_n485), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(G78gat), .ZN(G1335gat));
  INV_X1    g595(.A(new_n676), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n570), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n702), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT108), .Z(new_n800));
  AND2_X1   g599(.A1(new_n762), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n470), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n579), .A2(new_n631), .A3(new_n798), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n632), .B1(new_n573), .B2(new_n578), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT51), .B1(new_n809), .B2(new_n798), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n806), .A2(KEYINPUT109), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n470), .A2(new_n592), .A3(new_n702), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT110), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n803), .A2(new_n592), .B1(new_n814), .B2(new_n816), .ZN(G1336gat));
  NOR3_X1   g616(.A1(new_n782), .A2(G92gat), .A3(new_n436), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n812), .A2(new_n813), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n440), .B(new_n800), .C1(new_n745), .C2(new_n750), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G92gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n818), .B1(new_n806), .B2(new_n810), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n824), .B1(new_n826), .B2(KEYINPUT52), .ZN(new_n827));
  AOI211_X1 g626(.A(KEYINPUT111), .B(new_n820), .C1(new_n822), .C2(new_n825), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n823), .B1(new_n827), .B2(new_n828), .ZN(G1337gat));
  NAND2_X1  g628(.A1(new_n801), .A2(new_n725), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G99gat), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n576), .A2(new_n585), .A3(new_n702), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n814), .B2(new_n832), .ZN(G1338gat));
  NAND3_X1  g632(.A1(new_n742), .A2(new_n586), .A3(new_n485), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT112), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n812), .A2(new_n813), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n485), .B(new_n800), .C1(new_n745), .C2(new_n750), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G106gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n835), .B1(new_n806), .B2(new_n810), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n841), .B1(new_n843), .B2(KEYINPUT53), .ZN(new_n844));
  AOI211_X1 g643(.A(KEYINPUT113), .B(new_n837), .C1(new_n839), .C2(new_n842), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n840), .B1(new_n844), .B2(new_n845), .ZN(G1339gat));
  AND4_X1   g645(.A1(new_n571), .A2(new_n674), .A3(new_n677), .A4(new_n733), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n544), .A2(new_n546), .A3(new_n543), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n531), .B1(new_n530), .B2(new_n538), .ZN(new_n849));
  OAI22_X1  g648(.A1(new_n848), .A2(new_n849), .B1(new_n558), .B2(new_n559), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n569), .A2(new_n850), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n686), .A2(new_n693), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT54), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT55), .B1(new_n854), .B2(new_n694), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n687), .A2(new_n856), .A3(new_n688), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n695), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n698), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n853), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n856), .B1(new_n860), .B2(new_n685), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n689), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n681), .B1(new_n694), .B2(new_n856), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT55), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n747), .A2(new_n748), .A3(new_n851), .A4(new_n865), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n570), .A2(new_n865), .B1(new_n702), .B2(new_n851), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n749), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n865), .A2(new_n570), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n702), .A2(new_n851), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n870), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n866), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n741), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n847), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n440), .A2(new_n272), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n875), .A2(new_n434), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(new_n219), .A3(new_n571), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n875), .A2(new_n272), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n436), .A3(new_n574), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n570), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n880), .B1(new_n884), .B2(new_n219), .ZN(G1340gat));
  NOR3_X1   g684(.A1(new_n879), .A2(new_n220), .A3(new_n782), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n702), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n220), .ZN(G1341gat));
  OAI21_X1  g687(.A(G127gat), .B1(new_n879), .B2(new_n874), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n676), .A2(G127gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n882), .B2(new_n890), .ZN(G1342gat));
  NAND2_X1  g690(.A1(new_n881), .A2(new_n574), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n440), .A2(new_n632), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n892), .A2(G134gat), .A3(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n878), .A2(new_n631), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n895), .A2(new_n896), .B1(G134gat), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n899));
  INV_X1    g698(.A(new_n895), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(KEYINPUT56), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n895), .A2(KEYINPUT115), .A3(new_n896), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(G1343gat));
  NOR2_X1   g702(.A1(new_n725), .A2(new_n455), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n870), .A2(new_n871), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT114), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n867), .A2(new_n868), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n907), .A3(new_n749), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n741), .B1(new_n908), .B2(new_n866), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n470), .B(new_n904), .C1(new_n909), .C2(new_n847), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT118), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n571), .A2(G141gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n436), .A3(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n725), .A2(new_n877), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n921), .B1(new_n875), .B2(new_n455), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n455), .A2(new_n921), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OR3_X1    g724(.A1(new_n859), .A2(new_n864), .A3(KEYINPUT116), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT116), .B1(new_n859), .B2(new_n864), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n926), .A2(new_n570), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n631), .B1(new_n928), .B2(new_n871), .ZN(new_n929));
  INV_X1    g728(.A(new_n866), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n676), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n847), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(KEYINPUT117), .B(new_n676), .C1(new_n929), .C2(new_n930), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n925), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n570), .B(new_n920), .C1(new_n923), .C2(new_n935), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n936), .A2(G141gat), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n440), .A2(new_n571), .A3(G141gat), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n936), .A2(G141gat), .B1(new_n911), .B2(new_n938), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n919), .A2(new_n937), .B1(new_n939), .B2(new_n918), .ZN(G1344gat));
  NOR2_X1   g739(.A1(new_n733), .A2(G148gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n915), .A2(new_n436), .A3(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT59), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT57), .B1(new_n875), .B2(new_n455), .ZN(new_n944));
  INV_X1    g743(.A(new_n929), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n865), .A2(new_n631), .A3(new_n851), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n797), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n921), .B(new_n485), .C1(new_n947), .C2(new_n847), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n702), .A3(new_n920), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n943), .B1(new_n950), .B2(G148gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n943), .A2(G148gat), .ZN(new_n952));
  INV_X1    g751(.A(new_n920), .ZN(new_n953));
  INV_X1    g752(.A(new_n935), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(new_n922), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n952), .B1(new_n955), .B2(new_n702), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n942), .B1(new_n951), .B2(new_n956), .ZN(G1345gat));
  INV_X1    g756(.A(KEYINPUT119), .ZN(new_n958));
  INV_X1    g757(.A(G155gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n959), .B1(new_n955), .B2(new_n741), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n797), .A2(new_n959), .ZN(new_n961));
  AOI211_X1 g760(.A(new_n440), .B(new_n961), .C1(new_n912), .C2(new_n914), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n920), .B1(new_n923), .B2(new_n935), .ZN(new_n964));
  OAI21_X1  g763(.A(G155gat), .B1(new_n964), .B2(new_n874), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n915), .A2(new_n436), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n965), .B(KEYINPUT119), .C1(new_n966), .C2(new_n961), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n963), .A2(new_n967), .ZN(G1346gat));
  OAI21_X1  g767(.A(G162gat), .B1(new_n964), .B2(new_n749), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n894), .A2(G162gat), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n915), .A2(KEYINPUT120), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT120), .B1(new_n915), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1347gat));
  NAND2_X1  g772(.A1(new_n574), .A2(new_n440), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT122), .ZN(new_n975));
  OAI21_X1  g774(.A(KEYINPUT121), .B1(new_n875), .B2(new_n470), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n977), .B(new_n272), .C1(new_n909), .C2(new_n847), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n975), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n979), .A2(new_n554), .A3(new_n570), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n470), .A2(new_n436), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  OR3_X1    g781(.A1(new_n875), .A2(new_n434), .A3(new_n982), .ZN(new_n983));
  OR2_X1    g782(.A1(new_n983), .A2(new_n571), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n984), .A2(new_n985), .A3(G169gat), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n985), .B1(new_n984), .B2(G169gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n980), .B1(new_n986), .B2(new_n987), .ZN(G1348gat));
  INV_X1    g787(.A(G176gat), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n983), .A2(new_n989), .A3(new_n782), .ZN(new_n990));
  AOI21_X1  g789(.A(G176gat), .B1(new_n979), .B2(new_n702), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT124), .ZN(new_n992));
  OR2_X1    g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(G1349gat));
  OAI21_X1  g794(.A(G183gat), .B1(new_n983), .B2(new_n874), .ZN(new_n996));
  INV_X1    g795(.A(KEYINPUT125), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n976), .A2(new_n978), .ZN(new_n998));
  INV_X1    g797(.A(new_n975), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n797), .A2(new_n317), .ZN(new_n1000));
  AND4_X1   g799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n997), .B1(new_n979), .B2(new_n1000), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n996), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT60), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT60), .ZN(new_n1005));
  OAI211_X1 g804(.A(new_n1005), .B(new_n996), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(G1350gat));
  INV_X1    g806(.A(KEYINPUT61), .ZN(new_n1008));
  OAI21_X1  g807(.A(G190gat), .B1(new_n983), .B2(new_n632), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1011), .B1(new_n1010), .B2(new_n1009), .ZN(new_n1012));
  INV_X1    g811(.A(new_n749), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n979), .A2(new_n303), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1009), .A2(new_n1010), .A3(new_n1008), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .ZN(G1351gat));
  NOR2_X1   g815(.A1(new_n725), .A2(new_n982), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n949), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g817(.A(G197gat), .B1(new_n1018), .B2(new_n571), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n904), .A2(new_n440), .ZN(new_n1020));
  AOI21_X1  g819(.A(new_n1020), .B1(new_n976), .B2(new_n978), .ZN(new_n1021));
  INV_X1    g820(.A(G197gat), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n1021), .A2(new_n1022), .A3(new_n570), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1019), .A2(new_n1023), .ZN(G1352gat));
  INV_X1    g823(.A(KEYINPUT62), .ZN(new_n1025));
  INV_X1    g824(.A(KEYINPUT127), .ZN(new_n1026));
  NOR2_X1   g825(.A1(new_n733), .A2(G204gat), .ZN(new_n1027));
  NAND3_X1  g826(.A1(new_n1021), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g827(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g828(.A(new_n1026), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1030));
  OAI21_X1  g829(.A(new_n1025), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g830(.A(new_n1030), .ZN(new_n1032));
  NAND3_X1  g831(.A1(new_n1032), .A2(KEYINPUT62), .A3(new_n1028), .ZN(new_n1033));
  OAI21_X1  g832(.A(G204gat), .B1(new_n1018), .B2(new_n782), .ZN(new_n1034));
  NAND3_X1  g833(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(G1353gat));
  NAND3_X1  g834(.A1(new_n1021), .A2(new_n283), .A3(new_n797), .ZN(new_n1036));
  NAND3_X1  g835(.A1(new_n949), .A2(new_n797), .A3(new_n1017), .ZN(new_n1037));
  AND3_X1   g836(.A1(new_n1037), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1038));
  AOI21_X1  g837(.A(KEYINPUT63), .B1(new_n1037), .B2(G211gat), .ZN(new_n1039));
  OAI21_X1  g838(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(G1354gat));
  OAI21_X1  g839(.A(G218gat), .B1(new_n1018), .B2(new_n632), .ZN(new_n1041));
  NAND3_X1  g840(.A1(new_n1021), .A2(new_n284), .A3(new_n1013), .ZN(new_n1042));
  NAND2_X1  g841(.A1(new_n1041), .A2(new_n1042), .ZN(G1355gat));
endmodule


