

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761;

  NOR2_X1 U372 ( .A1(n438), .A2(n394), .ZN(n362) );
  AND2_X1 U373 ( .A1(n378), .A2(n375), .ZN(n384) );
  NOR2_X1 U374 ( .A1(n617), .A2(n432), .ZN(n428) );
  AND2_X1 U375 ( .A1(n391), .A2(n558), .ZN(n648) );
  OR2_X2 U376 ( .A1(n565), .A2(n352), .ZN(n414) );
  INV_X1 U377 ( .A(n356), .ZN(n352) );
  NOR2_X1 U378 ( .A1(n575), .A2(n607), .ZN(n576) );
  XNOR2_X1 U379 ( .A(n746), .B(n467), .ZN(n500) );
  BUF_X1 U380 ( .A(G107), .Z(n408) );
  XNOR2_X1 U381 ( .A(G128), .B(G143), .ZN(n452) );
  AND2_X2 U382 ( .A1(n365), .A2(n360), .ZN(n724) );
  XNOR2_X2 U383 ( .A(n503), .B(n502), .ZN(n678) );
  XNOR2_X2 U384 ( .A(n351), .B(KEYINPUT45), .ZN(n737) );
  NAND2_X1 U385 ( .A1(n384), .A2(n385), .ZN(n351) );
  NOR2_X2 U386 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X2 U387 ( .A1(n571), .A2(n577), .ZN(n608) );
  NAND2_X1 U388 ( .A1(n606), .A2(n673), .ZN(n617) );
  XNOR2_X2 U389 ( .A(n557), .B(KEYINPUT22), .ZN(n565) );
  XNOR2_X1 U390 ( .A(n542), .B(KEYINPUT35), .ZN(n398) );
  XNOR2_X2 U391 ( .A(G116), .B(G113), .ZN(n445) );
  NOR2_X2 U392 ( .A1(n544), .A2(n678), .ZN(n410) );
  INV_X2 U393 ( .A(n547), .ZN(n697) );
  NOR2_X2 U394 ( .A1(n692), .A2(n693), .ZN(n543) );
  XNOR2_X2 U395 ( .A(n506), .B(n443), .ZN(n573) );
  OR2_X2 U396 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X2 U397 ( .A(KEYINPUT90), .B(G110), .ZN(n449) );
  AND2_X1 U398 ( .A1(n363), .A2(n361), .ZN(n360) );
  AND2_X1 U399 ( .A1(n372), .A2(n371), .ZN(n370) );
  XNOR2_X1 U400 ( .A(n454), .B(n453), .ZN(n515) );
  AND2_X1 U401 ( .A1(n617), .A2(n432), .ZN(n430) );
  AND2_X1 U402 ( .A1(n616), .A2(n432), .ZN(n431) );
  NOR2_X1 U403 ( .A1(n756), .A2(KEYINPUT44), .ZN(n371) );
  XNOR2_X1 U404 ( .A(n614), .B(KEYINPUT42), .ZN(n760) );
  NOR2_X2 U405 ( .A1(n613), .A2(n386), .ZN(n658) );
  NOR2_X1 U406 ( .A1(n684), .A2(n682), .ZN(n612) );
  XOR2_X1 U407 ( .A(n644), .B(KEYINPUT62), .Z(n645) );
  XNOR2_X1 U408 ( .A(n493), .B(KEYINPUT21), .ZN(n690) );
  XNOR2_X1 U409 ( .A(n515), .B(n440), .ZN(n393) );
  XNOR2_X1 U410 ( .A(n447), .B(n446), .ZN(n494) );
  XNOR2_X1 U411 ( .A(n482), .B(n481), .ZN(n745) );
  XNOR2_X1 U412 ( .A(KEYINPUT64), .B(n736), .ZN(n749) );
  XNOR2_X1 U413 ( .A(KEYINPUT66), .B(KEYINPUT79), .ZN(n453) );
  XOR2_X1 U414 ( .A(KEYINPUT69), .B(G101), .Z(n466) );
  XOR2_X1 U415 ( .A(G122), .B(KEYINPUT16), .Z(n451) );
  XOR2_X1 U416 ( .A(G146), .B(G125), .Z(n480) );
  INV_X1 U417 ( .A(n398), .ZN(n372) );
  NAND2_X1 U418 ( .A1(n411), .A2(n427), .ZN(n433) );
  NOR2_X1 U419 ( .A1(n430), .A2(n431), .ZN(n411) );
  INV_X1 U420 ( .A(n514), .ZN(n425) );
  XOR2_X1 U421 ( .A(G902), .B(KEYINPUT15), .Z(n474) );
  XNOR2_X1 U422 ( .A(n393), .B(n465), .ZN(n746) );
  XNOR2_X1 U423 ( .A(n464), .B(G137), .ZN(n465) );
  XNOR2_X1 U424 ( .A(G134), .B(G131), .ZN(n464) );
  INV_X1 U425 ( .A(G469), .ZN(n442) );
  NOR2_X1 U426 ( .A1(G902), .A2(n723), .ZN(n473) );
  INV_X1 U427 ( .A(n554), .ZN(n434) );
  INV_X1 U428 ( .A(G953), .ZN(n736) );
  XOR2_X1 U429 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n529) );
  XNOR2_X1 U430 ( .A(G122), .B(KEYINPUT99), .ZN(n528) );
  XOR2_X1 U431 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n527) );
  XNOR2_X1 U432 ( .A(n495), .B(KEYINPUT96), .ZN(n416) );
  NOR2_X1 U433 ( .A1(G237), .A2(G953), .ZN(n496) );
  NAND2_X1 U434 ( .A1(n433), .A2(n353), .ZN(n438) );
  INV_X1 U435 ( .A(KEYINPUT78), .ZN(n456) );
  XNOR2_X1 U436 ( .A(n455), .B(KEYINPUT65), .ZN(n440) );
  INV_X1 U437 ( .A(KEYINPUT4), .ZN(n455) );
  AND2_X1 U438 ( .A1(n392), .A2(n355), .ZN(n373) );
  NOR2_X1 U439 ( .A1(n392), .A2(KEYINPUT84), .ZN(n383) );
  AND2_X1 U440 ( .A1(n377), .A2(n376), .ZN(n375) );
  NAND2_X1 U441 ( .A1(n433), .A2(n625), .ZN(n368) );
  XNOR2_X1 U442 ( .A(KEYINPUT38), .B(n607), .ZN(n680) );
  NOR2_X1 U443 ( .A1(n730), .A2(G902), .ZN(n490) );
  NAND2_X1 U444 ( .A1(n425), .A2(n426), .ZN(n424) );
  NAND2_X1 U445 ( .A1(KEYINPUT87), .A2(n514), .ZN(n423) );
  NAND2_X1 U446 ( .A1(n425), .A2(KEYINPUT87), .ZN(n421) );
  NAND2_X1 U447 ( .A1(n514), .A2(n426), .ZN(n420) );
  INV_X1 U448 ( .A(KEYINPUT1), .ZN(n441) );
  XOR2_X1 U449 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n487) );
  XNOR2_X1 U450 ( .A(KEYINPUT23), .B(KEYINPUT92), .ZN(n483) );
  XOR2_X1 U451 ( .A(KEYINPUT93), .B(KEYINPUT24), .Z(n484) );
  XNOR2_X1 U452 ( .A(G137), .B(G128), .ZN(n478) );
  XOR2_X1 U453 ( .A(G110), .B(G119), .Z(n479) );
  XOR2_X1 U454 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n482) );
  XNOR2_X1 U455 ( .A(n480), .B(G140), .ZN(n481) );
  XNOR2_X1 U456 ( .A(n466), .B(G146), .ZN(n467) );
  BUF_X1 U457 ( .A(n573), .Z(n574) );
  INV_X1 U458 ( .A(KEYINPUT85), .ZN(n508) );
  XNOR2_X1 U459 ( .A(n396), .B(KEYINPUT30), .ZN(n395) );
  INV_X1 U460 ( .A(n692), .ZN(n621) );
  INV_X1 U461 ( .A(KEYINPUT80), .ZN(n369) );
  INV_X1 U462 ( .A(KEYINPUT48), .ZN(n432) );
  INV_X1 U463 ( .A(KEYINPUT84), .ZN(n389) );
  XNOR2_X1 U464 ( .A(G134), .B(n408), .ZN(n516) );
  XNOR2_X1 U465 ( .A(G116), .B(G122), .ZN(n517) );
  XNOR2_X1 U466 ( .A(G113), .B(G104), .ZN(n526) );
  XNOR2_X1 U467 ( .A(G143), .B(G131), .ZN(n532) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n509) );
  OR2_X1 U469 ( .A1(G237), .A2(G902), .ZN(n507) );
  INV_X1 U470 ( .A(n679), .ZN(n397) );
  XNOR2_X1 U471 ( .A(n494), .B(n416), .ZN(n498) );
  NOR2_X1 U472 ( .A1(n368), .A2(n677), .ZN(n364) );
  NAND2_X1 U473 ( .A1(n354), .A2(n439), .ZN(n394) );
  XNOR2_X1 U474 ( .A(n403), .B(n402), .ZN(n505) );
  XNOR2_X1 U475 ( .A(n740), .B(n404), .ZN(n403) );
  INV_X1 U476 ( .A(n368), .ZN(n748) );
  NAND2_X1 U477 ( .A1(G214), .A2(n507), .ZN(n679) );
  AND2_X1 U478 ( .A1(n680), .A2(n608), .ZN(n609) );
  NOR2_X1 U479 ( .A1(n693), .A2(n546), .ZN(n570) );
  NAND2_X1 U480 ( .A1(n424), .A2(n423), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n414), .B(KEYINPUT83), .ZN(n391) );
  XNOR2_X1 U482 ( .A(n435), .B(n488), .ZN(n730) );
  XNOR2_X1 U483 ( .A(n745), .B(n436), .ZN(n435) );
  XNOR2_X1 U484 ( .A(n489), .B(n485), .ZN(n436) );
  XNOR2_X1 U485 ( .A(n632), .B(KEYINPUT123), .ZN(n634) );
  XNOR2_X1 U486 ( .A(n638), .B(n637), .ZN(n639) );
  XOR2_X1 U487 ( .A(KEYINPUT77), .B(G140), .Z(n469) );
  XOR2_X1 U488 ( .A(KEYINPUT88), .B(n629), .Z(n727) );
  NOR2_X1 U489 ( .A1(n697), .A2(n565), .ZN(n559) );
  AND2_X1 U490 ( .A1(n625), .A2(n504), .ZN(n353) );
  OR2_X1 U491 ( .A1(n626), .A2(n677), .ZN(n354) );
  AND2_X1 U492 ( .A1(n551), .A2(KEYINPUT84), .ZN(n355) );
  AND2_X1 U493 ( .A1(n562), .A2(n692), .ZN(n356) );
  AND2_X1 U494 ( .A1(n558), .A2(n389), .ZN(n357) );
  AND2_X1 U495 ( .A1(n421), .A2(n420), .ZN(n358) );
  INV_X1 U496 ( .A(KEYINPUT87), .ZN(n426) );
  XNOR2_X1 U497 ( .A(KEYINPUT89), .B(n474), .ZN(n626) );
  INV_X1 U498 ( .A(KEYINPUT82), .ZN(n439) );
  NAND2_X1 U499 ( .A1(n359), .A2(n437), .ZN(n366) );
  OR2_X2 U500 ( .A1(n737), .A2(n439), .ZN(n359) );
  NOR2_X1 U501 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U502 ( .A1(n737), .A2(n362), .ZN(n361) );
  NAND2_X1 U503 ( .A1(n737), .A2(n364), .ZN(n363) );
  NAND2_X1 U504 ( .A1(n366), .A2(n354), .ZN(n365) );
  NAND2_X1 U505 ( .A1(n367), .A2(n589), .ZN(n590) );
  NAND2_X1 U506 ( .A1(n662), .A2(KEYINPUT80), .ZN(n367) );
  INV_X1 U507 ( .A(n658), .ZN(n662) );
  NAND2_X1 U508 ( .A1(n658), .A2(n369), .ZN(n586) );
  XNOR2_X1 U509 ( .A(n547), .B(KEYINPUT6), .ZN(n599) );
  XNOR2_X2 U510 ( .A(n501), .B(G472), .ZN(n547) );
  NAND2_X1 U511 ( .A1(n398), .A2(KEYINPUT44), .ZN(n392) );
  INV_X1 U512 ( .A(n648), .ZN(n374) );
  NAND2_X1 U513 ( .A1(n573), .A2(n679), .ZN(n387) );
  NAND2_X1 U514 ( .A1(n418), .A2(n417), .ZN(n556) );
  XNOR2_X1 U515 ( .A(n612), .B(KEYINPUT41), .ZN(n709) );
  NAND2_X1 U516 ( .A1(n724), .A2(G210), .ZN(n627) );
  NAND2_X1 U517 ( .A1(n760), .A2(n759), .ZN(n615) );
  NAND2_X1 U518 ( .A1(n370), .A2(n379), .ZN(n378) );
  NAND2_X1 U519 ( .A1(n374), .A2(n373), .ZN(n380) );
  NAND2_X1 U520 ( .A1(n756), .A2(KEYINPUT44), .ZN(n376) );
  NAND2_X1 U521 ( .A1(n656), .A2(KEYINPUT44), .ZN(n377) );
  INV_X1 U522 ( .A(n656), .ZN(n379) );
  NAND2_X1 U523 ( .A1(n380), .A2(n381), .ZN(n385) );
  NAND2_X1 U524 ( .A1(n388), .A2(n390), .ZN(n382) );
  INV_X1 U525 ( .A(n401), .ZN(n386) );
  XNOR2_X2 U526 ( .A(n602), .B(KEYINPUT19), .ZN(n401) );
  XNOR2_X2 U527 ( .A(n387), .B(n508), .ZN(n602) );
  NAND2_X1 U528 ( .A1(n391), .A2(n357), .ZN(n388) );
  OR2_X1 U529 ( .A1(n551), .A2(KEYINPUT84), .ZN(n390) );
  XNOR2_X1 U530 ( .A(n393), .B(n459), .ZN(n402) );
  NAND2_X1 U531 ( .A1(n570), .A2(n395), .ZN(n571) );
  NOR2_X1 U532 ( .A1(n547), .A2(n397), .ZN(n396) );
  XNOR2_X1 U533 ( .A(n372), .B(G122), .ZN(G24) );
  NAND2_X1 U534 ( .A1(n401), .A2(n399), .ZN(n419) );
  INV_X1 U535 ( .A(n513), .ZN(n399) );
  NAND2_X1 U536 ( .A1(n401), .A2(n400), .ZN(n417) );
  NOR2_X1 U537 ( .A1(n513), .A2(n358), .ZN(n400) );
  XNOR2_X1 U538 ( .A(n458), .B(n460), .ZN(n404) );
  XNOR2_X2 U539 ( .A(n409), .B(n494), .ZN(n740) );
  XNOR2_X2 U540 ( .A(n407), .B(KEYINPUT32), .ZN(n756) );
  NOR2_X2 U541 ( .A1(n565), .A2(n564), .ZN(n407) );
  XNOR2_X1 U542 ( .A(n457), .B(n456), .ZN(n459) );
  NAND2_X1 U543 ( .A1(n419), .A2(n422), .ZN(n418) );
  XNOR2_X2 U544 ( .A(n470), .B(n451), .ZN(n409) );
  XNOR2_X1 U545 ( .A(n410), .B(KEYINPUT34), .ZN(n541) );
  NAND2_X1 U546 ( .A1(n724), .A2(G472), .ZN(n646) );
  NAND2_X1 U547 ( .A1(n412), .A2(n727), .ZN(n631) );
  XNOR2_X1 U548 ( .A(n627), .B(n628), .ZN(n412) );
  NAND2_X1 U549 ( .A1(n413), .A2(n727), .ZN(n636) );
  XNOR2_X1 U550 ( .A(n633), .B(n634), .ZN(n413) );
  XNOR2_X1 U551 ( .A(n415), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U552 ( .A1(n647), .A2(n727), .ZN(n415) );
  NAND2_X1 U553 ( .A1(n608), .A2(n572), .ZN(n575) );
  NAND2_X1 U554 ( .A1(n428), .A2(n429), .ZN(n427) );
  NOR2_X2 U555 ( .A1(n560), .A2(n621), .ZN(n656) );
  NAND2_X1 U556 ( .A1(n737), .A2(n748), .ZN(n676) );
  INV_X1 U557 ( .A(n616), .ZN(n429) );
  INV_X1 U558 ( .A(n580), .ZN(n689) );
  NAND2_X1 U559 ( .A1(n580), .A2(n434), .ZN(n693) );
  NAND2_X1 U560 ( .A1(n438), .A2(KEYINPUT82), .ZN(n437) );
  XNOR2_X2 U561 ( .A(n585), .B(n441), .ZN(n692) );
  XNOR2_X2 U562 ( .A(n473), .B(n442), .ZN(n585) );
  NAND2_X1 U563 ( .A1(n621), .A2(n689), .ZN(n561) );
  INV_X1 U564 ( .A(n689), .ZN(n558) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(n644) );
  AND2_X1 U566 ( .A1(G210), .A2(n507), .ZN(n443) );
  XNOR2_X1 U567 ( .A(G104), .B(G107), .ZN(n448) );
  INV_X1 U568 ( .A(KEYINPUT73), .ZN(n444) );
  XNOR2_X1 U569 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U570 ( .A(n470), .B(n471), .ZN(n472) );
  XNOR2_X1 U571 ( .A(n500), .B(n472), .ZN(n723) );
  INV_X1 U572 ( .A(KEYINPUT124), .ZN(n635) );
  XNOR2_X1 U573 ( .A(n445), .B(n444), .ZN(n447) );
  XOR2_X1 U574 ( .A(KEYINPUT3), .B(G119), .Z(n446) );
  INV_X1 U575 ( .A(n448), .ZN(n450) );
  XNOR2_X2 U576 ( .A(n450), .B(n449), .ZN(n470) );
  INV_X1 U577 ( .A(n452), .ZN(n454) );
  NAND2_X1 U578 ( .A1(G224), .A2(n749), .ZN(n457) );
  XOR2_X1 U579 ( .A(n466), .B(KEYINPUT17), .Z(n458) );
  XNOR2_X1 U580 ( .A(n480), .B(KEYINPUT18), .ZN(n460) );
  XOR2_X1 U581 ( .A(KEYINPUT55), .B(KEYINPUT86), .Z(n462) );
  XNOR2_X1 U582 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n461) );
  XNOR2_X1 U583 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U584 ( .A(n505), .B(n463), .ZN(n628) );
  NAND2_X1 U585 ( .A1(G227), .A2(n749), .ZN(n468) );
  XNOR2_X1 U586 ( .A(n469), .B(n468), .ZN(n471) );
  XOR2_X1 U587 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n477) );
  NAND2_X1 U588 ( .A1(n626), .A2(G234), .ZN(n475) );
  XNOR2_X1 U589 ( .A(n475), .B(KEYINPUT20), .ZN(n492) );
  NAND2_X1 U590 ( .A1(G217), .A2(n492), .ZN(n476) );
  XNOR2_X1 U591 ( .A(n477), .B(n476), .ZN(n491) );
  XNOR2_X1 U592 ( .A(n479), .B(n478), .ZN(n489) );
  XNOR2_X1 U593 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U594 ( .A1(G234), .A2(n749), .ZN(n486) );
  XNOR2_X1 U595 ( .A(n487), .B(n486), .ZN(n521) );
  NAND2_X1 U596 ( .A1(n521), .A2(G221), .ZN(n488) );
  XOR2_X1 U597 ( .A(n491), .B(n490), .Z(n580) );
  NAND2_X1 U598 ( .A1(n492), .A2(G221), .ZN(n493) );
  XOR2_X1 U599 ( .A(n690), .B(KEYINPUT95), .Z(n554) );
  XOR2_X1 U600 ( .A(KEYINPUT5), .B(KEYINPUT75), .Z(n495) );
  XNOR2_X1 U601 ( .A(n496), .B(KEYINPUT76), .ZN(n535) );
  AND2_X1 U602 ( .A1(G210), .A2(n535), .ZN(n497) );
  NOR2_X1 U603 ( .A1(n644), .A2(G902), .ZN(n501) );
  NAND2_X1 U604 ( .A1(n543), .A2(n599), .ZN(n503) );
  XOR2_X1 U605 ( .A(KEYINPUT102), .B(KEYINPUT33), .Z(n502) );
  INV_X1 U606 ( .A(n626), .ZN(n504) );
  XNOR2_X1 U607 ( .A(n509), .B(KEYINPUT91), .ZN(n510) );
  XOR2_X1 U608 ( .A(KEYINPUT14), .B(n510), .Z(n511) );
  NAND2_X1 U609 ( .A1(G952), .A2(n511), .ZN(n708) );
  NOR2_X1 U610 ( .A1(G953), .A2(n708), .ZN(n568) );
  NAND2_X1 U611 ( .A1(G902), .A2(n511), .ZN(n566) );
  OR2_X1 U612 ( .A1(n736), .A2(G898), .ZN(n742) );
  NOR2_X1 U613 ( .A1(n566), .A2(n742), .ZN(n512) );
  NOR2_X1 U614 ( .A1(n568), .A2(n512), .ZN(n513) );
  XNOR2_X1 U615 ( .A(KEYINPUT0), .B(KEYINPUT68), .ZN(n514) );
  INV_X1 U616 ( .A(n556), .ZN(n544) );
  XNOR2_X1 U617 ( .A(n516), .B(KEYINPUT100), .ZN(n520) );
  XOR2_X1 U618 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n518) );
  XNOR2_X1 U619 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U620 ( .A(n520), .B(n519), .Z(n523) );
  NAND2_X1 U621 ( .A1(G217), .A2(n521), .ZN(n522) );
  XNOR2_X1 U622 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U623 ( .A(n515), .B(n524), .ZN(n632) );
  NOR2_X1 U624 ( .A1(n632), .A2(G902), .ZN(n525) );
  XNOR2_X1 U625 ( .A(n525), .B(G478), .ZN(n549) );
  INV_X1 U626 ( .A(n549), .ZN(n552) );
  XNOR2_X1 U627 ( .A(KEYINPUT13), .B(G475), .ZN(n539) );
  XNOR2_X1 U628 ( .A(n527), .B(n526), .ZN(n531) );
  XNOR2_X1 U629 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U630 ( .A(n531), .B(n530), .Z(n533) );
  XNOR2_X1 U631 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U632 ( .A(n745), .B(n534), .Z(n537) );
  NAND2_X1 U633 ( .A1(G214), .A2(n535), .ZN(n536) );
  XNOR2_X1 U634 ( .A(n537), .B(n536), .ZN(n638) );
  NOR2_X1 U635 ( .A1(G902), .A2(n638), .ZN(n538) );
  XNOR2_X1 U636 ( .A(n539), .B(n538), .ZN(n553) );
  NAND2_X1 U637 ( .A1(n552), .A2(n553), .ZN(n540) );
  XNOR2_X1 U638 ( .A(n540), .B(KEYINPUT103), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n541), .A2(n572), .ZN(n542) );
  NAND2_X1 U640 ( .A1(n697), .A2(n543), .ZN(n701) );
  NOR2_X1 U641 ( .A1(n544), .A2(n701), .ZN(n545) );
  XNOR2_X1 U642 ( .A(n545), .B(KEYINPUT31), .ZN(n667) );
  INV_X1 U643 ( .A(n585), .ZN(n546) );
  AND2_X1 U644 ( .A1(n556), .A2(n570), .ZN(n548) );
  NAND2_X1 U645 ( .A1(n548), .A2(n547), .ZN(n652) );
  NAND2_X1 U646 ( .A1(n667), .A2(n652), .ZN(n550) );
  NAND2_X1 U647 ( .A1(n553), .A2(n549), .ZN(n665) );
  NOR2_X1 U648 ( .A1(n549), .A2(n553), .ZN(n657) );
  INV_X1 U649 ( .A(n657), .ZN(n668) );
  NAND2_X1 U650 ( .A1(n665), .A2(n668), .ZN(n683) );
  NAND2_X1 U651 ( .A1(n550), .A2(n683), .ZN(n551) );
  OR2_X1 U652 ( .A1(n553), .A2(n552), .ZN(n682) );
  NOR2_X1 U653 ( .A1(n682), .A2(n554), .ZN(n555) );
  NAND2_X1 U654 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U655 ( .A1(n559), .A2(n689), .ZN(n560) );
  XNOR2_X1 U656 ( .A(KEYINPUT101), .B(n561), .ZN(n563) );
  INV_X1 U657 ( .A(n599), .ZN(n562) );
  NAND2_X1 U658 ( .A1(n563), .A2(n562), .ZN(n564) );
  OR2_X1 U659 ( .A1(n566), .A2(n749), .ZN(n567) );
  NOR2_X1 U660 ( .A1(G900), .A2(n567), .ZN(n569) );
  NOR2_X1 U661 ( .A1(n569), .A2(n568), .ZN(n577) );
  INV_X1 U662 ( .A(n574), .ZN(n607) );
  XNOR2_X1 U663 ( .A(n576), .B(KEYINPUT104), .ZN(n757) );
  NAND2_X1 U664 ( .A1(KEYINPUT81), .A2(n683), .ZN(n587) );
  NOR2_X1 U665 ( .A1(n690), .A2(n577), .ZN(n578) );
  XOR2_X1 U666 ( .A(KEYINPUT72), .B(n578), .Z(n579) );
  NOR2_X1 U667 ( .A1(n580), .A2(n579), .ZN(n600) );
  AND2_X1 U668 ( .A1(n697), .A2(n600), .ZN(n583) );
  XOR2_X1 U669 ( .A(KEYINPUT105), .B(KEYINPUT28), .Z(n581) );
  XNOR2_X1 U670 ( .A(KEYINPUT106), .B(n581), .ZN(n582) );
  XNOR2_X1 U671 ( .A(n583), .B(n582), .ZN(n584) );
  NAND2_X1 U672 ( .A1(n585), .A2(n584), .ZN(n613) );
  NAND2_X1 U673 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U674 ( .A1(n757), .A2(n588), .ZN(n592) );
  OR2_X1 U675 ( .A1(n683), .A2(KEYINPUT81), .ZN(n589) );
  NAND2_X1 U676 ( .A1(KEYINPUT47), .A2(n590), .ZN(n591) );
  NAND2_X1 U677 ( .A1(n592), .A2(n591), .ZN(n597) );
  NAND2_X1 U678 ( .A1(n658), .A2(n683), .ZN(n593) );
  NAND2_X1 U679 ( .A1(KEYINPUT80), .A2(n593), .ZN(n594) );
  NOR2_X1 U680 ( .A1(KEYINPUT81), .A2(n594), .ZN(n595) );
  NOR2_X1 U681 ( .A1(KEYINPUT47), .A2(n595), .ZN(n596) );
  XNOR2_X1 U682 ( .A(n598), .B(KEYINPUT74), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U684 ( .A1(n665), .A2(n601), .ZN(n619) );
  INV_X1 U685 ( .A(n619), .ZN(n603) );
  NOR2_X1 U686 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U687 ( .A(n604), .B(KEYINPUT36), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n605), .A2(n621), .ZN(n673) );
  XNOR2_X1 U689 ( .A(n609), .B(KEYINPUT39), .ZN(n618) );
  NOR2_X1 U690 ( .A1(n665), .A2(n618), .ZN(n611) );
  XNOR2_X1 U691 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n610) );
  XNOR2_X1 U692 ( .A(n611), .B(n610), .ZN(n759) );
  NAND2_X1 U693 ( .A1(n680), .A2(n679), .ZN(n684) );
  OR2_X1 U694 ( .A1(n709), .A2(n613), .ZN(n614) );
  XNOR2_X1 U695 ( .A(n615), .B(KEYINPUT46), .ZN(n616) );
  OR2_X1 U696 ( .A1(n618), .A2(n668), .ZN(n674) );
  NAND2_X1 U697 ( .A1(n619), .A2(n679), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n622), .B(KEYINPUT43), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n574), .A2(n623), .ZN(n675) );
  INV_X1 U701 ( .A(n675), .ZN(n624) );
  AND2_X1 U702 ( .A1(n674), .A2(n624), .ZN(n625) );
  INV_X1 U703 ( .A(KEYINPUT2), .ZN(n677) );
  NOR2_X1 U704 ( .A1(n749), .A2(G952), .ZN(n629) );
  XOR2_X1 U705 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n630) );
  XNOR2_X1 U706 ( .A(n631), .B(n630), .ZN(G51) );
  NAND2_X1 U707 ( .A1(n724), .A2(G478), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(G63) );
  NAND2_X1 U709 ( .A1(n724), .A2(G475), .ZN(n640) );
  XOR2_X1 U710 ( .A(KEYINPUT59), .B(KEYINPUT67), .Z(n637) );
  XNOR2_X1 U711 ( .A(n640), .B(n639), .ZN(n641) );
  NAND2_X1 U712 ( .A1(n641), .A2(n727), .ZN(n643) );
  INV_X1 U713 ( .A(KEYINPUT60), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n643), .B(n642), .ZN(G60) );
  XNOR2_X1 U715 ( .A(n646), .B(n645), .ZN(n647) );
  XOR2_X1 U716 ( .A(n648), .B(G101), .Z(n649) );
  XNOR2_X1 U717 ( .A(KEYINPUT108), .B(n649), .ZN(G3) );
  NOR2_X1 U718 ( .A1(n665), .A2(n652), .ZN(n651) );
  XNOR2_X1 U719 ( .A(G104), .B(KEYINPUT109), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n651), .B(n650), .ZN(G6) );
  NOR2_X1 U721 ( .A1(n668), .A2(n652), .ZN(n654) );
  XNOR2_X1 U722 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U724 ( .A(n408), .B(n655), .ZN(G9) );
  XOR2_X1 U725 ( .A(G110), .B(n656), .Z(G12) );
  XOR2_X1 U726 ( .A(KEYINPUT29), .B(KEYINPUT110), .Z(n660) );
  NAND2_X1 U727 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U729 ( .A(G128), .B(n661), .ZN(G30) );
  NOR2_X1 U730 ( .A1(n665), .A2(n662), .ZN(n663) );
  XOR2_X1 U731 ( .A(KEYINPUT112), .B(n663), .Z(n664) );
  XNOR2_X1 U732 ( .A(G146), .B(n664), .ZN(G48) );
  NOR2_X1 U733 ( .A1(n665), .A2(n667), .ZN(n666) );
  XOR2_X1 U734 ( .A(G113), .B(n666), .Z(G15) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n670) );
  XNOR2_X1 U736 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n669) );
  XNOR2_X1 U737 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U738 ( .A(G116), .B(n671), .ZN(G18) );
  XOR2_X1 U739 ( .A(G125), .B(KEYINPUT37), .Z(n672) );
  XNOR2_X1 U740 ( .A(n673), .B(n672), .ZN(G27) );
  XNOR2_X1 U741 ( .A(G134), .B(n674), .ZN(G36) );
  XOR2_X1 U742 ( .A(G140), .B(n675), .Z(G42) );
  XNOR2_X1 U743 ( .A(n677), .B(n676), .ZN(n717) );
  BUF_X1 U744 ( .A(n678), .Z(n710) );
  NOR2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n687) );
  INV_X1 U747 ( .A(n683), .ZN(n685) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U749 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n710), .A2(n688), .ZN(n705) );
  NAND2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U752 ( .A(KEYINPUT49), .B(n691), .Z(n699) );
  NAND2_X1 U753 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U754 ( .A(n694), .B(KEYINPUT50), .ZN(n695) );
  XNOR2_X1 U755 ( .A(KEYINPUT115), .B(n695), .ZN(n696) );
  NOR2_X1 U756 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U757 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U758 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U759 ( .A(KEYINPUT51), .B(n702), .ZN(n703) );
  NOR2_X1 U760 ( .A1(n703), .A2(n709), .ZN(n704) );
  NOR2_X1 U761 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U762 ( .A(n706), .B(KEYINPUT52), .ZN(n707) );
  NOR2_X1 U763 ( .A1(n708), .A2(n707), .ZN(n713) );
  NOR2_X1 U764 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n711), .B(KEYINPUT116), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U767 ( .A(n714), .B(KEYINPUT117), .ZN(n715) );
  NOR2_X1 U768 ( .A1(G953), .A2(n715), .ZN(n716) );
  NAND2_X1 U769 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U770 ( .A(n718), .B(KEYINPUT118), .ZN(n719) );
  XOR2_X1 U771 ( .A(KEYINPUT53), .B(n719), .Z(G75) );
  XOR2_X1 U772 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n721) );
  XNOR2_X1 U773 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n720) );
  XNOR2_X1 U774 ( .A(n721), .B(n720), .ZN(n722) );
  XOR2_X1 U775 ( .A(n723), .B(n722), .Z(n726) );
  NAND2_X1 U776 ( .A1(n724), .A2(G469), .ZN(n725) );
  XNOR2_X1 U777 ( .A(n726), .B(n725), .ZN(n728) );
  INV_X1 U778 ( .A(n727), .ZN(n732) );
  NOR2_X1 U779 ( .A1(n728), .A2(n732), .ZN(G54) );
  NAND2_X1 U780 ( .A1(G217), .A2(n724), .ZN(n729) );
  XNOR2_X1 U781 ( .A(n729), .B(n730), .ZN(n731) );
  NOR2_X1 U782 ( .A1(n732), .A2(n731), .ZN(G66) );
  XOR2_X1 U783 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n734) );
  NAND2_X1 U784 ( .A1(G224), .A2(G953), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n734), .B(n733), .ZN(n735) );
  NAND2_X1 U786 ( .A1(n735), .A2(G898), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U788 ( .A1(n739), .A2(n738), .ZN(n744) );
  XNOR2_X1 U789 ( .A(n740), .B(G101), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U791 ( .A(n744), .B(n743), .Z(G69) );
  XOR2_X1 U792 ( .A(n746), .B(n745), .Z(n747) );
  XOR2_X1 U793 ( .A(KEYINPUT126), .B(n747), .Z(n751) );
  XOR2_X1 U794 ( .A(n751), .B(n748), .Z(n750) );
  NAND2_X1 U795 ( .A1(n750), .A2(n749), .ZN(n755) );
  XNOR2_X1 U796 ( .A(G227), .B(n751), .ZN(n752) );
  NAND2_X1 U797 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U798 ( .A1(n753), .A2(G953), .ZN(n754) );
  NAND2_X1 U799 ( .A1(n755), .A2(n754), .ZN(G72) );
  XOR2_X1 U800 ( .A(n756), .B(G119), .Z(G21) );
  XNOR2_X1 U801 ( .A(G143), .B(KEYINPUT111), .ZN(n758) );
  XNOR2_X1 U802 ( .A(n758), .B(n757), .ZN(G45) );
  XNOR2_X1 U803 ( .A(n759), .B(G131), .ZN(G33) );
  XOR2_X1 U804 ( .A(G137), .B(n760), .Z(n761) );
  XNOR2_X1 U805 ( .A(KEYINPUT127), .B(n761), .ZN(G39) );
endmodule

