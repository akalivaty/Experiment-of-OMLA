//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  INV_X1    g003(.A(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT90), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n202), .A2(KEYINPUT90), .A3(G1gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n202), .A2(G1gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(KEYINPUT91), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n212), .A2(new_n204), .A3(new_n207), .A4(new_n208), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT21), .ZN(new_n217));
  NAND2_X1  g016(.A1(G71gat), .A2(G78gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT95), .ZN(new_n221));
  INV_X1    g020(.A(G64gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G57gat), .ZN(new_n223));
  INV_X1    g022(.A(G57gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G64gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT95), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n218), .A2(new_n227), .A3(new_n219), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G71gat), .B(G78gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n221), .A2(new_n226), .A3(new_n230), .A4(new_n228), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n216), .B1(new_n217), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT96), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G127gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n217), .ZN(new_n238));
  XNOR2_X1  g037(.A(G183gat), .B(G211gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G231gat), .A2(G233gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G127gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n236), .B(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(new_n242), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(G155gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n250), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(new_n244), .B2(new_n247), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G134gat), .B(G162gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT17), .ZN(new_n257));
  XNOR2_X1  g056(.A(G43gat), .B(G50gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT14), .ZN(new_n259));
  INV_X1    g058(.A(G29gat), .ZN(new_n260));
  INV_X1    g059(.A(G36gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(KEYINPUT88), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G29gat), .A2(G36gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n263), .B1(new_n262), .B2(KEYINPUT88), .ZN(new_n267));
  OAI211_X1 g066(.A(KEYINPUT15), .B(new_n258), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n258), .A2(KEYINPUT15), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n258), .A2(KEYINPUT15), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n262), .A2(new_n263), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n265), .A4(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT89), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n268), .B2(new_n272), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n257), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OR2_X1    g076(.A1(G85gat), .A2(G92gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(G99gat), .A2(G106gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT8), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT7), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n281), .B1(G85gat), .B2(G92gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(G85gat), .A2(G92gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT7), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n278), .B(new_n280), .C1(new_n282), .C2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G99gat), .B(G106gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(KEYINPUT7), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n281), .A2(G85gat), .A3(G92gat), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n289), .A2(new_n290), .B1(KEYINPUT8), .B2(new_n279), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n286), .A3(new_n278), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n268), .A2(new_n272), .A3(KEYINPUT17), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AND3_X1   g094(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n276), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n274), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n289), .A2(new_n290), .ZN(new_n299));
  AND4_X1   g098(.A1(new_n286), .A2(new_n299), .A3(new_n278), .A4(new_n280), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n286), .B1(new_n291), .B2(new_n278), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n296), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(G190gat), .B(G218gat), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT97), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n295), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n309), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n295), .A2(new_n303), .A3(new_n311), .A4(new_n307), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n256), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n256), .A3(new_n312), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n314), .A2(KEYINPUT97), .A3(new_n304), .A4(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n315), .ZN(new_n317));
  OAI22_X1  g116(.A1(new_n317), .A2(new_n313), .B1(new_n306), .B2(new_n305), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n254), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G78gat), .B(G106gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT31), .B(G50gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326));
  INV_X1    g125(.A(G211gat), .ZN(new_n327));
  INV_X1    g126(.A(G218gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G211gat), .B(G218gat), .Z(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n334));
  INV_X1    g133(.A(G141gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(G148gat), .ZN(new_n336));
  INV_X1    g135(.A(G148gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n336), .B(new_n338), .C1(G141gat), .C2(new_n337), .ZN(new_n339));
  XNOR2_X1  g138(.A(G155gat), .B(G162gat), .ZN(new_n340));
  INV_X1    g139(.A(G155gat), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT2), .B1(new_n341), .B2(KEYINPUT77), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  INV_X1    g143(.A(new_n340), .ZN(new_n345));
  XNOR2_X1  g144(.A(G141gat), .B(G148gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(KEYINPUT2), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G22gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n343), .A2(new_n347), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT3), .B1(new_n332), .B2(new_n333), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n350), .B(new_n351), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n332), .A2(new_n333), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n353), .B1(new_n356), .B2(new_n344), .ZN(new_n357));
  OAI21_X1  g156(.A(G22gat), .B1(new_n357), .B2(new_n349), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n355), .A2(new_n358), .A3(G228gat), .A4(G233gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n355), .A2(new_n358), .B1(G228gat), .B2(G233gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n324), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(KEYINPUT81), .B(new_n324), .C1(new_n360), .C2(new_n361), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n361), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(new_n323), .A3(new_n359), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT82), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n367), .A2(new_n370), .A3(new_n323), .A4(new_n359), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G169gat), .ZN(new_n375));
  INV_X1    g174(.A(G176gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT23), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT23), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(G169gat), .B2(G176gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT24), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G190gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT65), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT65), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G190gat), .ZN(new_n388));
  AOI21_X1  g187(.A(G183gat), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n381), .B(KEYINPUT25), .C1(new_n384), .C2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT25), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n382), .A2(new_n383), .ZN(new_n392));
  NOR2_X1   g191(.A1(G183gat), .A2(G190gat), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT67), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n399), .A2(new_n375), .A3(new_n376), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT26), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT26), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n399), .A2(new_n402), .A3(new_n375), .A4(new_n376), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n380), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n388), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT27), .B(G183gat), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT28), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT28), .B1(new_n405), .B2(new_n406), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n382), .B(new_n404), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n398), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT73), .ZN(new_n411));
  NAND2_X1  g210(.A1(G226gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT73), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT74), .ZN(new_n417));
  INV_X1    g216(.A(new_n409), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT66), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n398), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n390), .A2(new_n397), .A3(KEYINPUT66), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n412), .B1(new_n422), .B2(KEYINPUT29), .ZN(new_n423));
  INV_X1    g222(.A(new_n332), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT74), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n411), .A2(new_n425), .A3(new_n413), .A4(new_n415), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n417), .A2(new_n423), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n413), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n411), .A2(new_n333), .A3(new_n412), .A4(new_n415), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n332), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G8gat), .B(G36gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(G64gat), .B(G92gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT75), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT75), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n431), .A2(new_n439), .A3(new_n435), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G127gat), .B(G134gat), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT68), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT1), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(G113gat), .B(G120gat), .Z(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n444), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n446), .B(new_n444), .C1(new_n443), .C2(new_n442), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(KEYINPUT4), .A3(new_n353), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n352), .A2(KEYINPUT3), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n450), .A3(new_n348), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n448), .A2(new_n347), .A3(new_n343), .A4(new_n449), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT4), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G225gat), .A2(G233gat), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT4), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n452), .A2(new_n454), .A3(new_n457), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n450), .A2(new_n352), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n455), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n450), .A2(KEYINPUT78), .A3(new_n352), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n459), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(new_n466), .A3(KEYINPUT5), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n452), .A2(new_n454), .A3(new_n457), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n459), .A2(KEYINPUT5), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G1gat), .B(G29gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(G85gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT0), .B(G57gat), .ZN(new_n474));
  XOR2_X1   g273(.A(new_n473), .B(new_n474), .Z(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT79), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n471), .A2(new_n476), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT79), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n467), .A2(new_n470), .A3(new_n480), .A4(new_n475), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n477), .A2(new_n478), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n476), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n431), .A2(KEYINPUT30), .A3(new_n435), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n431), .A2(new_n435), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n441), .A2(new_n484), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT80), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n488), .A2(new_n489), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n374), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n441), .A2(new_n485), .A3(new_n487), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n464), .A2(new_n465), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n458), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT39), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n468), .A2(new_n458), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(KEYINPUT83), .A3(KEYINPUT39), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n499), .A2(KEYINPUT39), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n475), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT40), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n467), .A2(new_n470), .A3(KEYINPUT84), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT84), .B1(new_n467), .B2(new_n470), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n476), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n493), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n427), .A2(KEYINPUT37), .A3(new_n430), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n434), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n431), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n510), .B1(new_n509), .B2(new_n434), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT38), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n483), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n507), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n439), .B1(new_n431), .B2(new_n435), .ZN(new_n520));
  AOI211_X1 g319(.A(KEYINPUT75), .B(new_n434), .C1(new_n427), .C2(new_n430), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n417), .A2(new_n423), .A3(new_n426), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n512), .B1(new_n523), .B2(new_n332), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n428), .A2(new_n429), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n524), .B1(new_n332), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT38), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n526), .A2(new_n527), .A3(new_n434), .A4(new_n513), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n516), .A2(new_n519), .A3(new_n522), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n529), .A3(new_n373), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT69), .B1(new_n422), .B2(new_n451), .ZN(new_n531));
  INV_X1    g330(.A(new_n421), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT66), .B1(new_n390), .B2(new_n397), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n409), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT69), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(new_n450), .ZN(new_n536));
  NAND2_X1  g335(.A1(G227gat), .A2(G233gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT64), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n422), .A2(new_n451), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n531), .A2(new_n536), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT34), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT32), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n531), .A2(new_n536), .A3(new_n540), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(new_n545), .B2(new_n538), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n538), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT33), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G15gat), .B(G43gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G71gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G99gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n546), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  AND4_X1   g354(.A1(KEYINPUT32), .A2(new_n547), .A3(KEYINPUT33), .A4(new_n554), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n543), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n547), .A2(KEYINPUT32), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT33), .B1(new_n545), .B2(new_n538), .ZN(new_n559));
  INV_X1    g358(.A(new_n554), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n549), .A2(new_n546), .A3(new_n554), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n562), .A3(new_n542), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n557), .A2(KEYINPUT36), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n557), .A2(new_n566), .A3(new_n563), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT36), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT72), .A4(new_n542), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT71), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n565), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n564), .A2(KEYINPUT71), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n492), .B(new_n530), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n567), .A2(new_n569), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT86), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n567), .A2(KEYINPUT86), .A3(new_n569), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n493), .A2(KEYINPUT35), .A3(new_n519), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n577), .A2(new_n373), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n486), .B1(new_n522), .B2(new_n438), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n581), .A2(KEYINPUT80), .A3(new_n484), .A4(new_n485), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n488), .A2(new_n489), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n373), .A2(new_n563), .A3(new_n557), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT35), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n320), .B1(new_n574), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n216), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n214), .A2(KEYINPUT92), .A3(new_n215), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n277), .A2(new_n590), .A3(new_n294), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n298), .A2(new_n215), .A3(new_n214), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT18), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n592), .A2(new_n597), .A3(new_n593), .A4(new_n594), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n216), .A2(new_n297), .A3(new_n274), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT93), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT93), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n216), .A2(new_n297), .A3(new_n602), .A4(new_n274), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n601), .A2(new_n594), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n593), .B(KEYINPUT13), .Z(new_n605));
  AOI21_X1  g404(.A(KEYINPUT94), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n604), .A2(KEYINPUT94), .A3(new_n605), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n599), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G169gat), .B(G197gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n599), .B(new_n614), .C1(new_n606), .C2(new_n607), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G230gat), .ZN(new_n620));
  INV_X1    g419(.A(G233gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n232), .A2(new_n288), .A3(new_n233), .A4(new_n292), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n218), .A2(new_n227), .A3(new_n219), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n227), .B1(new_n218), .B2(new_n219), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n230), .B1(new_n629), .B2(new_n226), .ZN(new_n630));
  INV_X1    g429(.A(new_n233), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n632), .A2(new_n302), .A3(KEYINPUT99), .A4(KEYINPUT10), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n234), .A2(new_n293), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT98), .B(KEYINPUT10), .Z(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n624), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n622), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n622), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n635), .A2(new_n624), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT100), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n647), .A2(KEYINPUT101), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n642), .A2(new_n645), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(KEYINPUT101), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n619), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n588), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n484), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  INV_X1    g456(.A(KEYINPUT102), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n493), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT16), .B(G8gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(KEYINPUT42), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(G8gat), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(KEYINPUT42), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(G1325gat));
  INV_X1    g464(.A(new_n577), .ZN(new_n666));
  INV_X1    g465(.A(new_n578), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(G15gat), .B1(new_n654), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n570), .A2(new_n571), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n564), .ZN(new_n671));
  INV_X1    g470(.A(new_n573), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n675), .A2(G15gat), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n669), .B1(new_n654), .B2(new_n676), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n654), .A2(new_n374), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(new_n351), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n373), .B1(new_n582), .B2(new_n583), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n508), .A2(new_n529), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n373), .B2(new_n684), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n685), .A2(new_n673), .B1(new_n586), .B2(new_n580), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n682), .B1(new_n686), .B2(new_n319), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n574), .A2(new_n587), .ZN(new_n688));
  INV_X1    g487(.A(new_n319), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(KEYINPUT44), .A3(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n254), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n653), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G29gat), .B1(new_n695), .B2(new_n484), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n686), .A2(new_n319), .A3(new_n693), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(new_n260), .A3(new_n655), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n699), .B2(new_n701), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n696), .B1(new_n702), .B2(new_n703), .ZN(G1328gat));
  NAND3_X1  g503(.A1(new_n697), .A2(new_n261), .A3(new_n493), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT46), .Z(new_n706));
  INV_X1    g505(.A(new_n493), .ZN(new_n707));
  OAI21_X1  g506(.A(G36gat), .B1(new_n695), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1329gat));
  OAI21_X1  g508(.A(G43gat), .B1(new_n695), .B2(new_n673), .ZN(new_n710));
  INV_X1    g509(.A(G43gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n697), .A2(new_n711), .A3(new_n668), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n710), .A2(new_n712), .A3(KEYINPUT47), .ZN(new_n713));
  INV_X1    g512(.A(new_n712), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n691), .A2(new_n675), .A3(new_n694), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(G43gat), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n713), .B1(new_n716), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  INV_X1    g517(.A(G50gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n697), .A2(new_n719), .A3(new_n374), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n718), .B1(new_n720), .B2(KEYINPUT107), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n687), .A2(new_n374), .A3(new_n694), .A4(new_n690), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G50gat), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n721), .B(new_n723), .C1(KEYINPUT107), .C2(new_n720), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n723), .A2(new_n720), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(G1331gat));
  INV_X1    g526(.A(new_n320), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n688), .A2(new_n728), .A3(new_n619), .A4(new_n652), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n484), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(new_n224), .ZN(G1332gat));
  NAND2_X1  g530(.A1(new_n729), .A2(KEYINPUT108), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n588), .A2(new_n733), .A3(new_n619), .A4(new_n652), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n707), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n736));
  NAND2_X1  g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n732), .A2(new_n734), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(new_n493), .A3(new_n737), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT109), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n740), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n742), .A2(new_n747), .ZN(G1333gat));
  XNOR2_X1  g547(.A(new_n673), .B(KEYINPUT103), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n732), .B2(new_n734), .ZN(new_n750));
  INV_X1    g549(.A(G71gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n668), .A2(new_n751), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n750), .A2(new_n751), .B1(new_n729), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n743), .A2(new_n374), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g556(.A1(new_n254), .A2(new_n618), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n687), .A2(new_n652), .A3(new_n690), .A4(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(G85gat), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n759), .A2(new_n760), .A3(new_n484), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n686), .B2(new_n319), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n688), .A2(KEYINPUT110), .A3(new_n689), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(new_n758), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT51), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n763), .A2(new_n767), .A3(new_n758), .A4(new_n764), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n766), .A2(new_n655), .A3(new_n652), .A4(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n761), .B1(new_n769), .B2(new_n760), .ZN(G1336gat));
  NOR2_X1   g569(.A1(new_n707), .A2(G92gat), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n766), .A2(new_n652), .A3(new_n768), .A4(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  OAI21_X1  g572(.A(G92gat), .B1(new_n759), .B2(new_n707), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n767), .A2(KEYINPUT111), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n765), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n776), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n763), .A2(new_n758), .A3(new_n764), .A4(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n777), .A2(new_n652), .A3(new_n771), .A4(new_n779), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n774), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n775), .B1(new_n781), .B2(new_n773), .ZN(G1337gat));
  INV_X1    g581(.A(new_n652), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n666), .A2(new_n667), .A3(G99gat), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT112), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n768), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G99gat), .B1(new_n759), .B2(new_n749), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1338gat));
  NOR2_X1   g587(.A1(new_n373), .A2(G106gat), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n766), .A2(new_n652), .A3(new_n768), .A4(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  OAI21_X1  g590(.A(G106gat), .B1(new_n759), .B2(new_n373), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n652), .A3(new_n779), .A4(new_n789), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(new_n792), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n795), .B2(new_n791), .ZN(G1339gat));
  NAND3_X1  g595(.A1(new_n634), .A2(new_n622), .A3(new_n637), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n639), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n798));
  AOI211_X1 g597(.A(KEYINPUT54), .B(new_n622), .C1(new_n634), .C2(new_n637), .ZN(new_n799));
  INV_X1    g598(.A(new_n645), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(KEYINPUT113), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n634), .A2(new_n637), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n804), .A3(new_n640), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n802), .B1(new_n805), .B2(new_n645), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n798), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n649), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(KEYINPUT55), .B(new_n798), .C1(new_n801), .C2(new_n806), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(KEYINPUT114), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT54), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n638), .ZN(new_n814));
  OAI21_X1  g613(.A(KEYINPUT113), .B1(new_n799), .B2(new_n800), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n805), .A2(new_n802), .A3(new_n645), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n812), .B1(new_n817), .B2(KEYINPUT55), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n809), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n604), .A2(new_n605), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n593), .B1(new_n592), .B2(new_n594), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n613), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n617), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n689), .A2(new_n820), .A3(new_n825), .ZN(new_n826));
  AOI22_X1  g625(.A1(new_n820), .A2(new_n618), .B1(new_n652), .B2(new_n825), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT115), .B(new_n826), .C1(new_n827), .C2(new_n689), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n810), .A2(KEYINPUT114), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n817), .A2(new_n812), .A3(KEYINPUT55), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n618), .A2(new_n809), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n825), .A2(new_n652), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n689), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n319), .A2(new_n819), .A3(new_n824), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n829), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n828), .A2(new_n837), .A3(new_n692), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n254), .A2(new_n319), .A3(new_n619), .A4(new_n783), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n666), .A2(new_n667), .A3(new_n374), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n493), .A2(new_n484), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n619), .ZN(new_n845));
  INV_X1    g644(.A(new_n839), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n835), .A2(new_n836), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n254), .B1(new_n847), .B2(KEYINPUT115), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(new_n837), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n484), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n707), .A3(new_n584), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n619), .A2(G113gat), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT116), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n845), .B1(new_n851), .B2(new_n853), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n844), .B2(new_n783), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n783), .A2(G120gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n851), .B2(new_n856), .ZN(G1341gat));
  NOR3_X1   g656(.A1(new_n844), .A2(new_n245), .A3(new_n692), .ZN(new_n858));
  INV_X1    g657(.A(new_n851), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n254), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n858), .B1(new_n860), .B2(new_n245), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n862), .A3(new_n689), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  INV_X1    g665(.A(new_n844), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT117), .B(new_n862), .C1(new_n867), .C2(new_n689), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n689), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(G134gat), .ZN(new_n871));
  OAI22_X1  g670(.A1(new_n865), .A2(new_n866), .B1(new_n868), .B2(new_n871), .ZN(G1343gat));
  NAND2_X1  g671(.A1(new_n673), .A2(new_n843), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n819), .A2(KEYINPUT118), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n832), .A2(new_n875), .A3(new_n809), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n874), .A2(new_n618), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n689), .B1(new_n877), .B2(new_n834), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n692), .B1(new_n878), .B2(new_n836), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n839), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n373), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT119), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  INV_X1    g683(.A(new_n882), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n884), .B(new_n885), .C1(new_n879), .C2(new_n839), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n840), .A2(new_n374), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n881), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n873), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n335), .B1(new_n890), .B2(new_n618), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n675), .A2(new_n373), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n892), .A2(new_n850), .A3(new_n707), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n893), .A2(new_n335), .A3(new_n618), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT58), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n886), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n882), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n884), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n889), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n873), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n618), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G141gat), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n893), .A2(new_n335), .A3(new_n618), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n895), .A2(new_n905), .ZN(G1344gat));
  NAND4_X1  g705(.A1(new_n893), .A2(KEYINPUT120), .A3(new_n337), .A4(new_n652), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n850), .A3(new_n337), .A4(new_n707), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(new_n783), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n839), .B(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT57), .B1(new_n913), .B2(new_n879), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n914), .A2(new_n374), .B1(new_n888), .B2(KEYINPUT57), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n783), .B1(new_n873), .B2(new_n916), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n915), .B(new_n917), .C1(new_n916), .C2(new_n873), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n337), .B1(new_n890), .B2(new_n652), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n911), .B(new_n919), .C1(KEYINPUT59), .C2(new_n920), .ZN(G1345gat));
  XOR2_X1   g720(.A(KEYINPUT77), .B(G155gat), .Z(new_n922));
  AOI21_X1  g721(.A(new_n922), .B1(new_n893), .B2(new_n254), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n254), .A2(new_n922), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n890), .B2(new_n924), .ZN(G1346gat));
  INV_X1    g724(.A(G162gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n893), .A2(new_n926), .A3(new_n689), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n890), .A2(new_n689), .ZN(new_n931));
  OAI22_X1  g730(.A1(new_n929), .A2(new_n930), .B1(new_n926), .B2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n707), .A2(new_n655), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n842), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G169gat), .B1(new_n934), .B2(new_n619), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT124), .B1(new_n840), .B2(new_n484), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  AOI211_X1 g736(.A(new_n937), .B(new_n655), .C1(new_n838), .C2(new_n839), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n493), .B(new_n584), .C1(new_n936), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n618), .A2(new_n375), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(G1348gat));
  NOR3_X1   g740(.A1(new_n934), .A2(new_n376), .A3(new_n783), .ZN(new_n942));
  INV_X1    g741(.A(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n652), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n944), .B2(new_n376), .ZN(G1349gat));
  NAND3_X1  g744(.A1(new_n842), .A2(new_n254), .A3(new_n933), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G183gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n254), .A2(new_n406), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n939), .B2(new_n948), .ZN(new_n949));
  OR2_X1    g748(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n950));
  NAND2_X1  g749(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n937), .B1(new_n849), .B2(new_n655), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n840), .A2(KEYINPUT124), .A3(new_n484), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n948), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n955), .A2(new_n493), .A3(new_n584), .A4(new_n956), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n957), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n947), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n952), .A2(new_n958), .ZN(G1350gat));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n405), .A3(new_n689), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n840), .A2(new_n841), .A3(new_n689), .A4(new_n933), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G190gat), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n964), .B1(new_n963), .B2(new_n965), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n960), .B1(new_n966), .B2(new_n967), .ZN(G1351gat));
  NAND2_X1  g767(.A1(new_n913), .A2(new_n879), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n969), .A2(new_n881), .A3(new_n374), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n888), .A2(KEYINPUT57), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n970), .A2(new_n971), .A3(new_n749), .A4(new_n933), .ZN(new_n972));
  OAI21_X1  g771(.A(G197gat), .B1(new_n972), .B2(new_n619), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n749), .A2(new_n374), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n974), .B1(new_n953), .B2(new_n954), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n493), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n619), .A2(G197gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(G1352gat));
  AND3_X1   g777(.A1(new_n970), .A2(new_n971), .A3(new_n933), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n979), .A2(KEYINPUT127), .A3(new_n652), .A4(new_n749), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n981), .B1(new_n972), .B2(new_n783), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n980), .A2(G204gat), .A3(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(G204gat), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n975), .A2(new_n984), .A3(new_n493), .A4(new_n652), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n983), .A2(new_n986), .A3(new_n987), .ZN(G1353gat));
  INV_X1    g787(.A(new_n976), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n989), .A2(new_n327), .A3(new_n254), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n915), .A2(new_n254), .A3(new_n749), .A4(new_n933), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  INV_X1    g791(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(G1354gat));
  NOR3_X1   g794(.A1(new_n972), .A2(new_n328), .A3(new_n319), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n989), .A2(new_n689), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n996), .B1(new_n997), .B2(new_n328), .ZN(G1355gat));
endmodule


