//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n560, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n616, new_n618, new_n619,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT69), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(KEYINPUT70), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT3), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT71), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n462), .A2(G137), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n460), .A2(KEYINPUT70), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n458), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n465), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n474), .A2(new_n481), .ZN(G160));
  AOI22_X1  g057(.A1(new_n471), .A2(KEYINPUT3), .B1(new_n463), .B2(new_n466), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(new_n475), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n475), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  AND2_X1   g068(.A1(KEYINPUT4), .A2(G138), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n462), .A2(new_n475), .A3(new_n467), .A4(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n475), .A2(G102), .A3(G2104), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n476), .A2(new_n477), .A3(G138), .A4(new_n475), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n483), .B2(G126), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n495), .B(new_n499), .C1(new_n502), .C2(new_n475), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G62), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT73), .A3(G62), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT74), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n512), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(KEYINPUT6), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(KEYINPUT72), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n524), .A2(G88), .A3(new_n513), .A4(new_n525), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n524), .A2(G50), .A3(G543), .A4(new_n525), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n518), .A2(new_n528), .ZN(G166));
  AOI22_X1  g104(.A1(new_n521), .A2(new_n523), .B1(KEYINPUT6), .B2(new_n520), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n534), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n524), .A2(new_n513), .A3(new_n525), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n535), .A2(new_n537), .A3(new_n540), .A4(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n539), .A2(G90), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n520), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n524), .A2(G543), .A3(new_n525), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G52), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n510), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n547), .A2(G43), .B1(new_n553), .B2(G651), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n539), .A2(G81), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  XOR2_X1   g134(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n560));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(new_n539), .A2(G91), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n547), .A2(new_n566), .A3(G53), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n566), .B1(new_n547), .B2(G53), .ZN(new_n568));
  OAI221_X1 g143(.A(new_n564), .B1(new_n520), .B2(new_n565), .C1(new_n567), .C2(new_n568), .ZN(G299));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n518), .A2(new_n570), .A3(new_n528), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n570), .B1(new_n518), .B2(new_n528), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n571), .A2(new_n572), .ZN(G303));
  NAND2_X1  g148(.A1(new_n539), .A2(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n547), .A2(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n538), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n530), .A2(KEYINPUT78), .A3(G86), .A4(new_n513), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n510), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n547), .A2(G48), .B1(new_n585), .B2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n520), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT79), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  OAI221_X1 g167(.A(new_n590), .B1(new_n591), .B2(new_n531), .C1(new_n592), .C2(new_n538), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(G66), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(G66), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n513), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G79), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n506), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(KEYINPUT81), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(KEYINPUT81), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n601), .A2(G651), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n539), .A2(KEYINPUT10), .A3(G92), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n538), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n604), .A2(new_n607), .B1(G54), .B2(new_n547), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT82), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n594), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n594), .B1(new_n611), .B2(G868), .ZN(G321));
  MUX2_X1   g188(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g189(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g190(.A(KEYINPUT83), .B(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n611), .B1(G860), .B2(new_n616), .ZN(G148));
  NAND2_X1  g192(.A1(new_n611), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g195(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n621));
  XNOR2_X1  g196(.A(G323), .B(new_n621), .ZN(G282));
  NAND2_X1  g197(.A1(new_n485), .A2(G123), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n488), .A2(G135), .ZN(new_n624));
  NOR2_X1   g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT86), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n472), .A2(new_n478), .A3(new_n475), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT85), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n629), .A2(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XOR2_X1   g212(.A(G2443), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT88), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT15), .B(G2435), .Z(new_n646));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n647));
  AOI22_X1  g222(.A1(new_n645), .A2(new_n646), .B1(KEYINPUT87), .B2(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(KEYINPUT87), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n648), .B(new_n649), .C1(new_n646), .C2(new_n645), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n641), .B(new_n650), .Z(new_n651));
  AND2_X1   g226(.A1(new_n651), .A2(G14), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2067), .B(G2678), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT17), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n661), .B(new_n662), .C1(new_n660), .C2(new_n656), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(KEYINPUT90), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(KEYINPUT90), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n676), .A2(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n667), .A2(new_n668), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(KEYINPUT20), .ZN(new_n680));
  INV_X1    g255(.A(new_n669), .ZN(new_n681));
  OR3_X1    g256(.A1(new_n673), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g257(.A1(new_n677), .A2(new_n679), .A3(new_n680), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1986), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1991), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n685), .B(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n690), .A2(G22), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G166), .B2(new_n690), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(KEYINPUT94), .ZN(new_n694));
  INV_X1    g269(.A(G1971), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n691), .A2(KEYINPUT94), .ZN(new_n696));
  AND3_X1   g271(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n695), .B1(new_n694), .B2(new_n696), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT34), .ZN(new_n700));
  MUX2_X1   g275(.A(G6), .B(G305), .S(G16), .Z(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(G288), .A2(G16), .ZN(new_n704));
  INV_X1    g279(.A(G23), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(G16), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(KEYINPUT33), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n704), .A2(new_n710), .A3(new_n707), .ZN(new_n711));
  AOI21_X1  g286(.A(G1976), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n710), .B1(new_n704), .B2(new_n707), .ZN(new_n713));
  AOI211_X1 g288(.A(KEYINPUT33), .B(new_n706), .C1(G288), .C2(G16), .ZN(new_n714));
  INV_X1    g289(.A(G1976), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n699), .A2(new_n700), .A3(new_n703), .A4(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n690), .A2(G24), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G290), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT93), .B(G1986), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n483), .A2(G119), .A3(G2105), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n483), .A2(G131), .A3(new_n475), .ZN(new_n725));
  OR2_X1    g300(.A1(G95), .A2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(KEYINPUT91), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n724), .A2(new_n725), .A3(new_n730), .A4(new_n727), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n723), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G25), .A2(G29), .ZN(new_n733));
  OR3_X1    g308(.A1(new_n732), .A2(KEYINPUT92), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT35), .B(G1991), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT92), .B1(new_n732), .B2(new_n733), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n735), .B1(new_n734), .B2(new_n736), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n718), .A2(new_n722), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(KEYINPUT95), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT95), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n718), .A2(new_n742), .A3(new_n739), .A4(new_n722), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT96), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n699), .A2(new_n703), .A3(new_n717), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT34), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n723), .A2(G26), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n485), .A2(G128), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n488), .A2(G140), .ZN(new_n753));
  OR2_X1    g328(.A1(G104), .A2(G2105), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT98), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n460), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n756), .B1(new_n755), .B2(new_n754), .C1(G116), .C2(new_n475), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n752), .A2(new_n753), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n751), .B1(new_n759), .B2(new_n723), .ZN(new_n760));
  MUX2_X1   g335(.A(new_n751), .B(new_n760), .S(KEYINPUT28), .Z(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT99), .B(G2067), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT36), .A4(new_n747), .ZN(new_n764));
  OR2_X1    g339(.A1(G16), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G286), .B2(new_n690), .ZN(new_n766));
  INV_X1    g341(.A(G1966), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT102), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n723), .A2(G35), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G162), .B2(new_n723), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(KEYINPUT29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(KEYINPUT29), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G2090), .ZN(new_n776));
  INV_X1    g351(.A(G2090), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n773), .A2(new_n777), .A3(new_n774), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n770), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT24), .A2(G34), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT24), .A2(G34), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n780), .A2(new_n723), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G160), .B2(new_n723), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G2084), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT101), .Z(new_n785));
  NAND2_X1  g360(.A1(G171), .A2(G16), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G5), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G1961), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OR2_X1    g364(.A1(G29), .A2(G32), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n485), .A2(G129), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n488), .A2(G141), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT26), .Z(new_n794));
  NAND3_X1  g369(.A1(new_n472), .A2(G105), .A3(new_n475), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n791), .A2(new_n792), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n790), .B1(new_n796), .B2(new_n723), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT27), .B(G1996), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n789), .B(new_n799), .C1(G2084), .C2(new_n783), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n723), .A2(G27), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G164), .B2(new_n723), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2078), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n690), .A2(G19), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n556), .B2(new_n690), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT97), .B(G1341), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  OR4_X1    g382(.A1(new_n785), .A2(new_n800), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n779), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n690), .A2(G4), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n611), .B2(new_n690), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n811), .A2(G1348), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n766), .A2(new_n767), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n788), .B2(new_n787), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT31), .B(G11), .Z(new_n815));
  INV_X1    g390(.A(G28), .ZN(new_n816));
  AOI21_X1  g391(.A(G29), .B1(new_n816), .B2(KEYINPUT30), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(KEYINPUT30), .B2(new_n816), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n818), .B1(new_n723), .B2(new_n627), .C1(new_n797), .C2(new_n798), .ZN(new_n819));
  OR3_X1    g394(.A1(new_n814), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n811), .A2(G1348), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n812), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT25), .Z(new_n824));
  AOI22_X1  g399(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n825));
  INV_X1    g400(.A(G139), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n824), .B1(new_n825), .B2(new_n475), .C1(new_n487), .C2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT100), .ZN(new_n828));
  MUX2_X1   g403(.A(G33), .B(new_n828), .S(G29), .Z(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(G2072), .Z(new_n830));
  INV_X1    g405(.A(KEYINPUT23), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n690), .A2(G20), .ZN(new_n832));
  AOI211_X1 g407(.A(new_n831), .B(new_n832), .C1(G299), .C2(G16), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n831), .B2(new_n832), .ZN(new_n834));
  INV_X1    g409(.A(G1956), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n809), .A2(new_n822), .A3(new_n830), .A4(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n750), .A2(new_n763), .A3(new_n764), .A4(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(G311));
  NAND2_X1  g415(.A1(new_n839), .A2(KEYINPUT103), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n837), .B1(new_n748), .B2(new_n749), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n842), .A2(new_n843), .A3(new_n763), .A4(new_n764), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n844), .ZN(G150));
  NAND2_X1  g420(.A1(new_n539), .A2(G93), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n547), .A2(G55), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n846), .B(new_n847), .C1(new_n520), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n611), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n556), .B(new_n849), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT39), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n853), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n851), .B1(new_n856), .B2(G860), .ZN(G145));
  XNOR2_X1  g432(.A(new_n627), .B(G160), .ZN(new_n858));
  INV_X1    g433(.A(G142), .ZN(new_n859));
  NOR2_X1   g434(.A1(G106), .A2(G2105), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(new_n475), .B2(G118), .ZN(new_n861));
  OAI22_X1  g436(.A1(new_n487), .A2(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(G130), .B2(new_n485), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n492), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n858), .B(new_n864), .Z(new_n865));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n462), .A2(G126), .A3(new_n467), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n500), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(G2105), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n495), .A2(new_n499), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n475), .B1(new_n867), .B2(new_n500), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n495), .A2(new_n499), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT104), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n759), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n871), .A2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(new_n758), .ZN(new_n877));
  INV_X1    g452(.A(new_n796), .ZN(new_n878));
  OR3_X1    g453(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n828), .B(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n878), .B1(new_n875), .B2(new_n877), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n828), .A2(new_n880), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n879), .B2(new_n882), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n631), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n884), .A2(new_n886), .A3(new_n631), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n888), .A2(new_n889), .A3(new_n728), .ZN(new_n890));
  INV_X1    g465(.A(new_n728), .ZN(new_n891));
  OR3_X1    g466(.A1(new_n884), .A2(new_n631), .A3(new_n886), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n892), .B2(new_n887), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n865), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n728), .B1(new_n888), .B2(new_n889), .ZN(new_n895));
  INV_X1    g470(.A(new_n865), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n887), .A3(new_n891), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT40), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n894), .A2(new_n898), .A3(new_n902), .A4(new_n899), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(G395));
  NOR2_X1   g479(.A1(new_n849), .A2(G868), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n518), .A2(new_n528), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(G288), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(G305), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n908), .B(G290), .Z(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT42), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(KEYINPUT106), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(KEYINPUT106), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n618), .B(new_n854), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n609), .A2(G299), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n609), .A2(G299), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT41), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n916), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n913), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n911), .A2(new_n912), .A3(new_n925), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n910), .B(KEYINPUT106), .C1(new_n922), .C2(new_n924), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n905), .B1(new_n928), .B2(G868), .ZN(G295));
  AOI21_X1  g504(.A(new_n905), .B1(new_n928), .B2(G868), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n854), .A2(KEYINPUT107), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n854), .A2(KEYINPUT107), .ZN(new_n933));
  XNOR2_X1  g508(.A(G286), .B(G301), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n932), .B2(new_n933), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n923), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n854), .B(KEYINPUT107), .ZN(new_n939));
  INV_X1    g514(.A(new_n934), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(new_n920), .A3(new_n935), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n908), .B(G290), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n899), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n938), .B2(new_n942), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n931), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n945), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n917), .A2(new_n949), .A3(new_n919), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n919), .A2(new_n949), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n941), .A2(new_n950), .A3(new_n935), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n938), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT109), .B1(new_n953), .B2(new_n909), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  AOI211_X1 g530(.A(new_n955), .B(new_n943), .C1(new_n938), .C2(new_n952), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n948), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n947), .B1(new_n957), .B2(new_n931), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT44), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT43), .B1(new_n945), .B2(new_n946), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n957), .B2(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n871), .B2(new_n874), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n481), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n468), .A2(new_n473), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n969), .B(G40), .C1(new_n970), .C2(G2105), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  OR3_X1    g548(.A1(new_n973), .A2(G1986), .A3(G290), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(G1986), .A3(G290), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT110), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT111), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n973), .B2(G1996), .ZN(new_n979));
  INV_X1    g554(.A(G1996), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n972), .A2(KEYINPUT111), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G2067), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n758), .B(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n980), .B2(new_n878), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n982), .A2(new_n878), .B1(new_n972), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n728), .B(new_n735), .Z(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(new_n973), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n977), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G2084), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n503), .A2(new_n991), .A3(new_n965), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n965), .B1(new_n872), .B2(new_n873), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT50), .ZN(new_n994));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n474), .A2(new_n995), .A3(new_n481), .ZN(new_n996));
  AND4_X1   g571(.A1(new_n990), .A2(new_n992), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT45), .B1(new_n503), .B2(new_n965), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(new_n999), .B2(new_n971), .ZN(new_n1000));
  INV_X1    g575(.A(new_n993), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT45), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT117), .B(new_n996), .C1(new_n1001), .C2(KEYINPUT45), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n997), .B1(new_n1004), .B2(new_n767), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT51), .B1(new_n1005), .B2(G168), .ZN(new_n1006));
  INV_X1    g581(.A(G8), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n1005), .B2(G168), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g584(.A(G286), .B(new_n997), .C1(new_n1004), .C2(new_n767), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT51), .B1(new_n1010), .B2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g587(.A(KEYINPUT45), .B(new_n965), .C1(new_n871), .C2(new_n874), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n971), .B1(new_n967), .B2(new_n993), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1971), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND4_X1   g590(.A1(new_n777), .A2(new_n992), .A3(new_n994), .A4(new_n996), .ZN(new_n1016));
  OAI21_X1  g591(.A(G8), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(G8), .B1(new_n571), .B2(new_n572), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT55), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1020), .B(G8), .C1(new_n571), .C2(new_n572), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(KEYINPUT116), .A2(G8), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1023), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1027), .B(G8), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n582), .A2(new_n1030), .A3(new_n586), .ZN(new_n1031));
  INV_X1    g606(.A(G48), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1033));
  OAI22_X1  g608(.A1(new_n531), .A2(new_n1032), .B1(new_n1033), .B2(new_n520), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n538), .A2(new_n579), .ZN(new_n1035));
  OAI21_X1  g610(.A(G1981), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT114), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1007), .B1(new_n1001), .B2(new_n996), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1031), .A2(new_n1036), .A3(new_n1043), .A4(KEYINPUT49), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1038), .A2(new_n1041), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n574), .A2(new_n575), .A3(G1976), .A4(new_n576), .ZN(new_n1046));
  XNOR2_X1  g621(.A(KEYINPUT113), .B(G1976), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(G288), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1042), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(G8), .B(new_n1046), .C1(new_n971), .C2(new_n993), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1050), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT112), .B1(new_n1050), .B2(KEYINPUT52), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1045), .B(new_n1049), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT124), .B1(new_n1029), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT124), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1056), .B(new_n1053), .C1(new_n1025), .C2(new_n1028), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1012), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G2078), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1013), .A2(new_n1014), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(G2078), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n968), .A2(new_n996), .A3(new_n1013), .A4(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n992), .A2(new_n994), .A3(new_n996), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n788), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT125), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1062), .A2(new_n1064), .A3(KEYINPUT125), .A4(new_n1066), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(G171), .A3(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1000), .A2(new_n1003), .A3(new_n1002), .A4(new_n1063), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1062), .A2(new_n1072), .A3(G301), .A4(new_n1066), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1073), .A2(KEYINPUT54), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1062), .A2(new_n1066), .A3(new_n1072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G171), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1062), .A2(new_n1064), .A3(G301), .A4(new_n1066), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT126), .B1(new_n1058), .B2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(G299), .B(KEYINPUT57), .Z(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(G2072), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1013), .A2(new_n1014), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1065), .A2(new_n835), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT119), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1091));
  XNOR2_X1  g666(.A(G299), .B(KEYINPUT57), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT122), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1084), .A2(new_n1087), .A3(new_n1088), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1097), .A3(new_n1092), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1090), .A2(new_n1094), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1348), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n971), .A2(new_n993), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1065), .A2(new_n1102), .B1(new_n983), .B2(new_n1103), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1104), .A2(new_n610), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n610), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n1108));
  AND3_X1   g683(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1013), .A2(new_n1014), .A3(new_n980), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT120), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT58), .B(G1341), .Z(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n971), .B2(new_n993), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1013), .A2(new_n1014), .A3(new_n1116), .A4(new_n980), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n556), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT59), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n1121), .A3(new_n556), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1089), .A2(new_n1093), .A3(KEYINPUT61), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1101), .A2(new_n1111), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1105), .A2(new_n1093), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(new_n1090), .A3(new_n1096), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1029), .A2(new_n1054), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n1056), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1029), .A2(KEYINPUT124), .A3(new_n1054), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1071), .A2(new_n1074), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1012), .A4(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1083), .A2(new_n1128), .A3(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1053), .B(KEYINPUT115), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1005), .A2(new_n1007), .A3(G286), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT63), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1137), .A2(new_n1138), .A3(new_n1141), .A4(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1029), .A2(new_n1141), .A3(new_n1054), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1142), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1045), .A2(new_n715), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1031), .B1(new_n1147), .B2(G288), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1144), .A2(new_n1146), .B1(new_n1042), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1077), .ZN(new_n1150));
  OAI221_X1 g725(.A(new_n1150), .B1(new_n1055), .B2(new_n1057), .C1(KEYINPUT62), .C2(new_n1012), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1140), .B(new_n1149), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n989), .B1(new_n1136), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n973), .B1(new_n878), .B2(new_n984), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT46), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n982), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n979), .A2(KEYINPUT46), .A3(new_n981), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1155), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT47), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n735), .B1(new_n729), .B2(new_n731), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n986), .A2(new_n1161), .B1(new_n983), .B2(new_n759), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n974), .B(KEYINPUT48), .Z(new_n1163));
  OAI22_X1  g738(.A1(new_n1162), .A2(new_n973), .B1(new_n988), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1154), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g741(.A1(G229), .A2(G401), .ZN(new_n1168));
  INV_X1    g742(.A(G319), .ZN(new_n1169));
  NOR2_X1   g743(.A1(G227), .A2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g744(.A(new_n1170), .B(KEYINPUT127), .Z(new_n1171));
  AND4_X1   g745(.A1(new_n900), .A2(new_n961), .A3(new_n1168), .A4(new_n1171), .ZN(G308));
  NAND4_X1  g746(.A1(new_n900), .A2(new_n961), .A3(new_n1168), .A4(new_n1171), .ZN(G225));
endmodule


