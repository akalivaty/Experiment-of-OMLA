//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(KEYINPUT5), .ZN(new_n202));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G155gat), .B(G162gat), .ZN(new_n205));
  XOR2_X1   g004(.A(G141gat), .B(G148gat), .Z(new_n206));
  INV_X1    g005(.A(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT76), .ZN(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n205), .B(new_n206), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215));
  OR2_X1    g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n213), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT75), .ZN(new_n219));
  AND2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n218), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n214), .A2(new_n215), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n215), .B1(new_n214), .B2(new_n224), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G120gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT69), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G120gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n235), .A3(G113gat), .ZN(new_n236));
  INV_X1    g035(.A(G113gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G120gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(KEYINPUT70), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n228), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT70), .B1(new_n236), .B2(new_n238), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n231), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n227), .A2(KEYINPUT77), .A3(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n216), .B(new_n217), .C1(new_n220), .C2(new_n221), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT76), .B(G155gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G162gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n248), .B2(KEYINPUT2), .ZN(new_n249));
  INV_X1    g048(.A(new_n224), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT3), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n214), .A2(new_n215), .A3(new_n224), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n244), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT77), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n204), .B1(new_n245), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n242), .A2(new_n243), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n214), .A2(new_n231), .A3(new_n224), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT79), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n236), .A2(new_n238), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(new_n239), .A3(new_n241), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT2), .ZN(new_n264));
  INV_X1    g063(.A(new_n246), .ZN(new_n265));
  INV_X1    g064(.A(new_n223), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n266), .B1(new_n205), .B2(new_n219), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n264), .A2(new_n265), .B1(new_n267), .B2(new_n218), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT79), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n263), .A2(new_n268), .A3(new_n269), .A4(new_n231), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n259), .A2(new_n270), .A3(KEYINPUT4), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n257), .A2(new_n258), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n271), .A2(KEYINPUT81), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT81), .B1(new_n271), .B2(new_n274), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n202), .B(new_n256), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n214), .A2(new_n224), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n244), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n259), .A2(new_n270), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n202), .B1(new_n280), .B2(new_n204), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT77), .B1(new_n227), .B2(new_n244), .ZN(new_n282));
  AND4_X1   g081(.A1(KEYINPUT77), .A2(new_n251), .A3(new_n244), .A4(new_n252), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n203), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n272), .A2(new_n273), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n259), .A2(new_n270), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n281), .B1(new_n284), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n277), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G1gat), .B(G29gat), .Z(new_n291));
  XNOR2_X1  g090(.A(G57gat), .B(G85gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n290), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n277), .A2(new_n289), .A3(new_n295), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT82), .ZN(new_n301));
  AND4_X1   g100(.A1(new_n301), .A2(new_n290), .A3(KEYINPUT6), .A4(new_n296), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n295), .B1(new_n277), .B2(new_n289), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n301), .B1(new_n303), .B2(KEYINPUT6), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n300), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G8gat), .B(G36gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(G64gat), .B(G92gat), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n306), .B(new_n307), .Z(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT27), .B(G183gat), .ZN(new_n312));
  INV_X1    g111(.A(G190gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT28), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(KEYINPUT28), .A3(new_n313), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT26), .ZN(new_n320));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G169gat), .ZN(new_n323));
  INV_X1    g122(.A(G176gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n318), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT24), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT68), .ZN(new_n331));
  NAND3_X1  g130(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n332));
  INV_X1    g131(.A(G183gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n313), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT68), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n321), .A2(new_n335), .A3(new_n329), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n331), .A2(new_n332), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT25), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n319), .B2(KEYINPUT23), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n341), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n338), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT23), .ZN(new_n344));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT67), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(KEYINPUT67), .A3(new_n345), .ZN(new_n349));
  AND4_X1   g148(.A1(new_n337), .A2(new_n343), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n346), .B1(new_n340), .B2(new_n342), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n313), .A3(KEYINPUT65), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT65), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(G183gat), .B2(G190gat), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n330), .A2(new_n352), .A3(new_n354), .A4(new_n332), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT25), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n328), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n311), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G197gat), .B(G204gat), .ZN(new_n360));
  AND2_X1   g159(.A1(G211gat), .A2(G218gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(KEYINPUT22), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(G211gat), .A2(G218gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n362), .B(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n340), .A2(new_n342), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n344), .A2(new_n345), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(new_n355), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n338), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n337), .A2(new_n343), .A3(new_n348), .A4(new_n349), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n370), .A2(new_n371), .B1(new_n318), .B2(new_n327), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(new_n310), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n359), .A2(new_n366), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n310), .B1(new_n372), .B2(KEYINPUT29), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n311), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n365), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n309), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n366), .B1(new_n359), .B2(new_n373), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(new_n376), .A3(new_n365), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n308), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(KEYINPUT30), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n379), .A2(new_n383), .A3(new_n380), .A4(new_n308), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n305), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387));
  INV_X1    g186(.A(G50gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n365), .A2(new_n358), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT3), .B1(new_n392), .B2(KEYINPUT84), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n365), .A2(new_n394), .A3(new_n358), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n268), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n365), .B1(new_n358), .B2(new_n252), .ZN(new_n397));
  INV_X1    g196(.A(G228gat), .ZN(new_n398));
  INV_X1    g197(.A(G233gat), .ZN(new_n399));
  OAI22_X1  g198(.A1(new_n396), .A2(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n397), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n226), .A2(new_n398), .A3(new_n399), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n401), .B(new_n402), .C1(new_n268), .C2(new_n392), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n391), .B1(new_n404), .B2(G22gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT85), .B(G22gat), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n400), .A2(KEYINPUT86), .A3(new_n406), .A4(new_n403), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n400), .A2(new_n406), .A3(new_n403), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n408), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n406), .B1(new_n400), .B2(new_n403), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n391), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n370), .A2(new_n371), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n416), .A2(new_n244), .A3(new_n328), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n244), .B1(new_n416), .B2(new_n328), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT72), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n244), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n357), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n372), .A2(new_n244), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT72), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n419), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT73), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT73), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n430), .A3(new_n427), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n425), .B(KEYINPUT64), .Z(new_n433));
  NAND3_X1  g232(.A1(new_n421), .A2(new_n422), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT32), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT33), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G15gat), .B(G43gat), .Z(new_n438));
  XNOR2_X1  g237(.A(G71gat), .B(G99gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n440), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n434), .B(KEYINPUT32), .C1(new_n436), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n433), .A2(KEYINPUT34), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n417), .B2(new_n418), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n432), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n431), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n430), .B1(new_n426), .B2(new_n427), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n444), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n415), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n386), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT35), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n452), .A2(KEYINPUT89), .A3(new_n448), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT89), .B1(new_n452), .B2(new_n448), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n305), .A2(new_n455), .A3(new_n385), .A4(new_n415), .ZN(new_n459));
  OAI22_X1  g258(.A1(new_n454), .A2(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n415), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n386), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n245), .A2(new_n255), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n275), .B2(new_n276), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT39), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n204), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n295), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n280), .A2(new_n204), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT39), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n470), .B1(new_n465), .B2(new_n204), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n463), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n465), .A2(new_n204), .ZN(new_n473));
  INV_X1    g272(.A(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(KEYINPUT40), .A3(new_n295), .A4(new_n467), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n385), .A2(new_n303), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT37), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n379), .B2(new_n380), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n481), .B2(new_n308), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT37), .B1(new_n374), .B2(new_n377), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(KEYINPUT88), .A3(new_n309), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n379), .A2(new_n480), .A3(new_n380), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT38), .ZN(new_n487));
  INV_X1    g286(.A(new_n381), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n379), .A2(new_n380), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(KEYINPUT37), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n308), .A2(KEYINPUT38), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n481), .A2(new_n489), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n488), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n415), .B(new_n478), .C1(new_n305), .C2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n451), .A2(new_n444), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n445), .B1(new_n432), .B2(new_n447), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n499), .B1(new_n502), .B2(KEYINPUT74), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT74), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n504), .B(KEYINPUT36), .C1(new_n500), .C2(new_n501), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n462), .A2(new_n498), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n460), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G8gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT16), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(G1gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT94), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n511), .B1(G1gat), .B2(new_n509), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n516));
  AND2_X1   g315(.A1(G43gat), .A2(G50gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(G43gat), .A2(G50gat), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT15), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT92), .B(G43gat), .Z(new_n520));
  AOI211_X1 g319(.A(KEYINPUT15), .B(new_n517), .C1(new_n520), .C2(new_n388), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n523), .A2(KEYINPUT14), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT91), .B(G36gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G29gat), .ZN(new_n526));
  INV_X1    g325(.A(G29gat), .ZN(new_n527));
  INV_X1    g326(.A(G36gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT90), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(new_n523), .A3(KEYINPUT14), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n524), .A2(new_n526), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n519), .B1(new_n521), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(new_n519), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n516), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT93), .A4(KEYINPUT17), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n515), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n515), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(new_n534), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n538), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT18), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n515), .B(new_n534), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n539), .B(KEYINPUT13), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n543), .B2(KEYINPUT18), .ZN(new_n551));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G197gat), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT11), .B(G169gat), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT12), .Z(new_n556));
  NOR3_X1   g355(.A1(new_n546), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n546), .B2(new_n551), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n507), .A2(KEYINPUT95), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT95), .B1(new_n507), .B2(new_n560), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(new_n209), .ZN(new_n565));
  XNOR2_X1  g364(.A(G183gat), .B(G211gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G57gat), .B(G64gat), .Z(new_n569));
  INV_X1    g368(.A(KEYINPUT96), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G71gat), .B(G78gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT9), .ZN(new_n574));
  INV_X1    g373(.A(G71gat), .ZN(new_n575));
  INV_X1    g374(.A(G78gat), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(new_n577), .A3(new_n569), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n569), .A2(new_n577), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(new_n571), .A3(new_n572), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n582));
  AND2_X1   g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G127gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n584), .A2(G127gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n581), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n578), .A2(KEYINPUT97), .A3(new_n580), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n515), .B1(new_n591), .B2(KEYINPUT21), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n586), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n592), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n584), .A2(G127gat), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n594), .B1(new_n595), .B2(new_n585), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n568), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n592), .B1(new_n586), .B2(new_n587), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n594), .A3(new_n585), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n599), .A3(new_n567), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n578), .A2(new_n580), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G99gat), .B(G106gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n603), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n610), .B(new_n611), .Z(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n581), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT10), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(KEYINPUT10), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n589), .B2(new_n590), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n602), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n613), .A2(new_n615), .ZN(new_n620));
  INV_X1    g419(.A(new_n602), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  NAND3_X1  g424(.A1(new_n619), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n619), .A2(new_n622), .ZN(new_n631));
  INV_X1    g430(.A(new_n625), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n612), .B1(new_n536), .B2(new_n537), .ZN(new_n635));
  XOR2_X1   g434(.A(G190gat), .B(G218gat), .Z(new_n636));
  AND2_X1   g435(.A1(G232gat), .A2(G233gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT41), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n534), .B2(new_n614), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n635), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n636), .B1(new_n635), .B2(new_n639), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n637), .A2(KEYINPUT41), .ZN(new_n643));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  XOR2_X1   g444(.A(new_n645), .B(KEYINPUT98), .Z(new_n646));
  NAND3_X1  g445(.A1(new_n641), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n645), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n641), .B2(new_n642), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n601), .A2(new_n634), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n601), .A2(new_n634), .A3(KEYINPUT100), .A4(new_n652), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n563), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n280), .A2(new_n204), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT5), .ZN(new_n660));
  INV_X1    g459(.A(new_n288), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(new_n256), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n202), .B(new_n203), .C1(new_n282), .C2(new_n283), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n271), .A2(new_n274), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT81), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n271), .A2(KEYINPUT81), .A3(new_n274), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n663), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI211_X1 g467(.A(KEYINPUT6), .B(new_n296), .C1(new_n662), .C2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT82), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n303), .A2(new_n301), .A3(KEYINPUT6), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n303), .A2(KEYINPUT6), .ZN(new_n672));
  AOI22_X1  g471(.A1(new_n670), .A2(new_n671), .B1(new_n672), .B2(new_n299), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  INV_X1    g474(.A(new_n385), .ZN(new_n676));
  INV_X1    g475(.A(new_n657), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n676), .B(new_n677), .C1(new_n561), .C2(new_n562), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n678), .A2(G8gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT16), .B(G8gat), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT42), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(KEYINPUT42), .B2(new_n681), .ZN(G1325gat));
  INV_X1    g482(.A(new_n658), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n503), .A2(new_n505), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G15gat), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n458), .A2(G15gat), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n684), .B2(new_n688), .ZN(G1326gat));
  NAND2_X1  g488(.A1(new_n658), .A2(new_n461), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT43), .B(G22gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  INV_X1    g491(.A(new_n601), .ZN(new_n693));
  INV_X1    g492(.A(new_n652), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n634), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT101), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n563), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(new_n527), .A3(new_n673), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  INV_X1    g498(.A(new_n460), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n386), .B2(new_n461), .ZN(new_n702));
  AOI211_X1 g501(.A(KEYINPUT102), .B(new_n415), .C1(new_n305), .C2(new_n385), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n498), .A2(new_n503), .A3(new_n505), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n705), .A3(KEYINPUT103), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n670), .A2(new_n671), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n676), .B1(new_n708), .B2(new_n300), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT102), .B1(new_n709), .B2(new_n415), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n701), .B(new_n461), .C1(new_n673), .C2(new_n676), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n498), .A2(new_n503), .A3(new_n505), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n707), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n700), .B1(new_n706), .B2(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n648), .A2(new_n651), .A3(KEYINPUT104), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT104), .B1(new_n648), .B2(new_n651), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(KEYINPUT44), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n652), .B1(new_n460), .B2(new_n506), .ZN(new_n723));
  OAI22_X1  g522(.A1(new_n715), .A2(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n560), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n630), .A2(new_n633), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n725), .A2(new_n601), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n305), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n699), .A2(new_n729), .ZN(G1328gat));
  INV_X1    g529(.A(new_n525), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n697), .A2(new_n676), .A3(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n525), .B1(new_n728), .B2(new_n385), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(new_n520), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n728), .B2(new_n686), .ZN(new_n738));
  INV_X1    g537(.A(new_n458), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n697), .A2(new_n739), .A3(new_n520), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT106), .B1(new_n728), .B2(new_n686), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n724), .A2(new_n745), .A3(new_n685), .A4(new_n727), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n744), .A2(new_n737), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n740), .A2(KEYINPUT47), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n743), .B1(new_n747), .B2(new_n748), .ZN(G1330gat));
  OAI21_X1  g548(.A(G50gat), .B1(new_n728), .B2(new_n415), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n415), .A2(G50gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT107), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n697), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n750), .A2(new_n753), .A3(KEYINPUT48), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1331gat));
  XNOR2_X1  g557(.A(new_n305), .B(KEYINPUT108), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n725), .A2(new_n601), .A3(new_n652), .A4(new_n726), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n715), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT109), .B(G57gat), .Z(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1332gat));
  OR3_X1    g562(.A1(new_n715), .A2(KEYINPUT110), .A3(new_n760), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT110), .B1(new_n715), .B2(new_n760), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n676), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT49), .B(G64gat), .Z(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(G1333gat));
  NOR2_X1   g569(.A1(new_n715), .A2(new_n760), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n458), .B(KEYINPUT111), .Z(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n575), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n764), .A2(new_n685), .A3(new_n765), .ZN(new_n775));
  AOI211_X1 g574(.A(KEYINPUT50), .B(new_n774), .C1(new_n775), .C2(G71gat), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(G71gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n773), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n776), .A2(new_n779), .ZN(G1334gat));
  NAND2_X1  g579(.A1(new_n766), .A2(new_n461), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g581(.A(new_n722), .B1(new_n507), .B2(new_n694), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT103), .B1(new_n704), .B2(new_n705), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n712), .A2(new_n713), .A3(new_n707), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n460), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n783), .B1(new_n786), .B2(new_n720), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n725), .A2(new_n693), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n634), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT112), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n724), .A2(new_n792), .A3(new_n789), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n791), .A2(new_n673), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n788), .A2(new_n652), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT51), .B1(new_n786), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  INV_X1    g596(.A(new_n795), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n715), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n673), .A2(new_n607), .A3(new_n726), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n794), .A2(new_n607), .B1(new_n800), .B2(new_n801), .ZN(G1336gat));
  NOR3_X1   g601(.A1(new_n634), .A2(G92gat), .A3(new_n385), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT113), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n724), .A2(new_n789), .ZN(new_n806));
  OAI21_X1  g605(.A(G92gat), .B1(new_n806), .B2(new_n385), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n809), .B(new_n803), .C1(new_n796), .C2(new_n799), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n805), .A2(new_n807), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n796), .ZN(new_n812));
  INV_X1    g611(.A(new_n799), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n804), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n791), .A2(new_n676), .A3(new_n793), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(G92gat), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n811), .B1(new_n816), .B2(new_n808), .ZN(G1337gat));
  AND3_X1   g616(.A1(new_n791), .A2(new_n685), .A3(new_n793), .ZN(new_n818));
  INV_X1    g617(.A(G99gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n739), .A2(new_n819), .A3(new_n726), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n818), .A2(new_n819), .B1(new_n800), .B2(new_n820), .ZN(G1338gat));
  XNOR2_X1  g620(.A(KEYINPUT114), .B(G106gat), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n822), .B1(new_n806), .B2(new_n415), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824));
  OR3_X1    g623(.A1(new_n634), .A2(G106gat), .A3(new_n415), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n823), .B(new_n824), .C1(new_n800), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n812), .B2(new_n813), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n791), .A2(new_n461), .A3(new_n793), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n822), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n826), .B1(new_n829), .B2(new_n824), .ZN(G1339gat));
  INV_X1    g629(.A(KEYINPUT104), .ZN(new_n831));
  INV_X1    g630(.A(new_n651), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n647), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n716), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n619), .A2(KEYINPUT54), .ZN(new_n836));
  INV_X1    g635(.A(new_n618), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n837), .B(new_n621), .C1(new_n620), .C2(KEYINPUT10), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT115), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n616), .A2(new_n618), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n841), .A3(new_n621), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n836), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n619), .A2(KEYINPUT54), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n632), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n835), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n843), .A2(new_n845), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n847), .A2(KEYINPUT55), .B1(new_n629), .B2(new_n628), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n560), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n538), .A2(new_n542), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n539), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n548), .A2(new_n549), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n555), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n558), .A2(new_n726), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n834), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n558), .A2(new_n853), .ZN(new_n856));
  INV_X1    g655(.A(new_n843), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n844), .A2(new_n632), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(KEYINPUT55), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n630), .A3(new_n846), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n719), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n693), .B1(new_n855), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n653), .A2(new_n560), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n461), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n673), .A2(new_n385), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n458), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G113gat), .B1(new_n868), .B2(new_n725), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n759), .B1(new_n862), .B2(new_n864), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n453), .A2(new_n676), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n560), .A2(new_n237), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n869), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT117), .ZN(G1340gat));
  OAI21_X1  g676(.A(G120gat), .B1(new_n868), .B2(new_n634), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n726), .A2(new_n233), .A3(new_n235), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n874), .B2(new_n879), .ZN(G1341gat));
  OAI21_X1  g679(.A(G127gat), .B1(new_n868), .B2(new_n693), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n693), .A2(G127gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n872), .B2(new_n882), .ZN(G1342gat));
  NOR3_X1   g682(.A1(new_n872), .A2(G134gat), .A3(new_n652), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT56), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n886), .A2(KEYINPUT118), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(KEYINPUT118), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n865), .A2(new_n694), .A3(new_n867), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT56), .B1(new_n889), .B2(G134gat), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n887), .B(new_n888), .C1(new_n890), .C2(new_n884), .ZN(G1343gat));
  NOR2_X1   g690(.A1(new_n685), .A2(new_n866), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n862), .A2(new_n864), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT57), .B1(new_n893), .B2(new_n461), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n461), .A2(KEYINPUT57), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n847), .A2(KEYINPUT119), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n897), .B1(new_n843), .B2(new_n845), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n896), .A2(new_n835), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n560), .A3(new_n848), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n694), .B1(new_n900), .B2(new_n854), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n693), .B1(new_n901), .B2(new_n861), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n895), .B1(new_n902), .B2(new_n864), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n892), .B1(new_n894), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G141gat), .B1(new_n904), .B2(new_n725), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n870), .A2(new_n385), .A3(new_n461), .A4(new_n686), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n906), .A2(G141gat), .A3(new_n725), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  XOR2_X1   g707(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n909));
  NAND3_X1  g708(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT120), .B(new_n892), .C1(new_n894), .C2(new_n903), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n560), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n907), .B1(new_n914), .B2(G141gat), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(G1344gat));
  OR3_X1    g716(.A1(new_n906), .A2(G148gat), .A3(new_n634), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G148gat), .ZN(new_n920));
  INV_X1    g719(.A(new_n913), .ZN(new_n921));
  OR3_X1    g720(.A1(new_n719), .A2(new_n856), .A3(new_n860), .ZN(new_n922));
  INV_X1    g721(.A(new_n854), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n859), .A2(new_n630), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n924), .B1(new_n559), .B2(new_n558), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n923), .B1(new_n925), .B2(new_n899), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n922), .B1(new_n926), .B2(new_n694), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n863), .B1(new_n927), .B2(new_n693), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n415), .B1(new_n862), .B2(new_n864), .ZN(new_n929));
  OAI22_X1  g728(.A1(new_n928), .A2(new_n895), .B1(new_n929), .B2(KEYINPUT57), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT120), .B1(new_n930), .B2(new_n892), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n921), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n920), .B1(new_n932), .B2(new_n726), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n856), .A2(new_n860), .A3(new_n652), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n693), .B1(new_n901), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT122), .B1(new_n657), .B2(new_n560), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT122), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n655), .A2(new_n937), .A3(new_n725), .A4(new_n656), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT57), .B1(new_n939), .B2(new_n461), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n895), .B1(new_n862), .B2(new_n864), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n726), .A3(new_n892), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n919), .B1(new_n943), .B2(G148gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n918), .B1(new_n933), .B2(new_n944), .ZN(G1345gat));
  NAND2_X1  g744(.A1(new_n912), .A2(new_n913), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n247), .B1(new_n946), .B2(new_n693), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n601), .A2(new_n210), .A3(new_n211), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n906), .B2(new_n948), .ZN(G1346gat));
  NOR3_X1   g748(.A1(new_n906), .A2(G162gat), .A3(new_n652), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT123), .Z(new_n951));
  OAI21_X1  g750(.A(G162gat), .B1(new_n946), .B2(new_n719), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1347gat));
  NAND4_X1  g752(.A1(new_n865), .A2(new_n676), .A3(new_n759), .A4(new_n772), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n954), .A2(new_n323), .A3(new_n725), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n673), .B1(new_n862), .B2(new_n864), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n956), .A2(new_n676), .A3(new_n415), .A4(new_n502), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n560), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n955), .B1(new_n323), .B2(new_n959), .ZN(G1348gat));
  OAI21_X1  g759(.A(G176gat), .B1(new_n954), .B2(new_n634), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n726), .A2(new_n324), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n957), .B2(new_n962), .ZN(G1349gat));
  OAI21_X1  g762(.A(G183gat), .B1(new_n954), .B2(new_n693), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n601), .A2(new_n312), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n957), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g766(.A1(new_n958), .A2(new_n313), .A3(new_n834), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n954), .A2(new_n652), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n970));
  AND4_X1   g769(.A1(KEYINPUT124), .A2(new_n969), .A3(new_n970), .A4(G190gat), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT124), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n313), .B1(new_n972), .B2(KEYINPUT61), .ZN(new_n973));
  AOI22_X1  g772(.A1(new_n969), .A2(new_n973), .B1(KEYINPUT124), .B2(new_n970), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n968), .B1(new_n971), .B2(new_n974), .ZN(G1351gat));
  INV_X1    g774(.A(new_n759), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n976), .A2(new_n385), .A3(new_n685), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n942), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(G197gat), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n978), .A2(new_n979), .A3(new_n725), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n686), .A2(new_n676), .A3(new_n461), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n981), .A2(KEYINPUT125), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(KEYINPUT125), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n982), .A2(new_n956), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(G197gat), .B1(new_n984), .B2(new_n560), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n980), .A2(new_n985), .ZN(G1352gat));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n987));
  INV_X1    g786(.A(G204gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n984), .A2(new_n988), .A3(new_n726), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n987), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n994), .A2(KEYINPUT62), .A3(new_n990), .ZN(new_n995));
  OAI21_X1  g794(.A(G204gat), .B1(new_n978), .B2(new_n634), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(G1353gat));
  OAI211_X1 g796(.A(new_n601), .B(new_n977), .C1(new_n940), .C2(new_n941), .ZN(new_n998));
  AOI21_X1  g797(.A(KEYINPUT63), .B1(new_n998), .B2(G211gat), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n693), .A2(G211gat), .ZN(new_n1001));
  AOI22_X1  g800(.A1(new_n999), .A2(new_n1000), .B1(new_n984), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n998), .A2(G211gat), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT63), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(KEYINPUT127), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1002), .B1(new_n1006), .B2(new_n1007), .ZN(G1354gat));
  OAI21_X1  g807(.A(G218gat), .B1(new_n978), .B2(new_n652), .ZN(new_n1009));
  INV_X1    g808(.A(G218gat), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n984), .A2(new_n1010), .A3(new_n834), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1009), .A2(new_n1011), .ZN(G1355gat));
endmodule


