//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  XNOR2_X1  g000(.A(KEYINPUT26), .B(G101), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G146), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(new_n193), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n203), .A3(new_n193), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(G143), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n199), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OR2_X1    g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n197), .A2(new_n199), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G137), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n209), .B1(new_n211), .B2(KEYINPUT11), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(G137), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  OAI211_X1 g028(.A(KEYINPUT65), .B(new_n214), .C1(new_n210), .C2(G137), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(KEYINPUT11), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n213), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n217), .A2(G131), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(G131), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n208), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n196), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n202), .A2(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n226));
  OAI21_X1  g040(.A(G143), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n224), .B1(new_n227), .B2(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n204), .A2(new_n205), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT66), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n193), .B1(new_n201), .B2(new_n203), .ZN(new_n232));
  OAI21_X1  g046(.A(G128), .B1(new_n232), .B2(new_n221), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n229), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n223), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G131), .ZN(new_n237));
  INV_X1    g051(.A(new_n211), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(new_n213), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n219), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n220), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT70), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT2), .A2(G113), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT2), .ZN(new_n244));
  INV_X1    g058(.A(G113), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT67), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT67), .B1(new_n244), .B2(new_n245), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n243), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(G116), .B(G119), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n249), .B(new_n243), .C1(new_n246), .C2(new_n247), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n223), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n233), .A2(new_n229), .A3(new_n234), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n234), .B1(new_n233), .B2(new_n229), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n219), .A2(new_n239), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(new_n220), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n242), .A2(new_n254), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n241), .A2(new_n253), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n254), .B(new_n220), .C1(new_n236), .C2(new_n240), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT69), .B1(new_n268), .B2(KEYINPUT28), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n270));
  AOI211_X1 g084(.A(new_n270), .B(new_n264), .C1(new_n266), .C2(new_n267), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n265), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n260), .B2(new_n220), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n273), .B(new_n220), .C1(new_n236), .C2(new_n240), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n253), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n192), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(new_n267), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT31), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n267), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n241), .A2(KEYINPUT30), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n275), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n284), .B2(new_n253), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT31), .A3(new_n278), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n192), .A2(new_n272), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(G472), .A2(G902), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n288), .B(KEYINPUT71), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT32), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n254), .B1(new_n260), .B2(new_n220), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT28), .B1(new_n291), .B2(new_n282), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n270), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT69), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n293), .A2(new_n295), .B1(new_n264), .B2(new_n263), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT31), .B1(new_n285), .B2(new_n278), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n254), .B1(new_n283), .B2(new_n275), .ZN(new_n298));
  NOR4_X1   g112(.A1(new_n298), .A2(new_n280), .A3(new_n192), .A4(new_n282), .ZN(new_n299));
  OAI22_X1  g113(.A1(new_n296), .A2(new_n278), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  INV_X1    g115(.A(new_n289), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n192), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n265), .A2(new_n292), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n294), .B1(new_n264), .B2(new_n263), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n305), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n278), .B(new_n265), .C1(new_n269), .C2(new_n271), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n192), .B1(new_n298), .B2(new_n282), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n304), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n290), .A2(new_n303), .B1(new_n316), .B2(G472), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n318), .A2(KEYINPUT16), .A3(G140), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT73), .B1(new_n321), .B2(G146), .ZN(new_n322));
  NAND2_X1  g136(.A1(G125), .A2(G140), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(G125), .A2(G140), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT16), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n319), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(new_n200), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n326), .A2(new_n327), .A3(G146), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n322), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G128), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n224), .A2(G119), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT24), .B(G110), .Z(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n334), .A2(KEYINPUT23), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(KEYINPUT23), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n339), .B(new_n340), .C1(G119), .C2(new_n224), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G110), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n332), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  OAI22_X1  g157(.A1(new_n341), .A2(G110), .B1(new_n336), .B2(new_n337), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n201), .A2(new_n203), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n320), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n331), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G953), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(G221), .A3(G234), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(G137), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT74), .B(KEYINPUT22), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n343), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n352), .B1(new_n343), .B2(new_n347), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OR3_X1    g169(.A1(new_n355), .A2(KEYINPUT25), .A3(G902), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(G234), .B2(new_n315), .ZN(new_n358));
  OAI21_X1  g172(.A(KEYINPUT25), .B1(new_n355), .B2(G902), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  OR3_X1    g174(.A1(new_n355), .A2(G902), .A3(new_n358), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n317), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G214), .B1(G237), .B2(G902), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n364), .B(KEYINPUT78), .Z(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n348), .A2(G952), .ZN(new_n367));
  NAND2_X1  g181(.A1(G234), .A2(G237), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  XOR2_X1   g184(.A(KEYINPUT21), .B(G898), .Z(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(G902), .A3(G953), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n208), .A2(G125), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(new_n318), .B2(new_n258), .ZN(new_n378));
  INV_X1    g192(.A(G224), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G953), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n378), .B(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(new_n385), .B2(G107), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  INV_X1    g201(.A(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G104), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n385), .A2(G107), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n386), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G101), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT75), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT75), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n391), .A2(new_n395), .A3(new_n392), .A4(G101), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n392), .B1(new_n391), .B2(G101), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n386), .A2(new_n389), .A3(new_n399), .A4(new_n390), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n253), .A3(new_n401), .ZN(new_n402));
  XOR2_X1   g216(.A(G110), .B(G122), .Z(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n333), .A2(G116), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT80), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n249), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n405), .A2(new_n410), .A3(G116), .A4(new_n333), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n408), .A2(G113), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n390), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n385), .A2(G107), .ZN(new_n414));
  OAI21_X1  g228(.A(G101), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n400), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n412), .A2(new_n252), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n402), .A2(new_n404), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n402), .A2(KEYINPUT82), .A3(new_n418), .A4(new_n404), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n402), .A2(new_n418), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT81), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n402), .A2(new_n426), .A3(new_n418), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(new_n403), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n384), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n402), .A2(new_n426), .A3(new_n418), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n426), .B1(new_n402), .B2(new_n418), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n430), .A2(new_n431), .A3(new_n404), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(KEYINPUT6), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n383), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n378), .A2(new_n380), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n412), .A2(new_n252), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n416), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT83), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n408), .A2(G113), .A3(new_n411), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n252), .B(new_n417), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n442), .A3(new_n416), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n403), .B(KEYINPUT8), .Z(new_n445));
  AOI22_X1  g259(.A1(new_n435), .A2(KEYINPUT7), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n381), .A2(KEYINPUT7), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n421), .A2(new_n422), .B1(new_n378), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(G902), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G210), .B1(G237), .B2(G902), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n434), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n434), .B2(new_n449), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n366), .B(new_n376), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n258), .A2(KEYINPUT10), .A3(new_n417), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n394), .A2(new_n396), .B1(new_n400), .B2(new_n398), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n205), .A2(KEYINPUT76), .A3(KEYINPUT1), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT76), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n224), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n456), .A2(new_n459), .B1(new_n227), .B2(new_n194), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n417), .B1(new_n460), .B2(new_n223), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT10), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n208), .A2(new_n455), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n218), .A2(new_n219), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n454), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G140), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n348), .A2(G227), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n466), .B(new_n467), .Z(new_n468));
  OAI211_X1 g282(.A(new_n255), .B(new_n416), .C1(new_n256), .C2(new_n257), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n461), .ZN(new_n470));
  INV_X1    g284(.A(new_n464), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT12), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT12), .ZN(new_n473));
  AOI211_X1 g287(.A(new_n473), .B(new_n464), .C1(new_n469), .C2(new_n461), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n465), .B(new_n468), .C1(new_n472), .C2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n468), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n454), .A2(new_n464), .A3(new_n463), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n464), .B1(new_n454), .B2(new_n463), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(KEYINPUT77), .A2(G469), .ZN(new_n481));
  OR2_X1    g295(.A1(KEYINPUT77), .A2(G469), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n480), .A2(new_n315), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n465), .B1(new_n472), .B2(new_n474), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n476), .ZN(new_n485));
  INV_X1    g299(.A(new_n478), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n465), .A3(new_n468), .ZN(new_n487));
  AOI21_X1  g301(.A(G902), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G469), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n483), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT9), .B(G234), .ZN(new_n491));
  OAI21_X1  g305(.A(G221), .B1(new_n491), .B2(G902), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OR2_X1    g307(.A1(G475), .A2(G902), .ZN(new_n494));
  XNOR2_X1  g308(.A(G113), .B(G122), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n385), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(KEYINPUT18), .A2(G131), .ZN(new_n498));
  INV_X1    g312(.A(G237), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n348), .A3(G214), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n193), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n325), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(G146), .A3(new_n323), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n502), .A3(new_n498), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT84), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT84), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n501), .A2(new_n508), .A3(new_n502), .A4(new_n498), .ZN(new_n509));
  AOI221_X4 g323(.A(new_n503), .B1(new_n346), .B2(new_n505), .C1(new_n507), .C2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(KEYINPUT19), .A3(new_n323), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT19), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n324), .B2(new_n325), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n331), .B1(new_n514), .B2(new_n195), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n500), .A2(new_n193), .ZN(new_n516));
  AOI21_X1  g330(.A(G143), .B1(new_n190), .B2(G214), .ZN(new_n517));
  OAI21_X1  g331(.A(G131), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n501), .A2(new_n237), .A3(new_n502), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n497), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n507), .A2(new_n509), .ZN(new_n522));
  INV_X1    g336(.A(new_n503), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n346), .A2(new_n505), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n501), .A2(new_n502), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n527), .B2(G131), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n518), .A2(new_n519), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n525), .B(new_n496), .C1(new_n530), .C2(new_n332), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT85), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT85), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n521), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n494), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT20), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT86), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT86), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n521), .A2(new_n531), .A3(new_n534), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n534), .B1(new_n521), .B2(new_n531), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n539), .B(KEYINPUT20), .C1(new_n542), .C2(new_n494), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT20), .B1(new_n494), .B2(KEYINPUT87), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n532), .B(new_n544), .C1(KEYINPUT87), .C2(new_n494), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n530), .A2(new_n332), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n496), .B1(new_n547), .B2(new_n525), .ZN(new_n548));
  INV_X1    g362(.A(new_n531), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n315), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G475), .ZN(new_n551));
  INV_X1    g365(.A(G478), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G128), .B(G143), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n210), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT89), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n210), .B1(new_n555), .B2(KEYINPUT13), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n193), .A2(G128), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n558), .B1(KEYINPUT13), .B2(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(G116), .B(G122), .Z(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT88), .ZN(new_n562));
  XNOR2_X1  g376(.A(G116), .B(G122), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT88), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(new_n388), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n388), .B1(new_n562), .B2(new_n565), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n557), .B(new_n560), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n555), .B(new_n210), .ZN(new_n570));
  INV_X1    g384(.A(G116), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(KEYINPUT14), .A3(G122), .ZN(new_n572));
  OAI211_X1 g386(.A(G107), .B(new_n572), .C1(new_n561), .C2(KEYINPUT14), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n491), .A2(new_n357), .A3(G953), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n569), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n575), .B1(new_n569), .B2(new_n574), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n315), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT90), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(KEYINPUT90), .B(new_n315), .C1(new_n576), .C2(new_n577), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n554), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n553), .B1(new_n578), .B2(new_n579), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n546), .A2(new_n551), .A3(new_n584), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n453), .A2(new_n493), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n363), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  INV_X1    g402(.A(new_n450), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n421), .A2(new_n422), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT6), .B1(new_n590), .B2(new_n432), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n428), .A2(new_n384), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n382), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n435), .A2(KEYINPUT7), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n444), .A2(new_n445), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n448), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n315), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n589), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT92), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n434), .A2(new_n449), .A3(new_n450), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n452), .A2(KEYINPUT92), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n601), .A2(new_n366), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n546), .A2(new_n551), .ZN(new_n604));
  INV_X1    g418(.A(new_n577), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n569), .A2(new_n574), .A3(new_n575), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT33), .ZN(new_n608));
  OR3_X1    g422(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT33), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n609), .A3(G478), .ZN(new_n610));
  NAND2_X1  g424(.A1(G478), .A2(G902), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(new_n552), .A3(new_n315), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n604), .A2(new_n376), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n603), .A2(KEYINPUT93), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n601), .A2(new_n366), .A3(new_n602), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(new_n615), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n287), .A2(new_n289), .ZN(new_n622));
  INV_X1    g436(.A(new_n362), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n490), .A2(new_n623), .A3(new_n492), .ZN(new_n624));
  INV_X1    g438(.A(G472), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n272), .A2(new_n192), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n281), .A2(new_n286), .ZN(new_n627));
  AOI21_X1  g441(.A(G902), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n625), .B1(new_n628), .B2(KEYINPUT91), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT91), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n287), .B2(G902), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n622), .B(new_n624), .C1(new_n629), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n621), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n385), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(new_n584), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n536), .A2(new_n537), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n538), .A2(new_n543), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n637), .A2(new_n639), .A3(new_n551), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n619), .A2(new_n375), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  INV_X1    g458(.A(new_n622), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n300), .A2(KEYINPUT91), .A3(new_n315), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n631), .A2(G472), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n343), .A2(new_n347), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n352), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n650), .B(new_n315), .C1(new_n357), .C2(G234), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n360), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n586), .A2(new_n645), .A3(new_n647), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  NAND2_X1  g469(.A1(new_n290), .A2(new_n303), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n309), .B1(new_n308), .B2(new_n305), .ZN(new_n657));
  AND4_X1   g471(.A1(new_n309), .A2(new_n265), .A3(new_n292), .A4(new_n305), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n315), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n312), .A2(new_n304), .A3(new_n313), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n493), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n369), .B(KEYINPUT95), .Z(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(new_n374), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n493), .A2(new_n640), .A3(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n662), .A2(new_n603), .A3(new_n652), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  NOR2_X1   g482(.A1(new_n285), .A2(new_n192), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n315), .B1(new_n268), .B2(new_n278), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n656), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n604), .A2(new_n637), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n673), .A2(new_n365), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n493), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n665), .B(KEYINPUT39), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT40), .Z(new_n679));
  INV_X1    g493(.A(new_n652), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n598), .A2(new_n600), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT38), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n675), .A2(new_n679), .A3(new_n680), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G143), .ZN(G45));
  INV_X1    g498(.A(new_n665), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n604), .A2(new_n614), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n662), .A2(new_n603), .A3(new_n652), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G146), .ZN(G48));
  NAND2_X1  g503(.A1(new_n480), .A2(new_n315), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n691), .A2(new_n483), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n492), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n317), .A2(new_n362), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n621), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT96), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n695), .B(new_n697), .ZN(G15));
  NAND2_X1  g512(.A1(new_n694), .A2(new_n641), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  NOR2_X1   g514(.A1(new_n317), .A2(new_n375), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n585), .A2(new_n680), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT97), .ZN(new_n703));
  INV_X1    g517(.A(new_n693), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n703), .B1(new_n603), .B2(new_n704), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n619), .A2(new_n693), .A3(KEYINPUT97), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n701), .B(new_n702), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT98), .B(G119), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G21));
  OAI21_X1  g523(.A(G472), .B1(new_n287), .B2(G902), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n297), .A2(new_n299), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n308), .A2(new_n278), .ZN(new_n712));
  OAI211_X1 g526(.A(KEYINPUT99), .B(new_n302), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT99), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n265), .A2(new_n292), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n281), .A2(new_n286), .B1(new_n715), .B2(new_n192), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n714), .B1(new_n716), .B2(new_n289), .ZN(new_n717));
  AND4_X1   g531(.A1(new_n623), .A2(new_n710), .A3(new_n713), .A4(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n619), .A2(new_n674), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n718), .A2(new_n376), .A3(new_n719), .A4(new_n704), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NAND4_X1  g535(.A1(new_n710), .A2(new_n652), .A3(new_n713), .A4(new_n717), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n686), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n705), .B2(new_n706), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT100), .B(G125), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G27));
  NOR3_X1   g540(.A1(new_n287), .A2(KEYINPUT32), .A3(new_n289), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n301), .B1(new_n300), .B2(new_n302), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n661), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n598), .A2(new_n366), .A3(new_n600), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n686), .A2(new_n493), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n731), .A3(new_n623), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(KEYINPUT101), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(KEYINPUT101), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n363), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT102), .B(G131), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G33));
  NOR3_X1   g553(.A1(new_n451), .A2(new_n452), .A3(new_n365), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n729), .A2(new_n623), .A3(new_n666), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  AND2_X1   g556(.A1(new_n485), .A2(new_n487), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n743), .A2(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(KEYINPUT45), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(G469), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(G469), .A2(G902), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n483), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n748), .A2(new_n753), .A3(new_n749), .ZN(new_n754));
  OAI211_X1 g568(.A(KEYINPUT103), .B(new_n483), .C1(new_n748), .C2(new_n749), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n748), .A2(new_n749), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT104), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n752), .A2(new_n754), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n492), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n604), .B2(KEYINPUT105), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n604), .A2(new_n613), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n647), .A2(new_n645), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n764), .A2(new_n765), .A3(new_n652), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n730), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n767), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n760), .A2(new_n677), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  NAND4_X1  g586(.A1(new_n317), .A2(new_n362), .A3(new_n687), .A4(new_n740), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT106), .Z(new_n774));
  AND3_X1   g588(.A1(new_n758), .A2(KEYINPUT47), .A3(new_n492), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT47), .B1(new_n758), .B2(new_n492), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  INV_X1    g592(.A(new_n692), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(KEYINPUT49), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(KEYINPUT49), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n623), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n763), .A2(new_n492), .A3(new_n366), .ZN(new_n783));
  OR4_X1    g597(.A1(new_n682), .A2(new_n782), .A3(new_n672), .A4(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n764), .A2(new_n663), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(new_n718), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n740), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT114), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n775), .A2(new_n776), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n779), .A2(new_n492), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n722), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n693), .A2(new_n730), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n785), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n673), .A2(new_n623), .A3(new_n370), .A4(new_n793), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n604), .A3(new_n614), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n682), .A2(new_n366), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n786), .A2(new_n704), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n791), .A2(new_n794), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n791), .A2(KEYINPUT51), .A3(new_n794), .A4(new_n802), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n786), .B1(new_n706), .B2(new_n705), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n785), .A2(new_n363), .A3(new_n793), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n807), .B(new_n367), .C1(new_n808), .C2(KEYINPUT48), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(KEYINPUT48), .B2(new_n808), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n805), .A2(new_n806), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT108), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT107), .B1(new_n604), .B2(new_n614), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n815), .B(new_n613), .C1(new_n546), .C2(new_n551), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n813), .B1(new_n817), .B2(new_n453), .ZN(new_n818));
  INV_X1    g632(.A(new_n453), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n819), .B(KEYINPUT108), .C1(new_n814), .C2(new_n816), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n632), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n587), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT109), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n637), .A2(new_n546), .A3(new_n551), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n453), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n624), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n647), .A2(new_n825), .A3(new_n645), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n823), .B1(new_n653), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n653), .A2(new_n823), .A3(new_n827), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n822), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n695), .A2(new_n707), .A3(new_n699), .A4(new_n720), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n582), .A2(new_n583), .A3(new_n665), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n639), .A2(new_n833), .A3(new_n551), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT110), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT110), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n639), .A2(new_n833), .A3(new_n836), .A4(new_n551), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n740), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n740), .A2(new_n835), .A3(KEYINPUT111), .A4(new_n837), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n662), .A2(new_n840), .A3(new_n652), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n792), .A2(new_n731), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(KEYINPUT112), .A3(new_n741), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n841), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n729), .A2(new_n676), .A3(new_n652), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n741), .B(new_n843), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n847), .A2(new_n848), .B1(new_n736), .B2(new_n734), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n831), .A2(new_n832), .A3(new_n844), .A4(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n493), .A2(new_n665), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n672), .A2(new_n719), .A3(new_n680), .A4(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n724), .A2(new_n667), .A3(new_n688), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT52), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n317), .A2(new_n493), .A3(new_n680), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n855), .B(new_n603), .C1(new_n666), .C2(new_n687), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n724), .A4(new_n852), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n812), .B1(new_n850), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n854), .A2(new_n858), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n653), .A2(new_n823), .A3(new_n827), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n587), .B(new_n821), .C1(new_n862), .C2(new_n828), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n707), .A2(new_n695), .A3(new_n699), .A4(new_n720), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n847), .A2(new_n848), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n866), .A2(new_n737), .A3(new_n844), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n861), .A2(KEYINPUT53), .A3(new_n865), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n860), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(KEYINPUT113), .B(new_n812), .C1(new_n850), .C2(new_n859), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n873));
  AOI211_X1 g687(.A(new_n613), .B(new_n795), .C1(new_n551), .C2(new_n546), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n860), .B2(new_n868), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n811), .A2(new_n873), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(G952), .A2(G953), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n784), .B1(new_n877), .B2(new_n878), .ZN(G75));
  NAND4_X1  g693(.A1(new_n870), .A2(G210), .A3(G902), .A4(new_n871), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n382), .B(KEYINPUT55), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n429), .A2(new_n433), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT115), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n348), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n889), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n885), .A2(new_n886), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n890), .A2(new_n892), .A3(new_n894), .ZN(G51));
  NAND2_X1  g709(.A1(new_n870), .A2(new_n871), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n875), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n747), .B(KEYINPUT57), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n480), .ZN(new_n900));
  OR3_X1    g714(.A1(new_n896), .A2(new_n315), .A3(new_n746), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n891), .B1(new_n900), .B2(new_n901), .ZN(G54));
  NAND4_X1  g716(.A1(new_n872), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n542), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n891), .ZN(G60));
  AND2_X1   g719(.A1(new_n608), .A2(new_n609), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n873), .A2(new_n876), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n611), .B(KEYINPUT59), .Z(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n906), .A2(new_n908), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n897), .A2(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n909), .A2(new_n892), .A3(new_n911), .ZN(G63));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT117), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT60), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n872), .A2(KEYINPUT118), .A3(new_n650), .A4(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n870), .A2(new_n871), .A3(new_n915), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n891), .B1(new_n917), .B2(new_n355), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n870), .A2(new_n650), .A3(new_n871), .A4(new_n915), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT118), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n916), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT116), .ZN(new_n923));
  XNOR2_X1  g737(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(G66));
  OAI21_X1  g741(.A(G953), .B1(new_n372), .B2(new_n379), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n865), .B2(G953), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n893), .B1(G898), .B2(new_n348), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  NAND4_X1  g745(.A1(new_n760), .A2(new_n363), .A3(new_n677), .A4(new_n719), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n777), .A2(new_n771), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n856), .A2(new_n724), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n856), .A2(KEYINPUT121), .A3(new_n724), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n936), .A2(new_n737), .A3(new_n741), .A4(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n348), .B1(new_n933), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n348), .A2(G900), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT123), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n514), .B(KEYINPUT120), .Z(new_n944));
  XNOR2_X1  g758(.A(new_n284), .B(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n939), .A2(new_n947), .A3(new_n941), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n943), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n348), .B1(G227), .B2(G900), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT124), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n936), .A2(new_n683), .A3(new_n937), .ZN(new_n953));
  AND2_X1   g767(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n777), .A2(new_n771), .ZN(new_n956));
  NOR2_X1   g770(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n953), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n678), .B1(new_n817), .B2(new_n824), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n363), .A3(new_n740), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n955), .A2(new_n956), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n348), .A3(new_n945), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n949), .A2(new_n952), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n950), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n963), .B(new_n965), .ZN(G72));
  XNOR2_X1  g780(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n625), .A2(new_n315), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n967), .B(new_n968), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n279), .A2(new_n313), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n970), .B(new_n971), .C1(new_n860), .C2(new_n868), .ZN(new_n972));
  INV_X1    g786(.A(new_n865), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n961), .A2(new_n973), .ZN(new_n974));
  AOI211_X1 g788(.A(new_n192), .B(new_n285), .C1(new_n974), .C2(new_n969), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n933), .A2(new_n938), .A3(new_n973), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n192), .B(new_n285), .C1(new_n976), .C2(new_n970), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n892), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n978), .A2(KEYINPUT126), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(KEYINPUT126), .ZN(new_n980));
  AOI211_X1 g794(.A(new_n972), .B(new_n975), .C1(new_n979), .C2(new_n980), .ZN(G57));
endmodule


