

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U553 ( .A(n597), .B(n596), .ZN(n646) );
  AND2_X1 U554 ( .A1(n595), .A2(G40), .ZN(n721) );
  AND2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n875) );
  INV_X2 U556 ( .A(G2105), .ZN(n523) );
  BUF_X2 U557 ( .A(n638), .Z(n640) );
  AND2_X2 U558 ( .A1(n721), .A2(n722), .ZN(n597) );
  AND2_X1 U559 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U560 ( .A(n648), .B(n647), .ZN(n701) );
  INV_X1 U561 ( .A(n646), .ZN(n638) );
  AND2_X1 U562 ( .A1(n527), .A2(n526), .ZN(G164) );
  NOR2_X1 U563 ( .A1(n656), .A2(n655), .ZN(n658) );
  XNOR2_X1 U564 ( .A(n658), .B(n657), .ZN(n659) );
  INV_X1 U565 ( .A(KEYINPUT5), .ZN(n536) );
  OR2_X1 U566 ( .A1(n518), .A2(n628), .ZN(n631) );
  XNOR2_X1 U567 ( .A(n637), .B(n636), .ZN(n645) );
  INV_X1 U568 ( .A(KEYINPUT29), .ZN(n636) );
  XNOR2_X1 U569 ( .A(n579), .B(n578), .ZN(n583) );
  INV_X1 U570 ( .A(KEYINPUT23), .ZN(n578) );
  XNOR2_X1 U571 ( .A(n581), .B(n580), .ZN(n582) );
  INV_X1 U572 ( .A(KEYINPUT65), .ZN(n580) );
  NAND2_X1 U573 ( .A1(n880), .A2(G137), .ZN(n585) );
  XOR2_X1 U574 ( .A(KEYINPUT71), .B(n541), .Z(G168) );
  AND2_X1 U575 ( .A1(n649), .A2(G1341), .ZN(n517) );
  AND2_X1 U576 ( .A1(n617), .A2(n616), .ZN(n518) );
  NAND2_X1 U577 ( .A1(n650), .A2(G8), .ZN(n651) );
  XNOR2_X1 U578 ( .A(n651), .B(KEYINPUT30), .ZN(n652) );
  NOR2_X1 U579 ( .A1(G1966), .A2(n701), .ZN(n675) );
  INV_X1 U580 ( .A(KEYINPUT87), .ZN(n647) );
  NOR2_X1 U581 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U582 ( .A1(G651), .A2(G543), .ZN(n785) );
  INV_X1 U583 ( .A(KEYINPUT17), .ZN(n519) );
  NOR2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XNOR2_X2 U585 ( .A(n520), .B(n519), .ZN(n880) );
  NAND2_X1 U586 ( .A1(n880), .A2(G138), .ZN(n527) );
  NAND2_X1 U587 ( .A1(G114), .A2(n875), .ZN(n522) );
  NOR2_X4 U588 ( .A1(n523), .A2(G2104), .ZN(n876) );
  NAND2_X1 U589 ( .A1(n876), .A2(G126), .ZN(n521) );
  AND2_X1 U590 ( .A1(n522), .A2(n521), .ZN(n525) );
  AND2_X2 U591 ( .A1(n523), .A2(G2104), .ZN(n879) );
  NAND2_X1 U592 ( .A1(G102), .A2(n879), .ZN(n524) );
  AND2_X1 U593 ( .A1(n525), .A2(n524), .ZN(n526) );
  INV_X1 U594 ( .A(G651), .ZN(n532) );
  NOR2_X1 U595 ( .A1(G543), .A2(n532), .ZN(n528) );
  XOR2_X2 U596 ( .A(KEYINPUT1), .B(n528), .Z(n789) );
  NAND2_X1 U597 ( .A1(G63), .A2(n789), .ZN(n530) );
  XOR2_X1 U598 ( .A(G543), .B(KEYINPUT0), .Z(n567) );
  NOR2_X2 U599 ( .A1(G651), .A2(n567), .ZN(n791) );
  NAND2_X1 U600 ( .A1(G51), .A2(n791), .ZN(n529) );
  NAND2_X1 U601 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U602 ( .A(KEYINPUT6), .B(n531), .ZN(n539) );
  NOR2_X1 U603 ( .A1(n567), .A2(n532), .ZN(n786) );
  NAND2_X1 U604 ( .A1(G76), .A2(n786), .ZN(n535) );
  NAND2_X1 U605 ( .A1(n785), .A2(G89), .ZN(n533) );
  XNOR2_X1 U606 ( .A(n533), .B(KEYINPUT4), .ZN(n534) );
  NAND2_X1 U607 ( .A1(n535), .A2(n534), .ZN(n537) );
  XNOR2_X1 U608 ( .A(n537), .B(n536), .ZN(n538) );
  NOR2_X1 U609 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U610 ( .A(KEYINPUT7), .B(n540), .Z(n541) );
  NAND2_X1 U611 ( .A1(G91), .A2(n785), .ZN(n543) );
  NAND2_X1 U612 ( .A1(G78), .A2(n786), .ZN(n542) );
  NAND2_X1 U613 ( .A1(n543), .A2(n542), .ZN(n546) );
  NAND2_X1 U614 ( .A1(G53), .A2(n791), .ZN(n544) );
  XNOR2_X1 U615 ( .A(KEYINPUT67), .B(n544), .ZN(n545) );
  NOR2_X1 U616 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X1 U617 ( .A1(n789), .A2(G65), .ZN(n547) );
  NAND2_X1 U618 ( .A1(n548), .A2(n547), .ZN(G299) );
  NAND2_X1 U619 ( .A1(G64), .A2(n789), .ZN(n550) );
  NAND2_X1 U620 ( .A1(G52), .A2(n791), .ZN(n549) );
  NAND2_X1 U621 ( .A1(n550), .A2(n549), .ZN(n555) );
  NAND2_X1 U622 ( .A1(G90), .A2(n785), .ZN(n552) );
  NAND2_X1 U623 ( .A1(G77), .A2(n786), .ZN(n551) );
  NAND2_X1 U624 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U625 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U626 ( .A1(n555), .A2(n554), .ZN(G171) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(n556) );
  XNOR2_X1 U628 ( .A(KEYINPUT72), .B(n556), .ZN(G286) );
  NAND2_X1 U629 ( .A1(G88), .A2(n785), .ZN(n558) );
  NAND2_X1 U630 ( .A1(G75), .A2(n786), .ZN(n557) );
  NAND2_X1 U631 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U632 ( .A1(G50), .A2(n791), .ZN(n559) );
  XNOR2_X1 U633 ( .A(KEYINPUT77), .B(n559), .ZN(n560) );
  NOR2_X1 U634 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U635 ( .A1(n789), .A2(G62), .ZN(n562) );
  NAND2_X1 U636 ( .A1(n563), .A2(n562), .ZN(G303) );
  NAND2_X1 U637 ( .A1(G49), .A2(n791), .ZN(n565) );
  NAND2_X1 U638 ( .A1(G74), .A2(G651), .ZN(n564) );
  NAND2_X1 U639 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U640 ( .A1(n789), .A2(n566), .ZN(n569) );
  NAND2_X1 U641 ( .A1(n567), .A2(G87), .ZN(n568) );
  NAND2_X1 U642 ( .A1(n569), .A2(n568), .ZN(G288) );
  NAND2_X1 U643 ( .A1(G73), .A2(n786), .ZN(n570) );
  XNOR2_X1 U644 ( .A(n570), .B(KEYINPUT2), .ZN(n577) );
  NAND2_X1 U645 ( .A1(G86), .A2(n785), .ZN(n572) );
  NAND2_X1 U646 ( .A1(G61), .A2(n789), .ZN(n571) );
  NAND2_X1 U647 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n791), .A2(G48), .ZN(n573) );
  XOR2_X1 U649 ( .A(KEYINPUT76), .B(n573), .Z(n574) );
  NOR2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U651 ( .A1(n577), .A2(n576), .ZN(G305) );
  NAND2_X1 U652 ( .A1(G101), .A2(n879), .ZN(n579) );
  NAND2_X1 U653 ( .A1(G113), .A2(n875), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U655 ( .A1(G125), .A2(n876), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n595) );
  BUF_X1 U658 ( .A(n595), .Z(G160) );
  NAND2_X1 U659 ( .A1(G85), .A2(n785), .ZN(n589) );
  NAND2_X1 U660 ( .A1(G72), .A2(n786), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n789), .A2(G60), .ZN(n590) );
  XOR2_X1 U663 ( .A(KEYINPUT66), .B(n590), .Z(n591) );
  NOR2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n791), .A2(G47), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(G290) );
  NOR2_X2 U667 ( .A1(G164), .A2(G1384), .ZN(n722) );
  INV_X1 U668 ( .A(KEYINPUT64), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G2072), .A2(n638), .ZN(n598) );
  XNOR2_X1 U670 ( .A(n598), .B(KEYINPUT27), .ZN(n600) );
  XOR2_X1 U671 ( .A(KEYINPUT90), .B(G1956), .Z(n1008) );
  NOR2_X1 U672 ( .A1(n640), .A2(n1008), .ZN(n599) );
  NOR2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n602) );
  INV_X1 U674 ( .A(KEYINPUT91), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n602), .B(n601), .ZN(n604) );
  INV_X1 U676 ( .A(G299), .ZN(n976) );
  NOR2_X1 U677 ( .A1(n604), .A2(n976), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n603), .B(KEYINPUT28), .ZN(n635) );
  NAND2_X1 U679 ( .A1(n976), .A2(n604), .ZN(n633) );
  NAND2_X1 U680 ( .A1(n640), .A2(G1996), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT26), .ZN(n617) );
  INV_X1 U682 ( .A(n638), .ZN(n649) );
  NAND2_X1 U683 ( .A1(n785), .A2(G81), .ZN(n606) );
  XNOR2_X1 U684 ( .A(n606), .B(KEYINPUT12), .ZN(n608) );
  NAND2_X1 U685 ( .A1(G68), .A2(n786), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(n610) );
  XOR2_X1 U687 ( .A(KEYINPUT68), .B(KEYINPUT13), .Z(n609) );
  XNOR2_X1 U688 ( .A(n610), .B(n609), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n789), .A2(G56), .ZN(n611) );
  XOR2_X1 U690 ( .A(KEYINPUT14), .B(n611), .Z(n612) );
  NOR2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n791), .A2(G43), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n984) );
  NOR2_X1 U694 ( .A1(n517), .A2(n984), .ZN(n616) );
  NAND2_X1 U695 ( .A1(G92), .A2(n785), .ZN(n619) );
  NAND2_X1 U696 ( .A1(G66), .A2(n789), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n624) );
  NAND2_X1 U698 ( .A1(G79), .A2(n786), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G54), .A2(n791), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U701 ( .A(KEYINPUT70), .B(n622), .ZN(n623) );
  NOR2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(KEYINPUT15), .ZN(n968) );
  NAND2_X1 U704 ( .A1(G2067), .A2(n640), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n649), .A2(G1348), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n968), .A2(n629), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n968), .A2(n629), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n632) );
  OR2_X2 U710 ( .A1(n635), .A2(n634), .ZN(n637) );
  NOR2_X1 U711 ( .A1(n638), .A2(G1961), .ZN(n639) );
  XOR2_X1 U712 ( .A(KEYINPUT88), .B(n639), .Z(n642) );
  XNOR2_X1 U713 ( .A(KEYINPUT25), .B(G2078), .ZN(n951) );
  NAND2_X1 U714 ( .A1(n640), .A2(n951), .ZN(n641) );
  NAND2_X1 U715 ( .A1(n642), .A2(n641), .ZN(n653) );
  NAND2_X1 U716 ( .A1(G171), .A2(n653), .ZN(n643) );
  XOR2_X1 U717 ( .A(KEYINPUT89), .B(n643), .Z(n644) );
  NAND2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n660) );
  NAND2_X1 U719 ( .A1(n646), .A2(G8), .ZN(n648) );
  NOR2_X1 U720 ( .A1(n649), .A2(G2084), .ZN(n672) );
  NOR2_X1 U721 ( .A1(n675), .A2(n672), .ZN(n650) );
  NOR2_X1 U722 ( .A1(n652), .A2(G168), .ZN(n656) );
  NOR2_X1 U723 ( .A1(G171), .A2(n653), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n654), .B(KEYINPUT92), .ZN(n655) );
  INV_X1 U725 ( .A(KEYINPUT31), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n660), .A2(n659), .ZN(n673) );
  AND2_X1 U727 ( .A1(G286), .A2(G8), .ZN(n661) );
  NAND2_X1 U728 ( .A1(n673), .A2(n661), .ZN(n670) );
  INV_X1 U729 ( .A(G8), .ZN(n668) );
  NOR2_X1 U730 ( .A1(n649), .A2(G2090), .ZN(n662) );
  XOR2_X1 U731 ( .A(KEYINPUT93), .B(n662), .Z(n664) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n701), .ZN(n663) );
  NOR2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U734 ( .A(n665), .B(KEYINPUT94), .ZN(n666) );
  NAND2_X1 U735 ( .A1(n666), .A2(G303), .ZN(n667) );
  OR2_X1 U736 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U737 ( .A(n671), .B(KEYINPUT32), .ZN(n679) );
  NAND2_X1 U738 ( .A1(G8), .A2(n672), .ZN(n677) );
  INV_X1 U739 ( .A(n673), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n697) );
  NOR2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n685) );
  NOR2_X1 U744 ( .A1(G1971), .A2(G303), .ZN(n680) );
  NOR2_X1 U745 ( .A1(n685), .A2(n680), .ZN(n975) );
  NAND2_X1 U746 ( .A1(n697), .A2(n975), .ZN(n681) );
  XNOR2_X1 U747 ( .A(KEYINPUT95), .B(n681), .ZN(n683) );
  NAND2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n974) );
  INV_X1 U749 ( .A(n701), .ZN(n693) );
  NAND2_X1 U750 ( .A1(n974), .A2(n693), .ZN(n682) );
  NOR2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U752 ( .A1(n684), .A2(KEYINPUT33), .ZN(n689) );
  NAND2_X1 U753 ( .A1(KEYINPUT33), .A2(n685), .ZN(n686) );
  NOR2_X1 U754 ( .A1(n701), .A2(n686), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n687), .B(KEYINPUT96), .ZN(n688) );
  NOR2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U757 ( .A(n690), .B(KEYINPUT97), .ZN(n691) );
  XNOR2_X1 U758 ( .A(G1981), .B(G305), .ZN(n970) );
  NOR2_X1 U759 ( .A1(n691), .A2(n970), .ZN(n705) );
  NOR2_X1 U760 ( .A1(G1981), .A2(G305), .ZN(n692) );
  XNOR2_X1 U761 ( .A(KEYINPUT24), .B(n692), .ZN(n694) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n703) );
  NOR2_X1 U763 ( .A1(G2090), .A2(G303), .ZN(n695) );
  XNOR2_X1 U764 ( .A(n695), .B(KEYINPUT98), .ZN(n696) );
  NAND2_X1 U765 ( .A1(n696), .A2(G8), .ZN(n698) );
  NAND2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U767 ( .A(KEYINPUT99), .B(n699), .Z(n700) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n739) );
  NAND2_X1 U771 ( .A1(G95), .A2(n879), .ZN(n707) );
  NAND2_X1 U772 ( .A1(G131), .A2(n880), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U774 ( .A1(G107), .A2(n875), .ZN(n709) );
  NAND2_X1 U775 ( .A1(G119), .A2(n876), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n866) );
  XNOR2_X1 U778 ( .A(KEYINPUT85), .B(G1991), .ZN(n947) );
  NOR2_X1 U779 ( .A1(n866), .A2(n947), .ZN(n720) );
  NAND2_X1 U780 ( .A1(G117), .A2(n875), .ZN(n713) );
  NAND2_X1 U781 ( .A1(G141), .A2(n880), .ZN(n712) );
  NAND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n879), .A2(G105), .ZN(n714) );
  XOR2_X1 U784 ( .A(KEYINPUT38), .B(n714), .Z(n715) );
  NOR2_X1 U785 ( .A1(n716), .A2(n715), .ZN(n718) );
  NAND2_X1 U786 ( .A1(n876), .A2(G129), .ZN(n717) );
  NAND2_X1 U787 ( .A1(n718), .A2(n717), .ZN(n888) );
  AND2_X1 U788 ( .A1(G1996), .A2(n888), .ZN(n719) );
  NOR2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n927) );
  INV_X1 U790 ( .A(n721), .ZN(n723) );
  NOR2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U792 ( .A(KEYINPUT81), .B(n724), .Z(n755) );
  INV_X1 U793 ( .A(n755), .ZN(n741) );
  NOR2_X1 U794 ( .A1(n927), .A2(n741), .ZN(n747) );
  XOR2_X1 U795 ( .A(n747), .B(KEYINPUT86), .Z(n737) );
  XNOR2_X1 U796 ( .A(G2067), .B(KEYINPUT37), .ZN(n753) );
  NAND2_X1 U797 ( .A1(n875), .A2(G116), .ZN(n725) );
  XOR2_X1 U798 ( .A(KEYINPUT83), .B(n725), .Z(n727) );
  NAND2_X1 U799 ( .A1(n876), .A2(G128), .ZN(n726) );
  NAND2_X1 U800 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U801 ( .A(n728), .B(KEYINPUT35), .ZN(n733) );
  NAND2_X1 U802 ( .A1(G104), .A2(n879), .ZN(n730) );
  NAND2_X1 U803 ( .A1(G140), .A2(n880), .ZN(n729) );
  NAND2_X1 U804 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U805 ( .A(KEYINPUT34), .B(n731), .Z(n732) );
  NAND2_X1 U806 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U807 ( .A(n734), .B(KEYINPUT36), .Z(n864) );
  OR2_X1 U808 ( .A1(n753), .A2(n864), .ZN(n735) );
  XNOR2_X1 U809 ( .A(KEYINPUT84), .B(n735), .ZN(n928) );
  NOR2_X1 U810 ( .A1(n928), .A2(n741), .ZN(n751) );
  INV_X1 U811 ( .A(n751), .ZN(n736) );
  NAND2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U813 ( .A(n740), .B(KEYINPUT100), .ZN(n744) );
  XOR2_X1 U814 ( .A(G1986), .B(G290), .Z(n987) );
  NOR2_X1 U815 ( .A1(n987), .A2(n741), .ZN(n742) );
  XOR2_X1 U816 ( .A(KEYINPUT82), .B(n742), .Z(n743) );
  NAND2_X1 U817 ( .A1(n744), .A2(n743), .ZN(n759) );
  NOR2_X1 U818 ( .A1(G1996), .A2(n888), .ZN(n922) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n745) );
  AND2_X1 U820 ( .A1(n947), .A2(n866), .ZN(n932) );
  NOR2_X1 U821 ( .A1(n745), .A2(n932), .ZN(n746) );
  NOR2_X1 U822 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U823 ( .A1(n922), .A2(n748), .ZN(n749) );
  XOR2_X1 U824 ( .A(KEYINPUT39), .B(n749), .Z(n750) );
  NOR2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U826 ( .A(KEYINPUT101), .B(n752), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n753), .A2(n864), .ZN(n925) );
  NAND2_X1 U828 ( .A1(n754), .A2(n925), .ZN(n756) );
  NAND2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U830 ( .A(n757), .B(KEYINPUT102), .ZN(n758) );
  NAND2_X1 U831 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U832 ( .A(n760), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U834 ( .A(G57), .ZN(G237) );
  INV_X1 U835 ( .A(G132), .ZN(G219) );
  INV_X1 U836 ( .A(G82), .ZN(G220) );
  NAND2_X1 U837 ( .A1(G7), .A2(G661), .ZN(n761) );
  XNOR2_X1 U838 ( .A(n761), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U839 ( .A(G223), .ZN(n822) );
  NAND2_X1 U840 ( .A1(n822), .A2(G567), .ZN(n762) );
  XOR2_X1 U841 ( .A(KEYINPUT11), .B(n762), .Z(G234) );
  INV_X1 U842 ( .A(G860), .ZN(n769) );
  OR2_X1 U843 ( .A1(n984), .A2(n769), .ZN(G153) );
  XNOR2_X1 U844 ( .A(G171), .B(KEYINPUT69), .ZN(G301) );
  NAND2_X1 U845 ( .A1(G868), .A2(G301), .ZN(n764) );
  INV_X1 U846 ( .A(G868), .ZN(n766) );
  NAND2_X1 U847 ( .A1(n968), .A2(n766), .ZN(n763) );
  NAND2_X1 U848 ( .A1(n764), .A2(n763), .ZN(G284) );
  NOR2_X1 U849 ( .A1(G868), .A2(G299), .ZN(n765) );
  XOR2_X1 U850 ( .A(KEYINPUT73), .B(n765), .Z(n768) );
  NOR2_X1 U851 ( .A1(G286), .A2(n766), .ZN(n767) );
  NOR2_X1 U852 ( .A1(n768), .A2(n767), .ZN(G297) );
  NAND2_X1 U853 ( .A1(n769), .A2(G559), .ZN(n770) );
  INV_X1 U854 ( .A(n968), .ZN(n895) );
  NAND2_X1 U855 ( .A1(n770), .A2(n895), .ZN(n771) );
  XNOR2_X1 U856 ( .A(n771), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U857 ( .A1(G868), .A2(n984), .ZN(n774) );
  NAND2_X1 U858 ( .A1(n895), .A2(G868), .ZN(n772) );
  NOR2_X1 U859 ( .A1(G559), .A2(n772), .ZN(n773) );
  NOR2_X1 U860 ( .A1(n774), .A2(n773), .ZN(G282) );
  XOR2_X1 U861 ( .A(G2100), .B(KEYINPUT74), .Z(n783) );
  NAND2_X1 U862 ( .A1(G111), .A2(n875), .ZN(n776) );
  NAND2_X1 U863 ( .A1(G135), .A2(n880), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n876), .A2(G123), .ZN(n777) );
  XOR2_X1 U866 ( .A(KEYINPUT18), .B(n777), .Z(n778) );
  NOR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n879), .A2(G99), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n929) );
  XOR2_X1 U870 ( .A(G2096), .B(n929), .Z(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(G156) );
  NAND2_X1 U872 ( .A1(G559), .A2(n895), .ZN(n784) );
  XNOR2_X1 U873 ( .A(n784), .B(n984), .ZN(n805) );
  NOR2_X1 U874 ( .A1(n805), .A2(G860), .ZN(n796) );
  NAND2_X1 U875 ( .A1(G93), .A2(n785), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G80), .A2(n786), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n795) );
  NAND2_X1 U878 ( .A1(G67), .A2(n789), .ZN(n790) );
  XOR2_X1 U879 ( .A(KEYINPUT75), .B(n790), .Z(n793) );
  NAND2_X1 U880 ( .A1(n791), .A2(G55), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n798) );
  XNOR2_X1 U883 ( .A(n796), .B(n798), .ZN(G145) );
  NOR2_X1 U884 ( .A1(G868), .A2(n798), .ZN(n797) );
  XNOR2_X1 U885 ( .A(n797), .B(KEYINPUT79), .ZN(n808) );
  XNOR2_X1 U886 ( .A(n976), .B(G305), .ZN(n799) );
  XOR2_X1 U887 ( .A(n799), .B(n798), .Z(n800) );
  XNOR2_X1 U888 ( .A(KEYINPUT19), .B(n800), .ZN(n802) );
  XNOR2_X1 U889 ( .A(G288), .B(KEYINPUT78), .ZN(n801) );
  XNOR2_X1 U890 ( .A(n802), .B(n801), .ZN(n803) );
  XNOR2_X1 U891 ( .A(n803), .B(G303), .ZN(n804) );
  XNOR2_X1 U892 ( .A(n804), .B(G290), .ZN(n892) );
  XNOR2_X1 U893 ( .A(n892), .B(n805), .ZN(n806) );
  NAND2_X1 U894 ( .A1(G868), .A2(n806), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n808), .A2(n807), .ZN(G295) );
  NAND2_X1 U896 ( .A1(G2078), .A2(G2084), .ZN(n809) );
  XOR2_X1 U897 ( .A(KEYINPUT20), .B(n809), .Z(n810) );
  NAND2_X1 U898 ( .A1(G2090), .A2(n810), .ZN(n811) );
  XNOR2_X1 U899 ( .A(KEYINPUT21), .B(n811), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n812), .A2(G2072), .ZN(n813) );
  XNOR2_X1 U901 ( .A(KEYINPUT80), .B(n813), .ZN(G158) );
  XNOR2_X1 U902 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U903 ( .A1(G220), .A2(G219), .ZN(n814) );
  XOR2_X1 U904 ( .A(KEYINPUT22), .B(n814), .Z(n815) );
  NOR2_X1 U905 ( .A1(G218), .A2(n815), .ZN(n816) );
  NAND2_X1 U906 ( .A1(G96), .A2(n816), .ZN(n826) );
  NAND2_X1 U907 ( .A1(n826), .A2(G2106), .ZN(n820) );
  NAND2_X1 U908 ( .A1(G69), .A2(G120), .ZN(n817) );
  NOR2_X1 U909 ( .A1(G237), .A2(n817), .ZN(n818) );
  NAND2_X1 U910 ( .A1(G108), .A2(n818), .ZN(n827) );
  NAND2_X1 U911 ( .A1(n827), .A2(G567), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n828) );
  NAND2_X1 U913 ( .A1(G661), .A2(G483), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n828), .A2(n821), .ZN(n825) );
  NAND2_X1 U915 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n822), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U918 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(G188) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n827), .A2(n826), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  INV_X1 U927 ( .A(n828), .ZN(G319) );
  XOR2_X1 U928 ( .A(G2678), .B(G2090), .Z(n830) );
  XNOR2_X1 U929 ( .A(G2072), .B(G2084), .ZN(n829) );
  XNOR2_X1 U930 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U931 ( .A(n831), .B(G2096), .Z(n833) );
  XNOR2_X1 U932 ( .A(G2078), .B(G2067), .ZN(n832) );
  XNOR2_X1 U933 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U934 ( .A(G2100), .B(KEYINPUT105), .Z(n835) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U937 ( .A(n837), .B(n836), .Z(G227) );
  XOR2_X1 U938 ( .A(G1981), .B(G1956), .Z(n839) );
  XNOR2_X1 U939 ( .A(G1966), .B(G1961), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n849) );
  XOR2_X1 U941 ( .A(KEYINPUT106), .B(KEYINPUT41), .Z(n841) );
  XNOR2_X1 U942 ( .A(G1991), .B(KEYINPUT107), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U944 ( .A(G1986), .B(G1976), .Z(n843) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1971), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U947 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U948 ( .A(KEYINPUT108), .B(G2474), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(G229) );
  NAND2_X1 U951 ( .A1(G124), .A2(n876), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U953 ( .A1(n875), .A2(G112), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U955 ( .A1(G100), .A2(n879), .ZN(n854) );
  NAND2_X1 U956 ( .A1(G136), .A2(n880), .ZN(n853) );
  NAND2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U958 ( .A1(n856), .A2(n855), .ZN(G162) );
  NAND2_X1 U959 ( .A1(G103), .A2(n879), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G139), .A2(n880), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G115), .A2(n875), .ZN(n860) );
  NAND2_X1 U963 ( .A1(G127), .A2(n876), .ZN(n859) );
  NAND2_X1 U964 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U965 ( .A(KEYINPUT47), .B(n861), .Z(n862) );
  NOR2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n915) );
  XOR2_X1 U967 ( .A(n864), .B(n915), .Z(n865) );
  XNOR2_X1 U968 ( .A(n865), .B(G162), .ZN(n869) );
  XNOR2_X1 U969 ( .A(G160), .B(G164), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U971 ( .A(n869), .B(n868), .Z(n874) );
  XOR2_X1 U972 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n871) );
  XNOR2_X1 U973 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n870) );
  XNOR2_X1 U974 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U975 ( .A(KEYINPUT48), .B(n872), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n890) );
  NAND2_X1 U977 ( .A1(G118), .A2(n875), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G130), .A2(n876), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U980 ( .A1(G106), .A2(n879), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G142), .A2(n880), .ZN(n881) );
  NAND2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U983 ( .A(n883), .B(KEYINPUT45), .Z(n884) );
  NOR2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n886), .B(n929), .ZN(n887) );
  XOR2_X1 U986 ( .A(n888), .B(n887), .Z(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U988 ( .A1(G37), .A2(n891), .ZN(G395) );
  XOR2_X1 U989 ( .A(G171), .B(n892), .Z(n893) );
  XNOR2_X1 U990 ( .A(n984), .B(n893), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n896), .B(G286), .ZN(n897) );
  NOR2_X1 U993 ( .A1(G37), .A2(n897), .ZN(G397) );
  XNOR2_X1 U994 ( .A(G2451), .B(G2443), .ZN(n907) );
  XOR2_X1 U995 ( .A(G2446), .B(G2430), .Z(n899) );
  XNOR2_X1 U996 ( .A(KEYINPUT104), .B(G2438), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U998 ( .A(G2435), .B(G2454), .Z(n901) );
  XNOR2_X1 U999 ( .A(G1341), .B(G1348), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1001 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U1002 ( .A(KEYINPUT103), .B(G2427), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(n908), .A2(G14), .ZN(n914) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n914), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n914), .ZN(G401) );
  XNOR2_X1 U1015 ( .A(G2072), .B(n915), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(G164), .B(G2078), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(KEYINPUT116), .ZN(n917) );
  NAND2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1019 ( .A(n919), .B(KEYINPUT50), .ZN(n920) );
  XOR2_X1 U1020 ( .A(KEYINPUT117), .B(n920), .Z(n941) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1023 ( .A(KEYINPUT51), .B(n923), .Z(n924) );
  XNOR2_X1 U1024 ( .A(n924), .B(KEYINPUT114), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n938) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(G160), .B(G2084), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT112), .B(n933), .Z(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(n936), .B(KEYINPUT113), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(KEYINPUT115), .B(n939), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(n942), .B(KEYINPUT118), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(n943), .B(KEYINPUT52), .ZN(n945) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n946), .A2(G29), .ZN(n997) );
  XNOR2_X1 U1041 ( .A(G2072), .B(G33), .ZN(n949) );
  XOR2_X1 U1042 ( .A(n947), .B(G25), .Z(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n958) );
  XOR2_X1 U1044 ( .A(G2067), .B(G26), .Z(n950) );
  NAND2_X1 U1045 ( .A1(n950), .A2(G28), .ZN(n956) );
  XOR2_X1 U1046 ( .A(n951), .B(G27), .Z(n953) );
  XNOR2_X1 U1047 ( .A(G32), .B(G1996), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(n954), .B(KEYINPUT119), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(n959), .B(KEYINPUT53), .ZN(n962) );
  XOR2_X1 U1053 ( .A(G2084), .B(G34), .Z(n960) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n960), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(G35), .B(G2090), .ZN(n963) );
  NOR2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1058 ( .A(KEYINPUT55), .B(n965), .Z(n966) );
  NOR2_X1 U1059 ( .A1(G29), .A2(n966), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(KEYINPUT120), .B(n967), .ZN(n995) );
  XOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .Z(n992) );
  XNOR2_X1 U1062 ( .A(n968), .B(G1348), .ZN(n973) );
  XOR2_X1 U1063 ( .A(G1966), .B(G168), .Z(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT57), .B(n971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n983) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(n976), .B(G1956), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(G1971), .A2(G303), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1072 ( .A(KEYINPUT121), .B(n981), .Z(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n990) );
  XOR2_X1 U1074 ( .A(G171), .B(G1961), .Z(n986) );
  XNOR2_X1 U1075 ( .A(n984), .B(G1341), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(KEYINPUT122), .B(n993), .ZN(n994) );
  NOR2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1082 ( .A1(n997), .A2(n996), .ZN(n1027) );
  XNOR2_X1 U1083 ( .A(G1971), .B(G22), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(G24), .B(G1986), .ZN(n998) );
  NOR2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XOR2_X1 U1086 ( .A(G1976), .B(G23), .Z(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XOR2_X1 U1088 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n1002) );
  XNOR2_X1 U1089 ( .A(n1003), .B(n1002), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G21), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(G5), .B(G1961), .ZN(n1004) );
  NOR2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1020) );
  XNOR2_X1 U1094 ( .A(n1008), .B(G20), .ZN(n1016) );
  XOR2_X1 U1095 ( .A(G1981), .B(G6), .Z(n1011) );
  XOR2_X1 U1096 ( .A(G19), .B(KEYINPUT124), .Z(n1009) );
  XNOR2_X1 U1097 ( .A(G1341), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(KEYINPUT59), .B(G1348), .Z(n1012) );
  XNOR2_X1 U1100 ( .A(G4), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(n1017), .B(KEYINPUT60), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(n1018), .B(KEYINPUT125), .Z(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1021), .Z(n1022) );
  XNOR2_X1 U1107 ( .A(n1022), .B(KEYINPUT127), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(G16), .B(KEYINPUT123), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(G11), .A2(n1025), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(n1028), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
  INV_X1 U1114 ( .A(G303), .ZN(G166) );
endmodule

