//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT65), .Z(new_n212));
  OR2_X1    g0012(.A1(new_n212), .A2(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT66), .ZN(new_n217));
  NOR2_X1   g0017(.A1(G58), .A2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n213), .A2(new_n214), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT67), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT68), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G107), .A2(G264), .ZN(new_n231));
  NAND4_X1  g0031(.A1(new_n228), .A2(new_n229), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n209), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT69), .Z(new_n235));
  OAI211_X1 g0035(.A(new_n224), .B(new_n235), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT70), .Z(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G226), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G223), .A3(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G222), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n259), .B1(new_n226), .B2(new_n258), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT71), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(new_n269), .A3(G274), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT71), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n264), .A2(new_n268), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(G226), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n265), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G190), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n208), .A2(G33), .B1(G1), .B2(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n203), .A2(G20), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT8), .B(G58), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n207), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n284), .A2(new_n286), .B1(G150), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n281), .B1(new_n282), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G13), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(G1), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G50), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n281), .B1(G1), .B2(new_n207), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(G50), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(KEYINPUT9), .ZN(new_n298));
  AOI211_X1 g0098(.A(new_n280), .B(new_n298), .C1(G200), .C2(new_n278), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(KEYINPUT9), .ZN(new_n300));
  XOR2_X1   g0100(.A(new_n300), .B(KEYINPUT72), .Z(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(KEYINPUT73), .A3(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(KEYINPUT73), .B1(new_n302), .B2(KEYINPUT10), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n304), .A2(new_n305), .B1(KEYINPUT10), .B2(new_n302), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n278), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(G169), .B2(new_n278), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(new_n297), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G68), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n291), .A2(G20), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT12), .ZN(new_n315));
  INV_X1    g0115(.A(new_n281), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n313), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n226), .B2(new_n285), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XOR2_X1   g0119(.A(KEYINPUT76), .B(KEYINPUT11), .Z(new_n320));
  OAI221_X1 g0120(.A(new_n315), .B1(new_n295), .B2(new_n313), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n319), .A2(new_n320), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT77), .ZN(new_n324));
  OAI211_X1 g0124(.A(G1), .B(G13), .C1(new_n255), .C2(new_n266), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(G238), .A3(new_n271), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n274), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT74), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n258), .A2(G232), .A3(G1698), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n258), .A2(G226), .A3(new_n260), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G97), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n264), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n274), .A2(KEYINPUT74), .A3(new_n326), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n329), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT13), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n329), .A2(new_n334), .A3(new_n335), .A4(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(G179), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  INV_X1    g0141(.A(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n341), .B1(new_n343), .B2(new_n339), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI211_X1 g0146(.A(KEYINPUT14), .B(new_n341), .C1(new_n343), .C2(new_n339), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n324), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT80), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n325), .A2(new_n350), .A3(G232), .A4(new_n271), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n274), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(KEYINPUT3), .A2(G33), .ZN(new_n353));
  NOR2_X1   g0153(.A1(KEYINPUT3), .A2(G33), .ZN(new_n354));
  OAI211_X1 g0154(.A(G226), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G87), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT79), .B1(new_n255), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT79), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(G33), .A3(G87), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(G223), .B(new_n260), .C1(new_n353), .C2(new_n354), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n355), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n264), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n325), .A2(G232), .A3(new_n271), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT80), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n352), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n341), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n366), .B2(G179), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT78), .ZN(new_n371));
  XNOR2_X1  g0171(.A(G58), .B(G68), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(G20), .ZN(new_n373));
  AND2_X1   g0173(.A1(G58), .A2(G68), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n371), .B(G20), .C1(new_n374), .C2(new_n218), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  INV_X1    g0177(.A(new_n287), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n373), .A2(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n256), .A2(new_n207), .A3(new_n257), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n353), .A2(new_n354), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n313), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n370), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT7), .B1(new_n383), .B2(new_n207), .ZN(new_n387));
  NOR4_X1   g0187(.A1(new_n353), .A2(new_n354), .A3(new_n381), .A4(G20), .ZN(new_n388));
  OAI21_X1  g0188(.A(G68), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n378), .A2(new_n377), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n374), .B2(new_n218), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT78), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n392), .B2(new_n375), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n393), .A3(KEYINPUT16), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n386), .A2(new_n316), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n293), .A2(new_n284), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n295), .B2(new_n284), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n369), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G200), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n362), .A2(new_n264), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n365), .A2(new_n274), .A3(new_n351), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n352), .A2(new_n279), .A3(new_n363), .A4(new_n365), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(new_n395), .A3(new_n398), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n343), .A2(new_n339), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G200), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n337), .A2(G190), .A3(new_n339), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n323), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n258), .A2(G238), .A3(G1698), .ZN(new_n417));
  INV_X1    g0217(.A(G107), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n417), .B1(new_n418), .B2(new_n258), .C1(new_n261), .C2(new_n241), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n264), .ZN(new_n420));
  INV_X1    g0220(.A(new_n225), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n275), .B1(new_n421), .B2(new_n276), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G169), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n307), .B2(new_n423), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT15), .B(G87), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n427), .A2(new_n286), .B1(G20), .B2(G77), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n378), .B2(new_n283), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n316), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n293), .A2(new_n226), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n430), .B(new_n431), .C1(new_n226), .C2(new_n295), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n423), .A2(G190), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n403), .B2(new_n423), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n433), .B1(new_n435), .B2(new_n432), .ZN(new_n436));
  OR4_X1    g0236(.A1(new_n349), .A2(new_n411), .A3(new_n416), .A4(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n312), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n427), .A2(new_n292), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n258), .A2(new_n207), .ZN(new_n440));
  OR2_X1    g0240(.A1(KEYINPUT81), .A2(G97), .ZN(new_n441));
  NAND2_X1  g0241(.A1(KEYINPUT81), .A2(G97), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n285), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n440), .A2(new_n313), .B1(new_n443), .B2(KEYINPUT19), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n441), .A2(new_n356), .A3(new_n418), .A4(new_n442), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT19), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n207), .B1(new_n332), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT84), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(KEYINPUT84), .A3(new_n447), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n444), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT85), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n281), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n383), .A2(G20), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n441), .A2(new_n442), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n286), .ZN(new_n456));
  AOI22_X1  g0256(.A1(G68), .A2(new_n454), .B1(new_n456), .B2(new_n446), .ZN(new_n457));
  INV_X1    g0257(.A(new_n450), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n457), .B1(new_n458), .B2(new_n448), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT85), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n439), .B1(new_n453), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n206), .A2(G45), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G250), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n267), .A2(G1), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G274), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n264), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n258), .A2(G238), .A3(new_n260), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n258), .A2(G244), .A3(G1698), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G116), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n466), .B1(new_n470), .B2(new_n264), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n471), .A2(new_n403), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n281), .B(new_n292), .C1(G1), .C2(new_n255), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G87), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n264), .ZN(new_n476));
  INV_X1    g0276(.A(new_n466), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(G190), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT86), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n471), .A2(new_n480), .A3(G190), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n461), .A2(new_n472), .A3(new_n475), .A4(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT87), .ZN(new_n484));
  INV_X1    g0284(.A(new_n439), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n474), .A2(new_n427), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n316), .B1(new_n459), .B2(KEYINPUT85), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n451), .A2(new_n452), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n485), .B(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n471), .A2(G179), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n341), .B2(new_n471), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n483), .A2(new_n484), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n484), .B1(new_n483), .B2(new_n492), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT82), .B1(new_n292), .B2(G97), .ZN(new_n496));
  OR3_X1    g0296(.A1(new_n292), .A2(KEYINPUT82), .A3(G97), .ZN(new_n497));
  INV_X1    g0297(.A(G97), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n496), .B(new_n497), .C1(new_n473), .C2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT6), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n498), .A2(new_n418), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G97), .A2(G107), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n455), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n418), .A2(KEYINPUT6), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(G20), .B1(G77), .B2(new_n287), .ZN(new_n507));
  OAI21_X1  g0307(.A(G107), .B1(new_n387), .B2(new_n388), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n499), .B1(new_n509), .B2(new_n316), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n266), .ZN(new_n512));
  NAND2_X1  g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n462), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G274), .ZN(new_n515));
  INV_X1    g0315(.A(new_n513), .ZN(new_n516));
  NOR2_X1   g0316(.A1(KEYINPUT5), .A2(G41), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n464), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n325), .ZN(new_n519));
  INV_X1    g0319(.A(G257), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(G244), .B1(new_n353), .B2(new_n354), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT4), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n522), .A2(new_n523), .B1(G33), .B2(G283), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n258), .A2(KEYINPUT4), .A3(G244), .A4(new_n260), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n523), .B1(new_n258), .B2(G250), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n524), .B(new_n525), .C1(new_n260), .C2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n521), .B1(new_n527), .B2(new_n264), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G169), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(G179), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n510), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI211_X1 g0332(.A(G190), .B(new_n521), .C1(new_n527), .C2(new_n264), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n524), .A2(new_n525), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n526), .A2(new_n260), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n264), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n521), .ZN(new_n537));
  AOI21_X1  g0337(.A(G200), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n510), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT83), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT83), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n510), .B(new_n541), .C1(new_n533), .C2(new_n538), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n532), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n258), .A2(G264), .A3(G1698), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n258), .A2(G257), .A3(new_n260), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n383), .A2(G303), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n264), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n514), .A2(new_n264), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n549), .A2(G270), .B1(G274), .B2(new_n514), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G169), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT21), .ZN(new_n553));
  OAI22_X1  g0353(.A1(new_n552), .A2(new_n553), .B1(new_n307), .B2(new_n551), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n455), .A2(new_n255), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G283), .ZN(new_n556));
  AOI21_X1  g0356(.A(G20), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(G116), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n207), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n316), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT20), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(KEYINPUT20), .B(new_n316), .C1(new_n557), .C2(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n473), .A2(G116), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n292), .A2(new_n558), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n554), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n562), .A2(new_n563), .B1(new_n566), .B2(new_n565), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n553), .B1(new_n570), .B2(new_n552), .ZN(new_n571));
  AOI21_X1  g0371(.A(G200), .B1(new_n548), .B2(new_n550), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n551), .A2(G190), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n569), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n258), .A2(G250), .A3(new_n260), .ZN(new_n576));
  OAI211_X1 g0376(.A(G257), .B(G1698), .C1(new_n353), .C2(new_n354), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G294), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n264), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n518), .A2(G264), .A3(new_n325), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n580), .A2(new_n515), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT89), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n549), .A2(KEYINPUT89), .A3(G264), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n580), .A2(new_n515), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n582), .A2(new_n279), .B1(new_n586), .B2(new_n403), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n473), .A2(new_n418), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n291), .A2(G20), .A3(new_n418), .ZN(new_n589));
  XNOR2_X1  g0389(.A(new_n589), .B(KEYINPUT25), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n207), .B(G87), .C1(new_n353), .C2(new_n354), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT22), .ZN(new_n593));
  OR3_X1    g0393(.A1(new_n469), .A2(KEYINPUT88), .A3(G20), .ZN(new_n594));
  OAI21_X1  g0394(.A(KEYINPUT88), .B1(new_n469), .B2(G20), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT23), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n207), .B2(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n418), .A2(KEYINPUT23), .A3(G20), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n594), .A2(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n593), .A2(KEYINPUT24), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n316), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT24), .B1(new_n593), .B2(new_n599), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n591), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n587), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n586), .A2(new_n307), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT90), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT90), .B1(new_n586), .B2(new_n307), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n580), .A2(new_n515), .A3(new_n581), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G169), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n604), .B1(new_n611), .B2(new_n603), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n543), .A2(new_n575), .A3(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n438), .A2(new_n495), .A3(new_n613), .ZN(G372));
  NAND4_X1  g0414(.A1(new_n461), .A2(new_n472), .A3(new_n475), .A4(new_n478), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT26), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n615), .A2(new_n492), .A3(new_n616), .A4(new_n532), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n543), .B1(new_n603), .B2(new_n587), .ZN(new_n618));
  INV_X1    g0418(.A(new_n603), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n605), .A2(new_n606), .B1(G169), .B2(new_n609), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(new_n608), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n569), .A2(new_n571), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n615), .B(new_n492), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n492), .B(new_n617), .C1(new_n618), .C2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n495), .A2(new_n532), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(KEYINPUT26), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n438), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n433), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n349), .B1(new_n415), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n410), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n402), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n310), .B1(new_n633), .B2(new_n306), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n629), .A2(new_n634), .ZN(G369));
  INV_X1    g0435(.A(new_n291), .ZN(new_n636));
  OR3_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .A3(G20), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT27), .B1(new_n636), .B2(G20), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(G343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n612), .B1(new_n619), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n621), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n643), .B1(new_n644), .B2(new_n642), .ZN(new_n645));
  XNOR2_X1  g0445(.A(new_n645), .B(KEYINPUT91), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n570), .A2(new_n642), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n575), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n622), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n647), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G330), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n649), .A2(new_n641), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n646), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n641), .B(KEYINPUT92), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n621), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n654), .A2(new_n656), .A3(new_n658), .ZN(G399));
  INV_X1    g0459(.A(new_n210), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(G41), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n445), .A2(G116), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n661), .A2(new_n206), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT93), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT93), .B1(new_n661), .B2(new_n221), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n613), .A2(new_n495), .A3(new_n657), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n548), .A2(new_n550), .A3(G179), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(new_n471), .A4(new_n528), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND4_X1   g0475(.A1(new_n471), .A2(new_n580), .A3(new_n584), .A4(new_n585), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(KEYINPUT30), .A3(new_n528), .A4(new_n671), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n471), .A2(G179), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n529), .A2(new_n678), .A3(new_n586), .A4(new_n551), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(KEYINPUT31), .B1(new_n680), .B2(new_n641), .ZN(new_n681));
  INV_X1    g0481(.A(new_n657), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(KEYINPUT31), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n652), .B1(new_n670), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n682), .B1(new_n625), .B2(new_n627), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g0487(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n626), .A2(KEYINPUT26), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n615), .A2(new_n492), .ZN(new_n691));
  INV_X1    g0491(.A(new_n532), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT26), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n492), .B(new_n693), .C1(new_n618), .C2(new_n623), .ZN(new_n694));
  OAI211_X1 g0494(.A(KEYINPUT29), .B(new_n642), .C1(new_n690), .C2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n685), .B1(new_n689), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n669), .B1(new_n696), .B2(G1), .ZN(G364));
  INV_X1    g0497(.A(new_n651), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n290), .A2(G20), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n206), .B1(new_n700), .B2(G45), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OR3_X1    g0502(.A1(new_n661), .A2(KEYINPUT95), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT95), .B1(new_n661), .B2(new_n702), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n699), .A2(new_n653), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT96), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n215), .B1(G20), .B2(new_n341), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(G179), .A2(G200), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n207), .B1(new_n711), .B2(G190), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n498), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n307), .A2(new_n403), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n207), .A2(G190), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n713), .B1(G68), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT98), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n403), .A2(G179), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n418), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n207), .A2(new_n279), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n714), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n722), .B1(G50), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G58), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n307), .A2(G200), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n715), .A2(new_n728), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT97), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n730), .A2(KEYINPUT97), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI221_X1 g0534(.A(new_n726), .B1(new_n727), .B2(new_n729), .C1(new_n734), .C2(new_n226), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n715), .A2(new_n711), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n736), .A2(KEYINPUT32), .A3(new_n377), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n723), .A2(new_n720), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G87), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT32), .B1(new_n736), .B2(new_n377), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(new_n258), .A3(new_n741), .ZN(new_n742));
  OR4_X1    g0542(.A1(new_n719), .A2(new_n735), .A3(new_n737), .A4(new_n742), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n736), .A2(KEYINPUT99), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n736), .A2(KEYINPUT99), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G329), .ZN(new_n748));
  INV_X1    g0548(.A(G294), .ZN(new_n749));
  INV_X1    g0549(.A(G303), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n383), .B1(new_n712), .B2(new_n749), .C1(new_n750), .C2(new_n738), .ZN(new_n751));
  XOR2_X1   g0551(.A(KEYINPUT33), .B(G317), .Z(new_n752));
  INV_X1    g0552(.A(G326), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n716), .A2(new_n752), .B1(new_n724), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G322), .ZN(new_n755));
  INV_X1    g0555(.A(G283), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n729), .A2(new_n755), .B1(new_n721), .B2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n751), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n748), .B(new_n758), .C1(new_n759), .C2(new_n734), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n710), .B1(new_n743), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n709), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n660), .A2(new_n383), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n766), .A2(G355), .B1(new_n558), .B2(new_n660), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n221), .A2(G45), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(new_n249), .B2(G45), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n660), .A2(new_n258), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n767), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n705), .B(new_n761), .C1(new_n765), .C2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n764), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n698), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n708), .A2(new_n775), .ZN(G396));
  NOR2_X1   g0576(.A1(new_n709), .A2(new_n762), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n705), .B1(new_n226), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n734), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n779), .A2(G116), .B1(new_n747), .B2(G311), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n721), .A2(new_n356), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n729), .A2(new_n749), .B1(new_n716), .B2(new_n756), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n781), .B(new_n782), .C1(G303), .C2(new_n725), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n258), .B(new_n713), .C1(G107), .C2(new_n739), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n780), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n383), .B1(new_n739), .B2(G50), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n786), .B1(new_n727), .B2(new_n712), .C1(new_n313), .C2(new_n721), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G132), .B2(new_n747), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G137), .A2(new_n725), .B1(new_n717), .B2(G150), .ZN(new_n789));
  INV_X1    g0589(.A(G143), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n789), .B1(new_n790), .B2(new_n729), .C1(new_n734), .C2(new_n377), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n788), .B1(new_n792), .B2(KEYINPUT34), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT34), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n785), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n796), .A2(KEYINPUT100), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n709), .B1(new_n796), .B2(KEYINPUT100), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n432), .A2(new_n641), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n435), .B2(new_n432), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n433), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n630), .A2(new_n642), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n778), .B1(new_n797), .B2(new_n798), .C1(new_n804), .C2(new_n763), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n686), .B(new_n803), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n706), .B1(new_n806), .B2(new_n685), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n806), .A2(new_n685), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n805), .B1(new_n808), .B2(new_n809), .ZN(G384));
  OAI211_X1 g0610(.A(G116), .B(new_n217), .C1(new_n506), .C2(KEYINPUT35), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(KEYINPUT35), .B2(new_n506), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT36), .ZN(new_n813));
  OR3_X1    g0613(.A1(new_n220), .A2(new_n226), .A3(new_n374), .ZN(new_n814));
  INV_X1    g0614(.A(G50), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G68), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n206), .B(G13), .C1(new_n814), .C2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n686), .A2(new_n804), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n802), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT38), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT103), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT102), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT16), .B1(new_n389), .B2(new_n393), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n281), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n386), .A2(KEYINPUT102), .A3(new_n316), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n826), .A3(new_n394), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n368), .B1(new_n827), .B2(new_n398), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n408), .A2(new_n395), .A3(new_n398), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n822), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n394), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n389), .A2(new_n393), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n281), .B1(new_n832), .B2(new_n370), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n833), .B2(KEYINPUT102), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n397), .B1(new_n834), .B2(new_n825), .ZN(new_n835));
  OAI211_X1 g0635(.A(KEYINPUT103), .B(new_n409), .C1(new_n835), .C2(new_n368), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n639), .B1(new_n827), .B2(new_n398), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n830), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT37), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT105), .ZN(new_n841));
  INV_X1    g0641(.A(new_n639), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n399), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n400), .A2(new_n409), .A3(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n840), .A2(new_n841), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n838), .B1(new_n402), .B2(new_n410), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n847), .B1(new_n839), .B2(KEYINPUT37), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(new_n841), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n821), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n827), .A2(new_n398), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n829), .B1(new_n857), .B2(new_n369), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n837), .B1(new_n858), .B2(KEYINPUT103), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n856), .B1(new_n859), .B2(new_n830), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT105), .B1(new_n860), .B2(new_n847), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n849), .A4(new_n851), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n324), .A2(new_n641), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n348), .A2(new_n415), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT101), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n348), .A2(KEYINPUT101), .A3(new_n415), .A4(new_n864), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n346), .A2(new_n347), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n324), .B(new_n641), .C1(new_n869), .C2(new_n416), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n820), .A2(new_n863), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n402), .B2(new_n842), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT106), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n863), .A2(new_n874), .A3(KEYINPUT39), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT39), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT107), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n844), .A2(new_n877), .A3(new_n846), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n877), .B1(new_n844), .B2(new_n846), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n878), .A2(new_n879), .A3(new_n847), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n843), .B1(new_n402), .B2(new_n410), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n821), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n862), .A2(new_n876), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n883), .A2(new_n874), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n876), .B1(new_n855), .B2(new_n862), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n875), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n349), .A2(new_n642), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n873), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n689), .A2(new_n438), .A3(new_n695), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n634), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n889), .B(new_n891), .Z(new_n892));
  NAND2_X1  g0692(.A1(new_n862), .A2(new_n882), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n680), .A2(KEYINPUT31), .A3(new_n641), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n681), .B2(KEYINPUT108), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT108), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n896), .B(KEYINPUT31), .C1(new_n680), .C2(new_n641), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n670), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n899), .A2(new_n804), .A3(KEYINPUT40), .A4(new_n871), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n804), .A3(new_n871), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n855), .B2(new_n862), .ZN(new_n904));
  OAI211_X1 g0704(.A(G330), .B(new_n902), .C1(new_n904), .C2(KEYINPUT40), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n438), .A2(G330), .A3(new_n899), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT109), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n905), .A2(KEYINPUT109), .A3(new_n906), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n900), .B1(new_n862), .B2(new_n882), .ZN(new_n911));
  INV_X1    g0711(.A(new_n903), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n850), .B1(new_n853), .B2(new_n841), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n913), .A2(KEYINPUT38), .A3(new_n861), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n913), .B2(new_n861), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n438), .A3(new_n899), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n909), .A2(new_n910), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n892), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n206), .B2(new_n700), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n892), .A2(new_n920), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n818), .B1(new_n922), .B2(new_n923), .ZN(G367));
  NOR2_X1   g0724(.A1(new_n771), .A2(new_n245), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n765), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n660), .B2(new_n427), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n705), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n712), .A2(new_n313), .ZN(new_n930));
  AOI22_X1  g0730(.A1(G58), .A2(new_n739), .B1(new_n717), .B2(G159), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n931), .B1(new_n790), .B2(new_n724), .C1(new_n734), .C2(new_n815), .ZN(new_n932));
  INV_X1    g0732(.A(G137), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n258), .B1(new_n736), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(G150), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n729), .A2(new_n935), .B1(new_n721), .B2(new_n226), .ZN(new_n936));
  OR4_X1    g0736(.A1(new_n930), .A2(new_n932), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n729), .A2(new_n750), .B1(new_n716), .B2(new_n749), .ZN(new_n938));
  INV_X1    g0738(.A(G317), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n504), .A2(new_n721), .B1(new_n736), .B2(new_n939), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n938), .B(new_n940), .C1(new_n779), .C2(G283), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n739), .A2(G116), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT46), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n258), .B(new_n944), .C1(G311), .C2(new_n725), .ZN(new_n945));
  INV_X1    g0745(.A(new_n712), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n942), .A2(new_n943), .B1(new_n946), .B2(G107), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT47), .B1(new_n937), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n937), .A2(KEYINPUT47), .A3(new_n948), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n709), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n461), .A2(new_n475), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n641), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n489), .B2(new_n491), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n691), .B2(new_n953), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n929), .B1(new_n949), .B2(new_n951), .C1(new_n955), .C2(new_n774), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n646), .B(new_n653), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(new_n655), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n540), .A2(new_n542), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n510), .B2(new_n657), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n692), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n532), .A2(new_n657), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n656), .B2(new_n658), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT44), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT110), .ZN(new_n968));
  INV_X1    g0768(.A(new_n654), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n965), .A2(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n656), .A2(new_n658), .A3(new_n964), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT45), .Z(new_n973));
  NAND2_X1  g0773(.A1(new_n654), .A2(KEYINPUT110), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n974), .B1(new_n971), .B2(new_n973), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n696), .B(new_n958), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n696), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n661), .B(KEYINPUT41), .Z(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n702), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n658), .B1(new_n656), .B2(KEYINPUT42), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n964), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n646), .A2(new_n655), .A3(new_n961), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n984), .A2(KEYINPUT42), .B1(new_n532), .B2(new_n657), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n983), .A2(new_n985), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n986));
  OR3_X1    g0786(.A1(new_n986), .A2(KEYINPUT43), .A3(new_n955), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n986), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n969), .A2(new_n964), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n988), .A2(new_n969), .A3(new_n964), .A4(new_n987), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n956), .B1(new_n981), .B2(new_n993), .ZN(G387));
  NAND2_X1  g0794(.A1(new_n958), .A2(new_n702), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n766), .A2(new_n663), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(G107), .B2(new_n210), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n242), .A2(G45), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT111), .Z(new_n999));
  AOI211_X1 g0799(.A(G45), .B(new_n663), .C1(G68), .C2(G77), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n283), .A2(G50), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n771), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n997), .B1(new_n999), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n706), .B1(new_n1004), .B2(new_n927), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT112), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n721), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n258), .B1(new_n1007), .B2(G116), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n734), .A2(new_n750), .B1(new_n939), .B2(new_n729), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT114), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(KEYINPUT114), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G322), .A2(new_n725), .B1(new_n717), .B2(G311), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT48), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n739), .A2(G294), .B1(new_n946), .B2(G283), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT49), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1008), .B1(new_n753), .B2(new_n736), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n1019), .B2(new_n1018), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n734), .A2(new_n313), .B1(new_n283), .B2(new_n716), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT113), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G77), .A2(new_n739), .B1(new_n1007), .B2(G97), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n815), .B2(new_n729), .C1(new_n935), .C2(new_n736), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n712), .A2(new_n426), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n258), .B1(new_n724), .B2(new_n377), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n709), .B1(new_n1021), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1006), .A2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT115), .Z(new_n1031));
  NOR2_X1   g0831(.A1(new_n646), .A2(new_n774), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n958), .A2(new_n696), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n661), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n958), .A2(new_n696), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n995), .B1(new_n1031), .B2(new_n1032), .C1(new_n1034), .C2(new_n1035), .ZN(G393));
  NAND2_X1  g0836(.A1(new_n971), .A2(new_n973), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n974), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n1033), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n977), .A2(new_n661), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n779), .A2(G294), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n724), .A2(new_n939), .B1(new_n729), .B2(new_n759), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT52), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n716), .A2(new_n750), .B1(new_n736), .B2(new_n755), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G283), .B2(new_n739), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n258), .B(new_n722), .C1(G116), .C2(new_n946), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n779), .A2(new_n284), .B1(G50), .B2(new_n717), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(KEYINPUT116), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n724), .A2(new_n935), .B1(new_n729), .B2(new_n377), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT51), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n738), .A2(new_n313), .B1(new_n736), .B2(new_n790), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n712), .A2(new_n226), .ZN(new_n1055));
  NOR4_X1   g0855(.A1(new_n1054), .A2(new_n781), .A3(new_n1055), .A4(new_n383), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1051), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1050), .A2(KEYINPUT116), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1049), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n709), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n771), .A2(new_n252), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n765), .B1(new_n210), .B2(new_n504), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1060), .B(new_n706), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n963), .B2(new_n764), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n702), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1042), .A2(new_n1066), .ZN(G390));
  INV_X1    g0867(.A(new_n802), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n686), .B2(new_n804), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n871), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n887), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n875), .B(new_n1071), .C1(new_n884), .C2(new_n885), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n642), .B(new_n801), .C1(new_n690), .C2(new_n694), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n802), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n871), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n893), .A3(new_n887), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n685), .A2(new_n804), .A3(new_n871), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n1072), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n899), .A2(G330), .A3(new_n804), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n871), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n702), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n777), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n706), .B1(new_n284), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n740), .A2(new_n383), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n724), .A2(new_n756), .B1(new_n716), .B2(new_n418), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n729), .A2(new_n558), .B1(new_n721), .B2(new_n313), .ZN(new_n1089));
  NOR4_X1   g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .A4(new_n1055), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n749), .B2(new_n746), .C1(new_n504), .C2(new_n734), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n258), .B1(new_n716), .B2(new_n933), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G159), .B2(new_n946), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n725), .A2(G128), .B1(new_n1007), .B2(G50), .ZN(new_n1094));
  INV_X1    g0894(.A(G132), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1094), .C1(new_n1095), .C2(new_n729), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n738), .A2(new_n935), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT53), .ZN(new_n1098));
  INV_X1    g0898(.A(G125), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT54), .B(G143), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n746), .C1(new_n734), .C2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1091), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1086), .B1(new_n1102), .B2(new_n709), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n886), .B2(new_n763), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1084), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n661), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n890), .A2(new_n906), .A3(new_n634), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n685), .A2(new_n804), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1070), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(KEYINPUT117), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1081), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1109), .A2(KEYINPUT117), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n820), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1074), .B1(new_n1070), .B2(new_n1079), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1077), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1107), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1083), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1106), .B1(new_n1117), .B2(KEYINPUT118), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1082), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1072), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n1120), .A3(new_n1116), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT118), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1116), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1105), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(G378));
  INV_X1    g0927(.A(KEYINPUT121), .ZN(new_n1128));
  XOR2_X1   g0928(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1129));
  NOR2_X1   g0929(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT73), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1130), .B1(new_n1133), .B2(new_n303), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n297), .A2(new_n639), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1134), .A2(new_n310), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1135), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n306), .B2(new_n311), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1129), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1135), .B1(new_n1134), .B2(new_n310), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n306), .A2(new_n311), .A3(new_n1137), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1129), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1128), .B1(new_n905), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n918), .A2(KEYINPUT121), .A3(G330), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n905), .A2(new_n1144), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1148), .A2(new_n889), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n889), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1107), .B1(new_n1083), .B2(new_n1116), .ZN(new_n1153));
  OAI21_X1  g0953(.A(KEYINPUT57), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n889), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1148), .A2(new_n889), .A3(new_n1149), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1107), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1121), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1154), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n661), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1144), .A2(new_n762), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n706), .B1(G50), .B2(new_n1085), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(G33), .A2(G41), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT119), .ZN(new_n1169));
  AOI211_X1 g0969(.A(G50), .B(new_n1169), .C1(new_n266), .C2(new_n383), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n729), .A2(new_n418), .B1(new_n721), .B2(new_n727), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n724), .A2(new_n558), .B1(new_n738), .B2(new_n226), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n266), .B(new_n383), .C1(new_n716), .C2(new_n498), .ZN(new_n1173));
  NOR4_X1   g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n930), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n756), .B2(new_n746), .C1(new_n426), .C2(new_n734), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT58), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1170), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(G128), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n724), .A2(new_n1099), .B1(new_n729), .B2(new_n1178), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1095), .A2(new_n716), .B1(new_n738), .B2(new_n1100), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(G150), .C2(new_n946), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n933), .B2(new_n734), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  INV_X1    g0983(.A(G124), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1169), .B1(new_n1184), .B2(new_n736), .C1(new_n377), .C2(new_n721), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT120), .Z(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1177), .B1(new_n1176), .B2(new_n1175), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1167), .B1(new_n1189), .B2(new_n709), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1159), .A2(new_n702), .B1(new_n1166), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1165), .A2(new_n1191), .ZN(G375));
  NAND2_X1  g0992(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n871), .A2(new_n763), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G294), .A2(new_n725), .B1(new_n739), .B2(G97), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n558), .B2(new_n716), .C1(new_n756), .C2(new_n729), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n734), .A2(new_n418), .B1(new_n746), .B2(new_n750), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n383), .B1(new_n721), .B2(new_n226), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1026), .A4(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT122), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(KEYINPUT122), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n258), .B1(new_n712), .B2(new_n815), .C1(new_n727), .C2(new_n721), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n724), .A2(new_n1095), .B1(new_n729), .B2(new_n933), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n377), .A2(new_n738), .B1(new_n716), .B2(new_n1100), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n1178), .B2(new_n746), .C1(new_n935), .C2(new_n734), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1201), .A2(new_n1202), .A3(new_n1207), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n706), .B1(G68), .B2(new_n1085), .C1(new_n1208), .C2(new_n710), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n1194), .A2(new_n701), .B1(new_n1195), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1194), .A2(new_n1107), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1212), .A2(new_n980), .A3(new_n1123), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1213), .ZN(G381));
  OR4_X1    g1014(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1165), .A2(new_n1126), .A3(new_n1191), .ZN(new_n1216));
  OR4_X1    g1016(.A1(G387), .A2(new_n1215), .A3(new_n1216), .A4(G381), .ZN(G407));
  OAI211_X1 g1017(.A(G407), .B(G213), .C1(G343), .C2(new_n1216), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT123), .ZN(G409));
  INV_X1    g1019(.A(G390), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1033), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n696), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n980), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n993), .B1(new_n1223), .B2(new_n701), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n956), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1220), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT126), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n956), .B(G390), .C1(new_n981), .C2(new_n993), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  XOR2_X1   g1029(.A(G393), .B(G396), .Z(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1230), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1226), .B(new_n1228), .C1(new_n1232), .C2(KEYINPUT126), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT61), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1123), .A2(new_n661), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1212), .A2(KEYINPUT60), .ZN(new_n1237));
  OR3_X1    g1037(.A1(new_n1193), .A2(KEYINPUT60), .A3(new_n1161), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(G384), .ZN(new_n1240));
  OR3_X1    g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n1210), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT125), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1239), .B2(new_n1210), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(G213), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(G343), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1246), .A2(G2897), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1243), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1239), .A2(new_n1240), .A3(new_n1210), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1248), .B1(new_n1242), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1251), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(KEYINPUT125), .A3(new_n1247), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1165), .A2(G378), .A3(new_n1191), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1159), .A2(new_n980), .A3(new_n1162), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1191), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1126), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1246), .B1(new_n1256), .B2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1234), .B(new_n1235), .C1(new_n1255), .C2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT124), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(new_n1263), .A3(new_n1251), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1246), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1106), .B1(new_n1154), .B2(new_n1163), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1191), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1266), .A2(new_n1126), .A3(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1259), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1265), .B(new_n1251), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT124), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1264), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1251), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1262), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1235), .B1(new_n1255), .B2(new_n1260), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT127), .B1(new_n1270), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT127), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1260), .A2(new_n1279), .A3(KEYINPUT62), .A4(new_n1251), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1264), .A2(new_n1271), .A3(new_n1277), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1276), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1275), .B1(new_n1283), .B2(new_n1234), .ZN(G405));
  NAND2_X1  g1084(.A1(new_n1234), .A2(new_n1253), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1231), .A2(new_n1251), .A3(new_n1233), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G375), .B(new_n1126), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1287), .B(new_n1288), .ZN(G402));
endmodule


