

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744;

  NOR2_X1 U372 ( .A1(n566), .A2(n567), .ZN(n732) );
  AND2_X1 U373 ( .A1(n586), .A2(n367), .ZN(n351) );
  OR2_X1 U374 ( .A1(n675), .A2(n393), .ZN(n389) );
  OR2_X1 U375 ( .A1(n478), .A2(n477), .ZN(n480) );
  XNOR2_X1 U376 ( .A(n406), .B(G107), .ZN(n511) );
  NAND2_X1 U377 ( .A1(n560), .A2(n561), .ZN(n670) );
  AND2_X1 U378 ( .A1(n592), .A2(n590), .ZN(n350) );
  XNOR2_X2 U379 ( .A(n461), .B(n353), .ZN(n579) );
  INV_X1 U380 ( .A(G116), .ZN(n406) );
  XNOR2_X1 U381 ( .A(n471), .B(n470), .ZN(n724) );
  NOR2_X1 U382 ( .A1(n709), .A2(n717), .ZN(n362) );
  XNOR2_X1 U383 ( .A(n386), .B(n359), .ZN(n709) );
  NOR2_X1 U384 ( .A1(n382), .A2(n601), .ZN(n381) );
  AND2_X1 U385 ( .A1(n589), .A2(KEYINPUT44), .ZN(n601) );
  XNOR2_X1 U386 ( .A(n583), .B(KEYINPUT22), .ZN(n595) );
  NOR2_X1 U387 ( .A1(n549), .A2(n543), .ZN(n546) );
  XNOR2_X1 U388 ( .A(n699), .B(n413), .ZN(n702) );
  OR2_X1 U389 ( .A1(n699), .A2(G902), .ZN(n397) );
  XNOR2_X1 U390 ( .A(n730), .B(G146), .ZN(n441) );
  XNOR2_X1 U391 ( .A(n482), .B(n370), .ZN(n730) );
  XNOR2_X1 U392 ( .A(n416), .B(G137), .ZN(n370) );
  INV_X2 U393 ( .A(G143), .ZN(n414) );
  INV_X1 U394 ( .A(n472), .ZN(n733) );
  NOR2_X2 U395 ( .A1(n595), .A2(n593), .ZN(n586) );
  NOR2_X2 U396 ( .A1(n626), .A2(n742), .ZN(n592) );
  XNOR2_X2 U397 ( .A(n351), .B(KEYINPUT32), .ZN(n742) );
  AND2_X1 U398 ( .A1(n650), .A2(n649), .ZN(n574) );
  XNOR2_X1 U399 ( .A(n740), .B(n578), .ZN(n591) );
  NOR2_X1 U400 ( .A1(n563), .A2(n632), .ZN(n565) );
  NAND2_X1 U401 ( .A1(n364), .A2(n363), .ZN(n563) );
  XNOR2_X1 U402 ( .A(n511), .B(n405), .ZN(n469) );
  INV_X1 U403 ( .A(KEYINPUT73), .ZN(n405) );
  NAND2_X1 U404 ( .A1(n369), .A2(n633), .ZN(n542) );
  XNOR2_X1 U405 ( .A(n524), .B(KEYINPUT104), .ZN(n369) );
  INV_X1 U406 ( .A(KEYINPUT1), .ZN(n395) );
  NOR2_X1 U407 ( .A1(G953), .A2(G237), .ZN(n498) );
  NOR2_X1 U408 ( .A1(n642), .A2(n357), .ZN(n363) );
  AND2_X1 U409 ( .A1(n515), .A2(G221), .ZN(n368) );
  XNOR2_X1 U410 ( .A(G119), .B(G110), .ZN(n448) );
  XOR2_X1 U411 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n449) );
  XOR2_X1 U412 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n508) );
  XNOR2_X1 U413 ( .A(G134), .B(G122), .ZN(n507) );
  XOR2_X1 U414 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n506) );
  XNOR2_X1 U415 ( .A(n398), .B(n445), .ZN(n729) );
  XOR2_X1 U416 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n445) );
  XNOR2_X1 U417 ( .A(n481), .B(G140), .ZN(n398) );
  AND2_X1 U418 ( .A1(n350), .A2(n591), .ZN(n382) );
  AND2_X1 U419 ( .A1(n593), .A2(n352), .ZN(n650) );
  NAND2_X1 U420 ( .A1(n650), .A2(n535), .ZN(n375) );
  XNOR2_X1 U421 ( .A(n464), .B(n373), .ZN(n372) );
  XNOR2_X1 U422 ( .A(n463), .B(n465), .ZN(n373) );
  NOR2_X1 U423 ( .A1(n462), .A2(n579), .ZN(n464) );
  XNOR2_X1 U424 ( .A(n441), .B(n425), .ZN(n460) );
  NAND2_X1 U425 ( .A1(n404), .A2(n402), .ZN(n407) );
  INV_X1 U426 ( .A(KEYINPUT4), .ZN(n415) );
  XNOR2_X1 U427 ( .A(n399), .B(G125), .ZN(n481) );
  INV_X1 U428 ( .A(G146), .ZN(n399) );
  XNOR2_X1 U429 ( .A(n489), .B(KEYINPUT39), .ZN(n530) );
  NAND2_X1 U430 ( .A1(n385), .A2(n667), .ZN(n549) );
  INV_X1 U431 ( .A(KEYINPUT108), .ZN(n544) );
  INV_X1 U432 ( .A(n576), .ZN(n391) );
  XNOR2_X1 U433 ( .A(n579), .B(n521), .ZN(n585) );
  XNOR2_X1 U434 ( .A(n504), .B(n503), .ZN(n560) );
  INV_X1 U435 ( .A(G469), .ZN(n396) );
  AND2_X1 U436 ( .A1(n580), .A2(n352), .ZN(n581) );
  XNOR2_X1 U437 ( .A(KEYINPUT16), .B(KEYINPUT72), .ZN(n468) );
  INV_X1 U438 ( .A(n593), .ZN(n654) );
  XNOR2_X1 U439 ( .A(G113), .B(G116), .ZN(n421) );
  INV_X1 U440 ( .A(KEYINPUT5), .ZN(n420) );
  XOR2_X1 U441 ( .A(KEYINPUT90), .B(KEYINPUT74), .Z(n419) );
  NAND2_X1 U442 ( .A1(n401), .A2(n409), .ZN(n400) );
  XNOR2_X1 U443 ( .A(n493), .B(n492), .ZN(n494) );
  NAND2_X1 U444 ( .A1(G234), .A2(G237), .ZN(n428) );
  OR2_X1 U445 ( .A1(G237), .A2(G902), .ZN(n486) );
  XNOR2_X1 U446 ( .A(G902), .B(KEYINPUT15), .ZN(n615) );
  INV_X1 U447 ( .A(n615), .ZN(n408) );
  XNOR2_X1 U448 ( .A(n417), .B(n383), .ZN(n467) );
  XNOR2_X1 U449 ( .A(n384), .B(G119), .ZN(n383) );
  INV_X1 U450 ( .A(G101), .ZN(n384) );
  INV_X1 U451 ( .A(G953), .ZN(n719) );
  XNOR2_X1 U452 ( .A(n454), .B(n453), .ZN(n716) );
  XNOR2_X1 U453 ( .A(n368), .B(n729), .ZN(n454) );
  XNOR2_X1 U454 ( .A(G137), .B(G128), .ZN(n451) );
  XOR2_X1 U455 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n447) );
  XNOR2_X1 U456 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n505) );
  XOR2_X1 U457 ( .A(G140), .B(G107), .Z(n437) );
  XNOR2_X1 U458 ( .A(G101), .B(G104), .ZN(n436) );
  AND2_X2 U459 ( .A1(n407), .A2(n408), .ZN(n715) );
  AND2_X1 U460 ( .A1(n613), .A2(n600), .ZN(n380) );
  AND2_X1 U461 ( .A1(n372), .A2(n371), .ZN(n366) );
  XNOR2_X1 U462 ( .A(n375), .B(KEYINPUT105), .ZN(n374) );
  INV_X1 U463 ( .A(n522), .ZN(n371) );
  XNOR2_X1 U464 ( .A(n549), .B(KEYINPUT19), .ZN(n572) );
  NAND2_X1 U465 ( .A1(n715), .A2(G217), .ZN(n379) );
  NAND2_X1 U466 ( .A1(n715), .A2(G475), .ZN(n386) );
  XNOR2_X1 U467 ( .A(n485), .B(n724), .ZN(n694) );
  XNOR2_X1 U468 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U469 ( .A1(n480), .A2(n479), .ZN(n484) );
  NOR2_X1 U470 ( .A1(n733), .A2(G952), .ZN(n717) );
  INV_X1 U471 ( .A(KEYINPUT40), .ZN(n531) );
  XNOR2_X1 U472 ( .A(n544), .B(KEYINPUT36), .ZN(n545) );
  NOR2_X1 U473 ( .A1(n392), .A2(n391), .ZN(n390) );
  AND2_X1 U474 ( .A1(n587), .A2(n649), .ZN(n367) );
  XNOR2_X1 U475 ( .A(n376), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U476 ( .A1(n378), .A2(n377), .ZN(n376) );
  INV_X1 U477 ( .A(n717), .ZN(n377) );
  XNOR2_X1 U478 ( .A(n379), .B(n360), .ZN(n378) );
  XOR2_X1 U479 ( .A(n653), .B(KEYINPUT88), .Z(n352) );
  XOR2_X1 U480 ( .A(G472), .B(KEYINPUT71), .Z(n353) );
  XNOR2_X1 U481 ( .A(n487), .B(n488), .ZN(n354) );
  INV_X1 U482 ( .A(n365), .ZN(n559) );
  NAND2_X1 U483 ( .A1(n374), .A2(n366), .ZN(n365) );
  NOR2_X1 U484 ( .A1(n566), .A2(n400), .ZN(n355) );
  AND2_X1 U485 ( .A1(n732), .A2(n718), .ZN(n356) );
  AND2_X1 U486 ( .A1(n558), .A2(n557), .ZN(n357) );
  XNOR2_X1 U487 ( .A(KEYINPUT80), .B(KEYINPUT45), .ZN(n358) );
  XOR2_X1 U488 ( .A(n708), .B(n707), .Z(n359) );
  XOR2_X1 U489 ( .A(n716), .B(KEYINPUT124), .Z(n360) );
  AND2_X1 U490 ( .A1(n408), .A2(G472), .ZN(n361) );
  INV_X1 U491 ( .A(KEYINPUT2), .ZN(n409) );
  NOR2_X1 U492 ( .A1(n704), .A2(n717), .ZN(n705) );
  NOR2_X1 U493 ( .A1(n697), .A2(n717), .ZN(n698) );
  XNOR2_X1 U494 ( .A(n362), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U495 ( .A1(n694), .A2(n615), .ZN(n410) );
  XNOR2_X1 U496 ( .A(n703), .B(n702), .ZN(n704) );
  AND2_X2 U497 ( .A1(n387), .A2(n390), .ZN(n577) );
  INV_X1 U498 ( .A(n548), .ZN(n364) );
  NAND2_X1 U499 ( .A1(n718), .A2(n732), .ZN(n403) );
  XNOR2_X2 U500 ( .A(n614), .B(n358), .ZN(n718) );
  XNOR2_X1 U501 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U502 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X2 U503 ( .A(n512), .B(n415), .ZN(n482) );
  NAND2_X1 U504 ( .A1(n381), .A2(n380), .ZN(n614) );
  INV_X1 U505 ( .A(n385), .ZN(n527) );
  XNOR2_X2 U506 ( .A(n410), .B(n354), .ZN(n385) );
  XNOR2_X1 U507 ( .A(n527), .B(KEYINPUT38), .ZN(n666) );
  NAND2_X1 U508 ( .A1(n576), .A2(n385), .ZN(n562) );
  NAND2_X1 U509 ( .A1(n403), .A2(KEYINPUT2), .ZN(n402) );
  XNOR2_X2 U510 ( .A(n573), .B(KEYINPUT0), .ZN(n602) );
  NAND2_X1 U511 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U512 ( .A1(n675), .A2(n394), .ZN(n388) );
  XNOR2_X2 U513 ( .A(n411), .B(KEYINPUT33), .ZN(n675) );
  AND2_X1 U514 ( .A1(n602), .A2(n575), .ZN(n392) );
  NOR2_X1 U515 ( .A1(n602), .A2(n575), .ZN(n393) );
  INV_X1 U516 ( .A(n575), .ZN(n394) );
  XNOR2_X2 U517 ( .A(n607), .B(n395), .ZN(n649) );
  XNOR2_X2 U518 ( .A(n397), .B(n396), .ZN(n607) );
  XNOR2_X2 U519 ( .A(n455), .B(n456), .ZN(n593) );
  INV_X1 U520 ( .A(n567), .ZN(n401) );
  NAND2_X1 U521 ( .A1(n355), .A2(n718), .ZN(n404) );
  NAND2_X1 U522 ( .A1(n407), .A2(n361), .ZN(n616) );
  AND2_X1 U523 ( .A1(n596), .A2(n574), .ZN(n411) );
  XNOR2_X1 U524 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n412) );
  XOR2_X1 U525 ( .A(n701), .B(n700), .Z(n413) );
  INV_X1 U526 ( .A(KEYINPUT94), .ZN(n492) );
  XNOR2_X1 U527 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U528 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U529 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U530 ( .A(n439), .B(n438), .ZN(n440) );
  INV_X1 U531 ( .A(KEYINPUT48), .ZN(n564) );
  XNOR2_X1 U532 ( .A(n502), .B(G475), .ZN(n503) );
  INV_X1 U533 ( .A(n572), .ZN(n550) );
  NOR2_X1 U534 ( .A1(n717), .A2(n618), .ZN(n619) );
  XNOR2_X1 U535 ( .A(n532), .B(n531), .ZN(n743) );
  XNOR2_X2 U536 ( .A(G953), .B(KEYINPUT64), .ZN(n472) );
  XOR2_X1 U537 ( .A(KEYINPUT82), .B(KEYINPUT62), .Z(n427) );
  XNOR2_X2 U538 ( .A(n414), .B(G128), .ZN(n512) );
  XOR2_X1 U539 ( .A(G131), .B(G134), .Z(n416) );
  XNOR2_X1 U540 ( .A(KEYINPUT68), .B(KEYINPUT3), .ZN(n417) );
  NAND2_X1 U541 ( .A1(n498), .A2(G210), .ZN(n418) );
  XNOR2_X1 U542 ( .A(n419), .B(n418), .ZN(n423) );
  XNOR2_X1 U543 ( .A(n467), .B(n424), .ZN(n425) );
  XOR2_X1 U544 ( .A(n460), .B(KEYINPUT109), .Z(n426) );
  XNOR2_X1 U545 ( .A(n427), .B(n426), .ZN(n617) );
  XNOR2_X1 U546 ( .A(n428), .B(KEYINPUT14), .ZN(n429) );
  AND2_X1 U547 ( .A1(G952), .A2(n429), .ZN(n682) );
  NAND2_X1 U548 ( .A1(n682), .A2(n719), .ZN(n569) );
  INV_X1 U549 ( .A(n569), .ZN(n433) );
  NAND2_X1 U550 ( .A1(n429), .A2(G902), .ZN(n430) );
  XNOR2_X1 U551 ( .A(n430), .B(KEYINPUT85), .ZN(n568) );
  NAND2_X1 U552 ( .A1(n472), .A2(n568), .ZN(n431) );
  NOR2_X1 U553 ( .A1(G900), .A2(n431), .ZN(n432) );
  NOR2_X1 U554 ( .A1(n433), .A2(n432), .ZN(n522) );
  XOR2_X1 U555 ( .A(KEYINPUT69), .B(G110), .Z(n476) );
  XOR2_X1 U556 ( .A(n476), .B(KEYINPUT76), .Z(n435) );
  NAND2_X1 U557 ( .A1(G227), .A2(n733), .ZN(n434) );
  XNOR2_X1 U558 ( .A(n435), .B(n434), .ZN(n439) );
  XNOR2_X1 U559 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U560 ( .A(n441), .B(n440), .ZN(n699) );
  INV_X1 U561 ( .A(n607), .ZN(n535) );
  XOR2_X1 U562 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n444) );
  NAND2_X1 U563 ( .A1(G234), .A2(n615), .ZN(n442) );
  XNOR2_X1 U564 ( .A(KEYINPUT20), .B(n442), .ZN(n457) );
  NAND2_X1 U565 ( .A1(n457), .A2(G217), .ZN(n443) );
  XNOR2_X1 U566 ( .A(n444), .B(n443), .ZN(n456) );
  NAND2_X1 U567 ( .A1(G234), .A2(n733), .ZN(n446) );
  XNOR2_X1 U568 ( .A(n447), .B(n446), .ZN(n515) );
  XNOR2_X1 U569 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U570 ( .A(n450), .B(KEYINPUT23), .Z(n452) );
  XNOR2_X1 U571 ( .A(n452), .B(n451), .ZN(n453) );
  NOR2_X1 U572 ( .A1(n716), .A2(G902), .ZN(n455) );
  XOR2_X1 U573 ( .A(KEYINPUT87), .B(KEYINPUT21), .Z(n459) );
  NAND2_X1 U574 ( .A1(n457), .A2(G221), .ZN(n458) );
  XNOR2_X1 U575 ( .A(n459), .B(n458), .ZN(n653) );
  NAND2_X1 U576 ( .A1(G214), .A2(n486), .ZN(n667) );
  INV_X1 U577 ( .A(n667), .ZN(n462) );
  NOR2_X1 U578 ( .A1(G902), .A2(n460), .ZN(n461) );
  INV_X1 U579 ( .A(KEYINPUT106), .ZN(n463) );
  INV_X1 U580 ( .A(KEYINPUT30), .ZN(n465) );
  INV_X1 U581 ( .A(KEYINPUT84), .ZN(n488) );
  XNOR2_X1 U582 ( .A(G113), .B(G104), .ZN(n466) );
  XNOR2_X1 U583 ( .A(n466), .B(G122), .ZN(n497) );
  XNOR2_X1 U584 ( .A(n467), .B(n497), .ZN(n471) );
  XNOR2_X1 U585 ( .A(n469), .B(n468), .ZN(n470) );
  INV_X1 U586 ( .A(n472), .ZN(n473) );
  NAND2_X1 U587 ( .A1(n473), .A2(G224), .ZN(n475) );
  XOR2_X1 U588 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n474) );
  XNOR2_X1 U589 ( .A(n475), .B(n474), .ZN(n478) );
  INV_X1 U590 ( .A(n476), .ZN(n477) );
  NAND2_X1 U591 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U592 ( .A(n482), .B(n481), .ZN(n483) );
  NAND2_X1 U593 ( .A1(G210), .A2(n486), .ZN(n487) );
  NAND2_X1 U594 ( .A1(n559), .A2(n666), .ZN(n489) );
  XOR2_X1 U595 ( .A(KEYINPUT12), .B(KEYINPUT95), .Z(n491) );
  XNOR2_X1 U596 ( .A(G143), .B(KEYINPUT11), .ZN(n490) );
  XNOR2_X1 U597 ( .A(n491), .B(n490), .ZN(n495) );
  XNOR2_X1 U598 ( .A(G131), .B(KEYINPUT96), .ZN(n493) );
  XOR2_X1 U599 ( .A(n497), .B(n496), .Z(n501) );
  NAND2_X1 U600 ( .A1(G214), .A2(n498), .ZN(n499) );
  XNOR2_X1 U601 ( .A(n729), .B(n499), .ZN(n500) );
  XNOR2_X1 U602 ( .A(n501), .B(n500), .ZN(n706) );
  NOR2_X1 U603 ( .A1(G902), .A2(n706), .ZN(n504) );
  XNOR2_X1 U604 ( .A(KEYINPUT13), .B(KEYINPUT97), .ZN(n502) );
  XNOR2_X1 U605 ( .A(n506), .B(n505), .ZN(n510) );
  XNOR2_X1 U606 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U607 ( .A(n510), .B(n509), .Z(n514) );
  XNOR2_X1 U608 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U609 ( .A(n514), .B(n513), .ZN(n517) );
  NAND2_X1 U610 ( .A1(n515), .A2(G217), .ZN(n516) );
  XOR2_X1 U611 ( .A(n517), .B(n516), .Z(n712) );
  NOR2_X1 U612 ( .A1(G902), .A2(n712), .ZN(n519) );
  XNOR2_X1 U613 ( .A(KEYINPUT102), .B(G478), .ZN(n518) );
  XOR2_X1 U614 ( .A(n519), .B(n518), .Z(n537) );
  AND2_X1 U615 ( .A1(n560), .A2(n537), .ZN(n520) );
  XOR2_X1 U616 ( .A(KEYINPUT103), .B(n520), .Z(n628) );
  AND2_X1 U617 ( .A1(n530), .A2(n628), .ZN(n644) );
  INV_X1 U618 ( .A(n644), .ZN(n529) );
  NOR2_X1 U619 ( .A1(n560), .A2(n537), .ZN(n633) );
  INV_X1 U620 ( .A(n633), .ZN(n637) );
  INV_X1 U621 ( .A(KEYINPUT6), .ZN(n521) );
  NOR2_X1 U622 ( .A1(n522), .A2(n653), .ZN(n523) );
  NAND2_X1 U623 ( .A1(n654), .A2(n523), .ZN(n533) );
  NOR2_X1 U624 ( .A1(n585), .A2(n533), .ZN(n524) );
  NOR2_X1 U625 ( .A1(n649), .A2(n542), .ZN(n525) );
  NAND2_X1 U626 ( .A1(n525), .A2(n667), .ZN(n526) );
  XNOR2_X1 U627 ( .A(KEYINPUT43), .B(n526), .ZN(n528) );
  NAND2_X1 U628 ( .A1(n528), .A2(n527), .ZN(n645) );
  NAND2_X1 U629 ( .A1(n529), .A2(n645), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n530), .A2(n633), .ZN(n532) );
  NOR2_X1 U631 ( .A1(n533), .A2(n579), .ZN(n534) );
  XNOR2_X1 U632 ( .A(KEYINPUT28), .B(n534), .ZN(n536) );
  NAND2_X1 U633 ( .A1(n536), .A2(n535), .ZN(n551) );
  NAND2_X1 U634 ( .A1(n667), .A2(n666), .ZN(n671) );
  INV_X1 U635 ( .A(n537), .ZN(n561) );
  NOR2_X1 U636 ( .A1(n671), .A2(n670), .ZN(n538) );
  XNOR2_X1 U637 ( .A(n538), .B(KEYINPUT41), .ZN(n664) );
  NOR2_X1 U638 ( .A1(n551), .A2(n664), .ZN(n539) );
  XNOR2_X1 U639 ( .A(KEYINPUT42), .B(n539), .ZN(n744) );
  NOR2_X1 U640 ( .A1(n743), .A2(n744), .ZN(n541) );
  INV_X1 U641 ( .A(KEYINPUT46), .ZN(n540) );
  XNOR2_X1 U642 ( .A(n541), .B(n540), .ZN(n548) );
  INV_X1 U643 ( .A(n649), .ZN(n594) );
  XOR2_X1 U644 ( .A(KEYINPUT107), .B(n542), .Z(n543) );
  XNOR2_X1 U645 ( .A(n546), .B(n545), .ZN(n547) );
  NOR2_X1 U646 ( .A1(n594), .A2(n547), .ZN(n642) );
  NOR2_X1 U647 ( .A1(n633), .A2(n628), .ZN(n672) );
  NAND2_X1 U648 ( .A1(n672), .A2(KEYINPUT78), .ZN(n552) );
  NOR2_X1 U649 ( .A1(n551), .A2(n550), .ZN(n634) );
  NAND2_X1 U650 ( .A1(n552), .A2(n634), .ZN(n553) );
  INV_X1 U651 ( .A(KEYINPUT47), .ZN(n554) );
  NAND2_X1 U652 ( .A1(n553), .A2(n554), .ZN(n558) );
  AND2_X1 U653 ( .A1(n554), .A2(KEYINPUT78), .ZN(n555) );
  NOR2_X1 U654 ( .A1(n672), .A2(n555), .ZN(n556) );
  NAND2_X1 U655 ( .A1(n556), .A2(n634), .ZN(n557) );
  NOR2_X1 U656 ( .A1(n561), .A2(n560), .ZN(n576) );
  NOR2_X1 U657 ( .A1(n365), .A2(n562), .ZN(n632) );
  NOR2_X1 U658 ( .A1(G898), .A2(n719), .ZN(n726) );
  NAND2_X1 U659 ( .A1(n726), .A2(n568), .ZN(n570) );
  NAND2_X1 U660 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U661 ( .A1(n572), .A2(n571), .ZN(n573) );
  INV_X1 U662 ( .A(n585), .ZN(n596) );
  XNOR2_X1 U663 ( .A(KEYINPUT70), .B(KEYINPUT34), .ZN(n575) );
  XNOR2_X2 U664 ( .A(n577), .B(KEYINPUT35), .ZN(n740) );
  INV_X1 U665 ( .A(KEYINPUT65), .ZN(n578) );
  AND2_X1 U666 ( .A1(n740), .A2(n578), .ZN(n588) );
  INV_X1 U667 ( .A(n579), .ZN(n659) );
  INV_X1 U668 ( .A(n602), .ZN(n582) );
  INV_X1 U669 ( .A(n670), .ZN(n580) );
  NAND2_X1 U670 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U671 ( .A1(n594), .A2(n586), .ZN(n584) );
  NOR2_X1 U672 ( .A1(n659), .A2(n584), .ZN(n626) );
  XOR2_X1 U673 ( .A(n585), .B(KEYINPUT77), .Z(n587) );
  NAND2_X1 U674 ( .A1(n588), .A2(n592), .ZN(n589) );
  INV_X1 U675 ( .A(KEYINPUT44), .ZN(n590) );
  NAND2_X1 U676 ( .A1(n594), .A2(n593), .ZN(n599) );
  NOR2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U678 ( .A(n597), .B(KEYINPUT81), .ZN(n598) );
  NOR2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n620) );
  INV_X1 U680 ( .A(n620), .ZN(n600) );
  XOR2_X1 U681 ( .A(n672), .B(KEYINPUT78), .Z(n612) );
  INV_X1 U682 ( .A(n650), .ZN(n648) );
  OR2_X1 U683 ( .A1(n648), .A2(n602), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n659), .A2(n649), .ZN(n647) );
  NOR2_X1 U685 ( .A1(n606), .A2(n647), .ZN(n604) );
  XNOR2_X1 U686 ( .A(KEYINPUT93), .B(KEYINPUT31), .ZN(n603) );
  XNOR2_X1 U687 ( .A(n604), .B(n603), .ZN(n605) );
  XOR2_X1 U688 ( .A(KEYINPUT92), .B(n605), .Z(n640) );
  NOR2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U690 ( .A(n608), .B(KEYINPUT89), .ZN(n609) );
  NOR2_X1 U691 ( .A1(n659), .A2(n609), .ZN(n610) );
  XNOR2_X1 U692 ( .A(KEYINPUT91), .B(n610), .ZN(n622) );
  NAND2_X1 U693 ( .A1(n640), .A2(n622), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U695 ( .A(n617), .B(n616), .Z(n618) );
  XOR2_X1 U696 ( .A(KEYINPUT63), .B(n619), .Z(G57) );
  XOR2_X1 U697 ( .A(G101), .B(n620), .Z(G3) );
  NOR2_X1 U698 ( .A1(n637), .A2(n622), .ZN(n621) );
  XOR2_X1 U699 ( .A(G104), .B(n621), .Z(G6) );
  INV_X1 U700 ( .A(n628), .ZN(n639) );
  NOR2_X1 U701 ( .A1(n639), .A2(n622), .ZN(n624) );
  XNOR2_X1 U702 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U704 ( .A(G107), .B(n625), .ZN(G9) );
  XOR2_X1 U705 ( .A(G110), .B(n626), .Z(n627) );
  XNOR2_X1 U706 ( .A(KEYINPUT110), .B(n627), .ZN(G12) );
  XOR2_X1 U707 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n630) );
  NAND2_X1 U708 ( .A1(n634), .A2(n628), .ZN(n629) );
  XNOR2_X1 U709 ( .A(n630), .B(n629), .ZN(n631) );
  XOR2_X1 U710 ( .A(G128), .B(n631), .Z(G30) );
  XOR2_X1 U711 ( .A(G143), .B(n632), .Z(G45) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U713 ( .A(n635), .B(KEYINPUT112), .ZN(n636) );
  XNOR2_X1 U714 ( .A(G146), .B(n636), .ZN(G48) );
  NOR2_X1 U715 ( .A1(n640), .A2(n637), .ZN(n638) );
  XOR2_X1 U716 ( .A(G113), .B(n638), .Z(G15) );
  NOR2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U718 ( .A(G116), .B(n641), .Z(G18) );
  XNOR2_X1 U719 ( .A(G125), .B(n642), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n643), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U721 ( .A(G134), .B(n644), .Z(G36) );
  XNOR2_X1 U722 ( .A(G140), .B(n645), .ZN(G42) );
  NOR2_X1 U723 ( .A1(n664), .A2(n675), .ZN(n646) );
  NOR2_X1 U724 ( .A1(G953), .A2(n646), .ZN(n685) );
  NOR2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n661) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n652) );
  XNOR2_X1 U727 ( .A(KEYINPUT113), .B(KEYINPUT50), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n652), .B(n651), .ZN(n657) );
  NAND2_X1 U729 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U730 ( .A(KEYINPUT49), .B(n655), .Z(n656) );
  NAND2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U734 ( .A(KEYINPUT51), .B(n662), .Z(n663) );
  NOR2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U736 ( .A(KEYINPUT114), .B(n665), .ZN(n679) );
  NOR2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U738 ( .A(KEYINPUT115), .B(n668), .Z(n669) );
  NOR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n676) );
  NOR2_X1 U742 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U743 ( .A(KEYINPUT116), .B(n677), .ZN(n678) );
  NOR2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U745 ( .A(n680), .B(KEYINPUT52), .ZN(n681) );
  XNOR2_X1 U746 ( .A(n681), .B(KEYINPUT117), .ZN(n683) );
  NAND2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n692) );
  NOR2_X1 U749 ( .A1(KEYINPUT2), .A2(n732), .ZN(n686) );
  XNOR2_X1 U750 ( .A(n686), .B(KEYINPUT79), .ZN(n688) );
  NAND2_X1 U751 ( .A1(KEYINPUT2), .A2(n356), .ZN(n687) );
  NAND2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n690) );
  NOR2_X1 U753 ( .A1(KEYINPUT2), .A2(n718), .ZN(n689) );
  NOR2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U756 ( .A(KEYINPUT53), .B(n693), .ZN(G75) );
  NAND2_X1 U757 ( .A1(n715), .A2(G210), .ZN(n696) );
  XNOR2_X1 U758 ( .A(n694), .B(n412), .ZN(n695) );
  XNOR2_X1 U759 ( .A(KEYINPUT56), .B(n698), .ZN(G51) );
  NAND2_X1 U760 ( .A1(n715), .A2(G469), .ZN(n703) );
  XOR2_X1 U761 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n701) );
  XNOR2_X1 U762 ( .A(KEYINPUT119), .B(KEYINPUT118), .ZN(n700) );
  XNOR2_X1 U763 ( .A(KEYINPUT120), .B(n705), .ZN(G54) );
  XNOR2_X1 U764 ( .A(KEYINPUT121), .B(KEYINPUT83), .ZN(n708) );
  XNOR2_X1 U765 ( .A(n706), .B(KEYINPUT59), .ZN(n707) );
  XOR2_X1 U766 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n711) );
  NAND2_X1 U767 ( .A1(n715), .A2(G478), .ZN(n710) );
  XNOR2_X1 U768 ( .A(n711), .B(n710), .ZN(n713) );
  XNOR2_X1 U769 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U770 ( .A1(n717), .A2(n714), .ZN(G63) );
  NAND2_X1 U771 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U772 ( .A1(G953), .A2(G224), .ZN(n720) );
  XNOR2_X1 U773 ( .A(KEYINPUT61), .B(n720), .ZN(n721) );
  NAND2_X1 U774 ( .A1(n721), .A2(G898), .ZN(n722) );
  NAND2_X1 U775 ( .A1(n723), .A2(n722), .ZN(n728) );
  XNOR2_X1 U776 ( .A(n724), .B(G110), .ZN(n725) );
  NOR2_X1 U777 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U778 ( .A(n728), .B(n727), .ZN(G69) );
  XOR2_X1 U779 ( .A(n730), .B(n729), .Z(n731) );
  XNOR2_X1 U780 ( .A(KEYINPUT126), .B(n731), .ZN(n735) );
  XOR2_X1 U781 ( .A(n735), .B(n732), .Z(n734) );
  NAND2_X1 U782 ( .A1(n734), .A2(n733), .ZN(n739) );
  XNOR2_X1 U783 ( .A(G227), .B(n735), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U785 ( .A1(G953), .A2(n737), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n739), .A2(n738), .ZN(G72) );
  XOR2_X1 U787 ( .A(G122), .B(n740), .Z(n741) );
  XNOR2_X1 U788 ( .A(n741), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U789 ( .A(n742), .B(G119), .Z(G21) );
  XOR2_X1 U790 ( .A(n743), .B(G131), .Z(G33) );
  XOR2_X1 U791 ( .A(G137), .B(n744), .Z(G39) );
endmodule

