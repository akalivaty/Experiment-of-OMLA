//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G224), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(G143), .B2(new_n193), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n198), .A2(KEYINPUT65), .A3(G146), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n195), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT0), .A2(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n198), .A2(G146), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT64), .B1(new_n193), .B2(G143), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n198), .A3(G146), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n202), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n201), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI22_X1  g023(.A1(new_n200), .A2(new_n201), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G125), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n195), .B(new_n213), .C1(new_n197), .C2(new_n199), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n193), .A2(G143), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n215), .B2(KEYINPUT1), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n206), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n211), .B1(G125), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n218), .A2(KEYINPUT88), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT88), .B1(new_n210), .B2(G125), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n192), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n219), .A2(new_n192), .A3(new_n220), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n225));
  INV_X1    g039(.A(G104), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT80), .A2(G104), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n230));
  INV_X1    g044(.A(G101), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT80), .A2(G104), .ZN(new_n232));
  NOR2_X1   g046(.A1(KEYINPUT80), .A2(G104), .ZN(new_n233));
  OAI21_X1  g047(.A(G107), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n226), .A2(G107), .ZN(new_n235));
  AND2_X1   g049(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n230), .A2(new_n231), .A3(new_n234), .A4(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT2), .ZN(new_n241));
  INV_X1    g055(.A(G113), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n243), .A2(new_n244), .B1(KEYINPUT2), .B2(G113), .ZN(new_n245));
  INV_X1    g059(.A(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G116), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G119), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n248), .A2(G119), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT5), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n242), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT5), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n245), .A2(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n232), .A2(new_n233), .A3(G107), .ZN(new_n256));
  INV_X1    g070(.A(G107), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G104), .ZN(new_n258));
  OAI21_X1  g072(.A(G101), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n239), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(KEYINPUT86), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT3), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n232), .A2(new_n233), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(new_n257), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n238), .A2(new_n234), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n262), .B(G101), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT83), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n234), .B(new_n238), .C1(new_n256), .C2(new_n263), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT83), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n262), .A4(G101), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n257), .A2(G104), .ZN(new_n272));
  OR2_X1    g086(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g087(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n257), .B1(new_n227), .B2(new_n228), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n231), .B1(new_n277), .B2(new_n230), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT4), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(G101), .B1(new_n265), .B2(new_n266), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT82), .B1(new_n281), .B2(new_n239), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n268), .B(new_n271), .C1(new_n280), .C2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n245), .B(new_n250), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n261), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(G110), .B(G122), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n287), .B(KEYINPUT87), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT6), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT86), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n260), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n268), .A2(new_n271), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n269), .A2(G101), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n279), .B1(new_n295), .B2(new_n278), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n262), .B1(new_n281), .B2(KEYINPUT82), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n293), .B1(new_n298), .B2(new_n284), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n290), .A2(new_n291), .B1(new_n299), .B2(new_n287), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n296), .A2(new_n297), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n268), .A2(new_n271), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n284), .ZN(new_n303));
  AOI211_X1 g117(.A(new_n291), .B(new_n288), .C1(new_n303), .C2(new_n261), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n224), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT7), .B1(new_n191), .B2(G953), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n219), .A2(new_n220), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n287), .B(KEYINPUT8), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n239), .A2(new_n259), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(new_n255), .ZN(new_n311));
  INV_X1    g125(.A(new_n260), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n218), .A2(new_n307), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n303), .A2(new_n261), .A3(new_n287), .ZN(new_n317));
  AOI21_X1  g131(.A(G902), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n190), .B1(new_n306), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n223), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n221), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n288), .B1(new_n303), .B2(new_n261), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n317), .B1(new_n323), .B2(KEYINPUT6), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n324), .B2(new_n304), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n189), .A3(new_n318), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n188), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G221), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT9), .B(G234), .Z(new_n329));
  INV_X1    g143(.A(G902), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT11), .ZN(new_n333));
  INV_X1    g147(.A(G134), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(G137), .ZN(new_n335));
  INV_X1    g149(.A(G137), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT11), .A3(G134), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(G137), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G131), .ZN(new_n340));
  INV_X1    g154(.A(G131), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n335), .A2(new_n337), .A3(new_n341), .A4(new_n338), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n204), .B1(new_n198), .B2(G146), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n193), .A2(KEYINPUT64), .A3(G143), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n215), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n216), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT65), .B1(new_n198), .B2(G146), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n196), .A2(new_n193), .A3(G143), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n194), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n346), .A2(new_n347), .B1(new_n350), .B2(new_n213), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n214), .B1(new_n350), .B2(new_n216), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n239), .A2(new_n354), .A3(new_n259), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n310), .A2(new_n353), .B1(new_n355), .B2(new_n352), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n343), .B(new_n356), .C1(new_n283), .C2(new_n210), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n340), .A2(new_n342), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n239), .A2(new_n354), .A3(new_n259), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n217), .B1(new_n239), .B2(new_n259), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT12), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT12), .B(new_n358), .C1(new_n359), .C2(new_n360), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n357), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT84), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n357), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G953), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G227), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(KEYINPUT79), .ZN(new_n372));
  XNOR2_X1  g186(.A(G110), .B(G140), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n367), .A2(new_n369), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n374), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n357), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n207), .A2(new_n208), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n346), .A2(new_n378), .B1(new_n350), .B2(new_n207), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n301), .A2(new_n302), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n343), .B1(new_n380), .B2(new_n356), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n375), .A2(G469), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n357), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n374), .B1(new_n385), .B2(new_n381), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n357), .A2(new_n365), .A3(new_n376), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT72), .B(G902), .Z(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT85), .B(G469), .Z(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(G469), .A2(G902), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(G475), .A2(G902), .ZN(new_n395));
  XNOR2_X1  g209(.A(G113), .B(G122), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(new_n226), .ZN(new_n397));
  INV_X1    g211(.A(G237), .ZN(new_n398));
  AND4_X1   g212(.A1(G143), .A2(new_n398), .A3(new_n370), .A4(G214), .ZN(new_n399));
  NOR2_X1   g213(.A1(G237), .A2(G953), .ZN(new_n400));
  AOI21_X1  g214(.A(G143), .B1(new_n400), .B2(G214), .ZN(new_n401));
  OAI21_X1  g215(.A(G131), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT17), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n398), .A2(new_n370), .A3(G214), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n198), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n400), .A2(G143), .A3(G214), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n341), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT16), .ZN(new_n409));
  INV_X1    g223(.A(G140), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(G125), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT75), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT75), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n413), .A2(new_n409), .A3(new_n410), .A4(G125), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(G125), .ZN(new_n415));
  INV_X1    g229(.A(G125), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G140), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n412), .B(new_n414), .C1(new_n418), .C2(new_n409), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n193), .ZN(new_n420));
  XNOR2_X1  g234(.A(G125), .B(G140), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT16), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n422), .A2(G146), .A3(new_n412), .A4(new_n414), .ZN(new_n423));
  OAI211_X1 g237(.A(KEYINPUT17), .B(G131), .C1(new_n399), .C2(new_n401), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n408), .A2(new_n420), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT90), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n399), .A2(new_n401), .ZN(new_n427));
  NAND2_X1  g241(.A1(KEYINPUT18), .A2(G131), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n415), .A2(new_n417), .A3(new_n193), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n416), .A2(G140), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n410), .A2(G125), .ZN(new_n431));
  OAI21_X1  g245(.A(G146), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n427), .A2(new_n428), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(KEYINPUT18), .B(G131), .C1(new_n399), .C2(new_n401), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n426), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n429), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n405), .A2(new_n406), .A3(new_n428), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n434), .A2(new_n436), .A3(new_n426), .A4(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n397), .B(new_n425), .C1(new_n435), .C2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT90), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n438), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n418), .A2(KEYINPUT19), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT19), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n421), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n447), .A3(new_n193), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT91), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n402), .A2(new_n407), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT91), .A4(new_n193), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n450), .A2(new_n423), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n397), .B1(new_n444), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n395), .B1(new_n441), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(KEYINPUT20), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n450), .A2(new_n452), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n451), .A2(new_n423), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n459), .A2(new_n460), .B1(new_n438), .B2(new_n443), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n440), .B1(new_n461), .B2(new_n397), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n458), .B1(new_n462), .B2(new_n395), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n212), .A2(G143), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n198), .A2(G128), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n334), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n198), .A2(G128), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n212), .A2(G143), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(G134), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT13), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n471), .A3(G134), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G122), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G116), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n248), .A2(G122), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n475), .A2(new_n476), .A3(G107), .ZN(new_n477));
  AOI21_X1  g291(.A(G107), .B1(new_n475), .B2(new_n476), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n468), .A2(new_n469), .A3(new_n471), .A4(G134), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n473), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT92), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT92), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n473), .A2(new_n479), .A3(new_n483), .A4(new_n480), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n248), .A2(G122), .ZN(new_n486));
  NAND2_X1  g300(.A1(KEYINPUT14), .A2(G107), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n477), .A2(new_n478), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G116), .B(G122), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(KEYINPUT14), .A3(G107), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n467), .A3(new_n470), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT93), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n475), .A2(new_n476), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n257), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n490), .A2(G107), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n495), .B(new_n496), .C1(new_n486), .C2(new_n487), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n467), .A2(new_n470), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n491), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n329), .A2(G217), .A3(new_n370), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n485), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n485), .B2(new_n501), .ZN(new_n505));
  OAI211_X1 g319(.A(KEYINPUT94), .B(new_n390), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n485), .A2(new_n501), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n502), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n485), .A2(new_n501), .A3(new_n503), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n508), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n513), .A2(KEYINPUT94), .A3(new_n390), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n397), .B1(new_n444), .B2(new_n425), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n330), .B1(new_n441), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G475), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G952), .ZN(new_n521));
  AOI211_X1 g335(.A(G953), .B(new_n521), .C1(G234), .C2(G237), .ZN(new_n522));
  AOI211_X1 g336(.A(new_n370), .B(new_n390), .C1(G234), .C2(G237), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT21), .B(G898), .Z(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n522), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NOR4_X1   g340(.A1(new_n464), .A2(new_n516), .A3(new_n520), .A4(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n327), .A2(new_n332), .A3(new_n394), .A4(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT76), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n420), .A2(new_n423), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT23), .B1(new_n212), .B2(G119), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT73), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n246), .A2(G128), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT23), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n533), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n246), .A2(G128), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT23), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n539), .B(new_n542), .C1(KEYINPUT73), .C2(new_n534), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(G110), .A3(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT24), .B(G110), .Z(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n540), .A3(new_n535), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n531), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n545), .B1(new_n540), .B2(new_n535), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n541), .A2(new_n543), .ZN(new_n549));
  INV_X1    g363(.A(G110), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n423), .A2(new_n429), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT22), .B(G137), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n370), .A2(G221), .A3(G234), .ZN(new_n555));
  XOR2_X1   g369(.A(new_n554), .B(new_n555), .Z(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n547), .B(new_n556), .C1(new_n551), .C2(new_n552), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n390), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT25), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n558), .A2(KEYINPUT25), .A3(new_n390), .A4(new_n559), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G217), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(new_n390), .B2(G234), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n530), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n566), .ZN(new_n568));
  AOI211_X1 g382(.A(KEYINPUT76), .B(new_n568), .C1(new_n562), .C2(new_n563), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n566), .A2(G902), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n558), .A2(new_n559), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n567), .A2(new_n569), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(G472), .A2(G902), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT28), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n334), .A2(G137), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n336), .A2(G134), .ZN(new_n580));
  OAI21_X1  g394(.A(G131), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n342), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n358), .A2(new_n379), .B1(new_n217), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n285), .B1(new_n584), .B2(KEYINPUT67), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n379), .A2(new_n358), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n217), .A2(new_n583), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT67), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n578), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT68), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n584), .A2(new_n285), .ZN(new_n592));
  OAI22_X1  g406(.A1(new_n343), .A2(new_n210), .B1(new_n351), .B2(new_n582), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n284), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT28), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT67), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n285), .A3(new_n588), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT68), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n578), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n591), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n400), .A2(G210), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT30), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n593), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT30), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n284), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n592), .A3(new_n606), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT31), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n608), .A2(KEYINPUT69), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT69), .B1(new_n608), .B2(new_n615), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n577), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT32), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT69), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n284), .B1(new_n593), .B2(new_n597), .ZN(new_n622));
  AOI211_X1 g436(.A(KEYINPUT68), .B(KEYINPUT28), .C1(new_n622), .C2(new_n588), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n600), .B1(new_n599), .B2(new_n578), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n606), .B1(new_n625), .B2(new_n596), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n613), .B(KEYINPUT31), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n621), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n608), .A2(new_n615), .A3(KEYINPUT69), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(KEYINPUT32), .A3(new_n577), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT70), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n623), .B2(new_n624), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n591), .A2(KEYINPUT70), .A3(new_n601), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n607), .B1(new_n595), .B2(KEYINPUT28), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n635), .A2(KEYINPUT29), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT71), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n625), .A2(new_n635), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n612), .A2(new_n592), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT29), .B1(new_n640), .B2(new_n607), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n389), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n637), .A2(KEYINPUT71), .ZN(new_n644));
  OAI21_X1  g458(.A(G472), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n620), .A2(new_n631), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n529), .A2(new_n576), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G101), .ZN(G3));
  NAND2_X1  g462(.A1(new_n320), .A2(new_n326), .ZN(new_n649));
  INV_X1    g463(.A(new_n526), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT33), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n504), .B2(new_n505), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n511), .A2(KEYINPUT33), .A3(new_n512), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(new_n390), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G478), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n513), .A2(new_n507), .A3(new_n390), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n519), .B1(new_n456), .B2(new_n463), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n649), .A2(new_n187), .A3(new_n650), .A4(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n389), .B1(new_n628), .B2(new_n629), .ZN(new_n661));
  INV_X1    g475(.A(G472), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n618), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n394), .A2(new_n576), .A3(new_n332), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT34), .B(G104), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G6));
  AND3_X1   g481(.A1(new_n325), .A2(new_n189), .A3(new_n318), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n189), .B1(new_n325), .B2(new_n318), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n187), .B(new_n650), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n455), .A2(new_n457), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT95), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n462), .A2(new_n458), .A3(new_n395), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n455), .A2(KEYINPUT95), .A3(new_n457), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n516), .A2(new_n674), .A3(new_n519), .A4(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT96), .B1(new_n670), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT96), .ZN(new_n678));
  INV_X1    g492(.A(new_n676), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n327), .A2(new_n678), .A3(new_n650), .A4(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n376), .B1(new_n366), .B2(KEYINPUT84), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n382), .B1(new_n682), .B2(new_n369), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n389), .B1(new_n386), .B2(new_n387), .ZN(new_n684));
  AOI22_X1  g498(.A1(new_n683), .A2(G469), .B1(new_n684), .B2(new_n391), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n331), .B1(new_n685), .B2(new_n393), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n390), .B1(new_n616), .B2(new_n617), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G472), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n686), .A2(new_n688), .A3(new_n576), .A4(new_n618), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n681), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G107), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G9));
  NAND2_X1  g507(.A1(new_n564), .A2(new_n566), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT76), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n564), .A2(new_n530), .A3(new_n566), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n557), .A2(KEYINPUT36), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n553), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n573), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n695), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n618), .B(new_n700), .C1(new_n661), .C2(new_n662), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n528), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT98), .B(KEYINPUT37), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G110), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n702), .B(new_n704), .ZN(G12));
  NAND2_X1  g519(.A1(new_n394), .A2(new_n332), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n187), .B1(new_n668), .B2(new_n669), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(G900), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n522), .B1(new_n523), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n676), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n646), .A2(new_n708), .A3(new_n700), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G128), .ZN(G30));
  XOR2_X1   g527(.A(new_n710), .B(KEYINPUT39), .Z(new_n714));
  NAND2_X1  g528(.A1(new_n686), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT40), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n649), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n658), .A2(new_n516), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n720), .A2(new_n188), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n700), .ZN(new_n723));
  INV_X1    g537(.A(new_n613), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n595), .B2(new_n607), .ZN(new_n725));
  OAI21_X1  g539(.A(G472), .B1(new_n725), .B2(G902), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n620), .A2(new_n631), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n717), .A2(new_n722), .A3(new_n723), .A4(new_n727), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n728), .A2(KEYINPUT100), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(KEYINPUT100), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G143), .ZN(G45));
  INV_X1    g546(.A(new_n710), .ZN(new_n733));
  AND4_X1   g547(.A1(new_n658), .A2(new_n655), .A3(new_n656), .A4(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n646), .A2(new_n708), .A3(new_n700), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  INV_X1    g550(.A(new_n660), .ZN(new_n737));
  INV_X1    g551(.A(G469), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n392), .B(new_n332), .C1(new_n738), .C2(new_n684), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n737), .A2(new_n646), .A3(new_n576), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  NAND3_X1  g557(.A1(new_n646), .A2(new_n576), .A3(new_n740), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n681), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n248), .ZN(G18));
  NAND2_X1  g560(.A1(new_n700), .A2(new_n527), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n707), .A2(new_n747), .A3(new_n739), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n646), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  NAND2_X1  g564(.A1(new_n576), .A2(KEYINPUT101), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n633), .A2(new_n596), .A3(new_n634), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n615), .B1(new_n752), .B2(new_n606), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n577), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n695), .A2(new_n696), .A3(new_n574), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT101), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND4_X1   g571(.A1(new_n688), .A2(new_n751), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n721), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n650), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n707), .A2(new_n739), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  NOR2_X1   g577(.A1(new_n707), .A2(new_n739), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n687), .A2(G472), .B1(new_n577), .B2(new_n753), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n764), .A2(new_n700), .A3(new_n765), .A4(new_n734), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G125), .ZN(G27));
  AND2_X1   g581(.A1(new_n751), .A2(new_n757), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n393), .B(KEYINPUT102), .Z(new_n769));
  NAND3_X1  g583(.A1(new_n384), .A2(new_n392), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n332), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n320), .A2(new_n187), .A3(new_n326), .A4(new_n734), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AND4_X1   g587(.A1(KEYINPUT42), .A2(new_n768), .A3(new_n646), .A4(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n646), .A2(new_n773), .A3(new_n576), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT42), .B1(new_n775), .B2(KEYINPUT103), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT103), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n646), .A2(new_n773), .A3(new_n777), .A4(new_n576), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n774), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n341), .ZN(G33));
  NAND3_X1  g594(.A1(new_n320), .A2(new_n187), .A3(new_n326), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT104), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n676), .B2(new_n710), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n674), .A2(new_n675), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n520), .B1(new_n515), .B2(new_n509), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(KEYINPUT104), .A3(new_n785), .A4(new_n733), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n781), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n771), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n646), .A2(new_n576), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  OR2_X1    g605(.A1(new_n683), .A2(KEYINPUT45), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n683), .A2(KEYINPUT45), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(G469), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n769), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT46), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT105), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n769), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n392), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT105), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n795), .A2(new_n801), .A3(new_n796), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n798), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n331), .ZN(new_n805));
  INV_X1    g619(.A(new_n658), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n657), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT106), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(KEYINPUT43), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n657), .A2(new_n806), .B1(new_n808), .B2(KEYINPUT43), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n810), .B1(new_n811), .B2(new_n809), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(KEYINPUT107), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n663), .B(new_n700), .C1(new_n814), .C2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT44), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n781), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n805), .A2(new_n819), .A3(new_n714), .A4(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(KEYINPUT108), .B(G137), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(G39));
  OAI21_X1  g637(.A(KEYINPUT47), .B1(new_n804), .B2(new_n331), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n803), .A2(new_n825), .A3(new_n332), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n646), .A2(new_n576), .A3(new_n772), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  OAI21_X1  g643(.A(new_n392), .B1(new_n738), .B2(new_n684), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n807), .A2(new_n188), .A3(new_n331), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n727), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n720), .A3(new_n835), .A4(new_n768), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n776), .A2(new_n778), .ZN(new_n837));
  INV_X1    g651(.A(new_n774), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n758), .A2(new_n761), .B1(new_n748), .B2(new_n646), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n741), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n745), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n839), .A2(new_n842), .A3(KEYINPUT114), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n712), .A2(new_n766), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT110), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n712), .A2(KEYINPUT110), .A3(new_n766), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n770), .A2(new_n332), .A3(new_n733), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n187), .B(new_n759), .C1(new_n668), .C2(new_n669), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n727), .A3(new_n723), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n846), .A2(new_n735), .A3(new_n847), .A4(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n712), .A2(new_n735), .A3(new_n851), .A4(new_n766), .ZN(new_n854));
  XNOR2_X1  g668(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n665), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n520), .B(new_n464), .C1(new_n515), .C2(new_n509), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n327), .A2(new_n650), .A3(new_n859), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n689), .A2(new_n860), .B1(new_n528), .B2(new_n701), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n647), .B(new_n858), .C1(new_n861), .C2(KEYINPUT109), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT109), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n687), .A2(G472), .B1(new_n630), .B2(new_n577), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n708), .A2(new_n527), .A3(new_n864), .A4(new_n700), .ZN(new_n865));
  INV_X1    g679(.A(new_n664), .ZN(new_n866));
  INV_X1    g680(.A(new_n670), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n864), .A4(new_n859), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n863), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n516), .A2(new_n520), .A3(new_n710), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n700), .A2(new_n784), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n871), .A2(new_n781), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n646), .A2(new_n872), .A3(new_n686), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n773), .A2(new_n700), .A3(new_n765), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n790), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n862), .A2(new_n869), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n840), .B(new_n741), .C1(new_n681), .C2(new_n744), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n877), .B1(new_n779), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n843), .A2(new_n857), .A3(new_n876), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT53), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n790), .A2(new_n873), .A3(new_n874), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n646), .A2(new_n576), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n665), .B1(new_n883), .B2(new_n529), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n860), .A2(new_n663), .A3(new_n664), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT109), .B1(new_n885), .B2(new_n702), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n865), .A2(new_n868), .A3(new_n863), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n882), .A2(new_n884), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n888), .A2(new_n779), .A3(new_n878), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n854), .B(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT54), .B1(new_n881), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n720), .A2(new_n188), .A3(new_n740), .ZN(new_n895));
  INV_X1    g709(.A(new_n522), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n813), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n895), .A2(KEYINPUT50), .A3(new_n758), .A4(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT50), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n758), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n720), .A2(new_n188), .A3(new_n740), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n781), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n812), .A2(new_n904), .A3(new_n522), .A4(new_n740), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n765), .A2(new_n700), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT116), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT116), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n904), .A2(new_n576), .A3(new_n522), .A4(new_n740), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n727), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n657), .A2(new_n658), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n907), .A2(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n830), .A2(new_n332), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n824), .B2(new_n826), .ZN(new_n916));
  INV_X1    g730(.A(new_n900), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n904), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n913), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT51), .B1(new_n913), .B2(KEYINPUT115), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI221_X1 g735(.A(new_n913), .B1(KEYINPUT115), .B2(KEYINPUT51), .C1(new_n916), .C2(new_n918), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n917), .A2(new_n764), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n521), .B(G953), .C1(new_n910), .C2(new_n659), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n768), .A2(new_n646), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n925), .A2(new_n740), .A3(new_n904), .A4(new_n897), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT117), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT48), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n923), .B(new_n924), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n921), .A2(new_n922), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT112), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n889), .A2(new_n857), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(KEYINPUT53), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT53), .B1(new_n889), .B2(new_n857), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT112), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n779), .A2(new_n878), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n892), .A2(new_n938), .A3(KEYINPUT53), .A4(new_n876), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT113), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT113), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n889), .A2(new_n941), .A3(KEYINPUT53), .A4(new_n892), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n935), .A2(new_n937), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  AOI211_X1 g757(.A(new_n894), .B(new_n932), .C1(new_n943), .C2(KEYINPUT54), .ZN(new_n944));
  NOR2_X1   g758(.A1(G952), .A2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n836), .B1(new_n944), .B2(new_n945), .ZN(G75));
  NAND4_X1  g760(.A1(new_n881), .A2(new_n389), .A3(new_n190), .A4(new_n893), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT56), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n324), .A2(new_n304), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n224), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n325), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT118), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(KEYINPUT56), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n947), .A2(new_n948), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n947), .B2(new_n948), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n370), .A2(G952), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(G51));
  XOR2_X1   g772(.A(new_n769), .B(KEYINPUT57), .Z(new_n959));
  AND3_X1   g773(.A1(new_n881), .A2(KEYINPUT54), .A3(new_n893), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(new_n894), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n388), .B(KEYINPUT119), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n881), .A2(new_n389), .A3(new_n893), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n794), .B(KEYINPUT120), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n957), .B1(new_n963), .B2(new_n966), .ZN(G54));
  AND2_X1   g781(.A1(KEYINPUT58), .A2(G475), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n964), .A2(new_n462), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n462), .B1(new_n964), .B2(new_n968), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n957), .ZN(G60));
  NAND2_X1  g785(.A1(new_n652), .A2(new_n653), .ZN(new_n972));
  XNOR2_X1  g786(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n507), .A2(new_n330), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n960), .B2(new_n894), .ZN(new_n977));
  INV_X1    g791(.A(new_n957), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n940), .B(new_n942), .C1(KEYINPUT112), .C2(new_n936), .ZN(new_n980));
  INV_X1    g794(.A(new_n937), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT54), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n894), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n975), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n979), .B1(new_n986), .B2(new_n972), .ZN(G63));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(KEYINPUT123), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(KEYINPUT123), .ZN(new_n990));
  XNOR2_X1  g804(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n565), .A2(new_n330), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n881), .A2(new_n893), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n558), .A2(new_n559), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n881), .A2(new_n698), .A3(new_n893), .A4(new_n993), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n978), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n989), .B(new_n990), .C1(new_n996), .C2(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n997), .A2(new_n978), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n994), .A2(new_n995), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1000), .A2(KEYINPUT123), .A3(new_n988), .A4(new_n1001), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n999), .A2(new_n1002), .ZN(G66));
  OAI21_X1  g817(.A(G953), .B1(new_n525), .B2(new_n191), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n878), .A2(new_n862), .A3(new_n869), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n949), .B1(G898), .B2(new_n370), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1006), .B(new_n1007), .ZN(G69));
  AND3_X1   g822(.A1(new_n846), .A2(new_n735), .A3(new_n847), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n729), .A2(new_n1009), .A3(new_n730), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(KEYINPUT124), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1011), .A2(KEYINPUT124), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1012), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n828), .A2(new_n821), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n904), .B1(new_n659), .B2(new_n859), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n1018), .A2(new_n715), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n883), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n610), .A2(new_n611), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n445), .A2(new_n447), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1022), .B(new_n1023), .Z(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1025), .A2(G953), .ZN(new_n1026));
  AOI21_X1  g840(.A(KEYINPUT125), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(G227), .B1(new_n1025), .B2(KEYINPUT125), .ZN(new_n1028));
  OAI21_X1  g842(.A(G953), .B1(new_n1028), .B2(new_n709), .ZN(new_n1029));
  INV_X1    g843(.A(new_n849), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n805), .A2(new_n714), .A3(new_n925), .A4(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1031), .A2(new_n839), .A3(new_n790), .A4(new_n1009), .ZN(new_n1032));
  NOR3_X1   g846(.A1(new_n1032), .A2(new_n1016), .A3(G953), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n709), .A2(new_n370), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1025), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AND3_X1   g849(.A1(new_n1027), .A2(new_n1029), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1029), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1036), .A2(new_n1037), .ZN(G72));
  XNOR2_X1  g852(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n662), .A2(new_n330), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1005), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1041), .B1(new_n1021), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1043), .A2(new_n606), .A3(new_n640), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n606), .B1(new_n612), .B2(new_n592), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n943), .B(new_n1041), .C1(new_n724), .C2(new_n1045), .ZN(new_n1046));
  OR2_X1    g860(.A1(new_n1032), .A2(new_n1016), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1041), .B1(new_n1047), .B2(new_n1042), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n640), .A2(new_n606), .ZN(new_n1049));
  XNOR2_X1  g863(.A(new_n1049), .B(KEYINPUT127), .ZN(new_n1050));
  AOI21_X1  g864(.A(new_n957), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  AND3_X1   g865(.A1(new_n1044), .A2(new_n1046), .A3(new_n1051), .ZN(G57));
endmodule


