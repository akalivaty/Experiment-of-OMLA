//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  INV_X1    g001(.A(G116), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT67), .B1(new_n188), .B2(G119), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G119), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT2), .B(G113), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n189), .A2(new_n192), .A3(KEYINPUT68), .A4(new_n193), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT69), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n189), .A2(new_n192), .A3(new_n193), .ZN(new_n201));
  INV_X1    g015(.A(new_n197), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n200), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n194), .A2(KEYINPUT69), .A3(new_n197), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n199), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT70), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n200), .A3(new_n202), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT69), .B1(new_n194), .B2(new_n197), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT70), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(new_n199), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G137), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT11), .A3(G134), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n214), .A2(new_n216), .A3(new_n220), .A4(new_n217), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G143), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n223), .A2(KEYINPUT65), .A3(G146), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n224), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT0), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(G143), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n223), .A2(G146), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n233), .A2(new_n234), .B1(new_n230), .B2(new_n231), .ZN(new_n235));
  AND3_X1   g049(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n229), .A2(new_n232), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n234), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT66), .A2(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT66), .A2(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(G143), .B2(new_n226), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n240), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(G128), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n223), .A2(KEYINPUT65), .A3(G146), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT65), .B1(new_n223), .B2(G146), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n233), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n213), .A2(G137), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n215), .A2(G134), .ZN(new_n254));
  OAI21_X1  g068(.A(G131), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n221), .A2(new_n255), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n222), .A2(new_n239), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n206), .A2(new_n211), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n206), .A2(KEYINPUT71), .A3(new_n211), .A4(new_n257), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n239), .A2(new_n222), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n252), .A2(new_n256), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT30), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n264), .B1(new_n262), .B2(new_n263), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n209), .A2(new_n210), .A3(new_n199), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n210), .B1(new_n209), .B2(new_n199), .ZN(new_n268));
  OAI22_X1  g082(.A1(new_n265), .A2(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n260), .A2(new_n261), .A3(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT72), .B(KEYINPUT27), .Z(new_n271));
  NOR2_X1   g085(.A1(G237), .A2(G953), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G210), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n271), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G101), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n187), .B1(new_n270), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n258), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n277), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n206), .A2(new_n211), .ZN(new_n282));
  INV_X1    g096(.A(new_n257), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n260), .A2(new_n284), .A3(new_n261), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n281), .B1(new_n285), .B2(KEYINPUT28), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n278), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(KEYINPUT28), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n267), .A2(new_n268), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT28), .B1(new_n289), .B2(new_n257), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n290), .A2(new_n187), .A3(new_n276), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT73), .B(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G472), .B1(new_n287), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT31), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n270), .A2(new_n296), .A3(new_n277), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n260), .A2(new_n269), .A3(new_n261), .A4(new_n277), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT31), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n290), .B1(new_n285), .B2(KEYINPUT28), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n297), .B(new_n299), .C1(new_n300), .C2(new_n277), .ZN(new_n301));
  NOR2_X1   g115(.A1(G472), .A2(G902), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT32), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n288), .A2(new_n280), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n276), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n298), .B(new_n296), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n303), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n295), .B(new_n306), .C1(new_n310), .C2(KEYINPUT32), .ZN(new_n311));
  INV_X1    g125(.A(G217), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n293), .B2(G234), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  OR2_X1    g128(.A1(KEYINPUT66), .A2(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT66), .A2(G128), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n315), .A2(KEYINPUT23), .A3(G119), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n231), .A2(G119), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT23), .B1(new_n231), .B2(G119), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n317), .A2(KEYINPUT75), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n243), .A2(new_n321), .A3(KEYINPUT23), .A4(G119), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT78), .B(G110), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n231), .A2(G119), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n243), .B2(G119), .ZN(new_n326));
  INV_X1    g140(.A(G110), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT24), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT24), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G110), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n331), .B1(new_n328), .B2(new_n330), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI22_X1  g149(.A1(new_n323), .A2(new_n324), .B1(new_n326), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(KEYINPUT76), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(G125), .A3(G140), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(KEYINPUT16), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT16), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n338), .B2(G140), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G146), .ZN(new_n346));
  XNOR2_X1  g160(.A(G125), .B(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n226), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n336), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n327), .B1(new_n320), .B2(new_n322), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n226), .A3(new_n344), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n346), .A2(new_n352), .B1(new_n335), .B2(new_n326), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT77), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n334), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n326), .A2(new_n355), .A3(new_n332), .ZN(new_n356));
  INV_X1    g170(.A(new_n352), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n226), .B1(new_n342), .B2(new_n344), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n359), .A2(new_n350), .A3(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n349), .B1(new_n354), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT22), .B(G137), .ZN(new_n363));
  INV_X1    g177(.A(G953), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n364), .A2(G221), .A3(G234), .ZN(new_n365));
  XOR2_X1   g179(.A(new_n363), .B(new_n365), .Z(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n349), .B(new_n366), .C1(new_n354), .C2(new_n361), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n293), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT25), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n368), .A2(KEYINPUT25), .A3(new_n293), .A4(new_n369), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n314), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(new_n369), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n313), .A2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n311), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT92), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT9), .B(G234), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n382), .A2(new_n312), .A3(G953), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n384), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n315), .A2(G143), .A3(new_n316), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n223), .A2(G128), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n213), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT79), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G107), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G122), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G116), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n188), .A2(G122), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n395), .A2(new_n399), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n390), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT89), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT13), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n389), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n388), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n389), .A2(new_n404), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n388), .A2(new_n403), .A3(new_n405), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n402), .B1(new_n410), .B2(G134), .ZN(new_n411));
  AOI21_X1  g225(.A(KEYINPUT14), .B1(new_n396), .B2(G116), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n396), .A2(G116), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT90), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n398), .A2(KEYINPUT14), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT90), .ZN(new_n417));
  OAI21_X1  g231(.A(G107), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n388), .A2(new_n389), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G134), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n390), .ZN(new_n421));
  INV_X1    g235(.A(new_n401), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n418), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n381), .B(new_n387), .C1(new_n411), .C2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n402), .ZN(new_n425));
  INV_X1    g239(.A(new_n409), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n426), .A2(new_n406), .A3(new_n407), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n425), .B1(new_n427), .B2(new_n213), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n387), .A2(new_n381), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n385), .A2(KEYINPUT92), .A3(new_n386), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n418), .A2(new_n421), .A3(new_n422), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n428), .A2(new_n429), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT93), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n424), .A2(new_n432), .A3(new_n433), .A4(new_n293), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT15), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n434), .A2(new_n435), .A3(G478), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(G478), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n424), .A2(new_n432), .A3(new_n293), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT93), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n434), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n436), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n272), .A2(G143), .A3(G214), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(G143), .B1(new_n272), .B2(G214), .ZN(new_n445));
  OAI21_X1  g259(.A(G131), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n272), .A2(G214), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n223), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n220), .A3(new_n443), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n446), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT88), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n357), .A2(new_n358), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n446), .A2(new_n449), .A3(new_n454), .A4(new_n450), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n446), .A2(new_n450), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n452), .A2(new_n453), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G113), .B(G122), .ZN(new_n458));
  INV_X1    g272(.A(G104), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(KEYINPUT18), .A2(G131), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n444), .A2(new_n445), .A3(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n448), .A2(new_n443), .B1(KEYINPUT18), .B2(G131), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n339), .A2(G146), .A3(new_n341), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n348), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n465), .B2(new_n466), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n457), .A2(new_n460), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n464), .A2(new_n468), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT19), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n347), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n339), .A2(KEYINPUT19), .A3(new_n341), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n226), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n346), .A2(new_n475), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n476), .A2(KEYINPUT87), .B1(new_n446), .B2(new_n449), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n346), .A2(new_n478), .A3(new_n475), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n471), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n470), .B1(new_n480), .B2(new_n460), .ZN(new_n481));
  NOR2_X1   g295(.A1(G475), .A2(G902), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n442), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n442), .A3(new_n482), .ZN(new_n485));
  INV_X1    g299(.A(G902), .ZN(new_n486));
  INV_X1    g300(.A(new_n470), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n460), .B1(new_n457), .B2(new_n469), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n484), .A2(new_n485), .B1(G475), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G952), .ZN(new_n491));
  AOI211_X1 g305(.A(G953), .B(new_n491), .C1(G234), .C2(G237), .ZN(new_n492));
  AOI211_X1 g306(.A(new_n364), .B(new_n293), .C1(G234), .C2(G237), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT21), .B(G898), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n441), .A2(new_n490), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G469), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT3), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n391), .B1(new_n499), .B2(G104), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(G104), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n392), .A3(new_n394), .ZN(new_n504));
  INV_X1    g318(.A(G101), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(G104), .B2(G107), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n395), .B2(G104), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n229), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n245), .A2(KEYINPUT80), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G128), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n245), .A2(KEYINPUT80), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n509), .B1(new_n514), .B2(new_n251), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n252), .B1(new_n506), .B2(new_n508), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n222), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT12), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT10), .ZN(new_n519));
  INV_X1    g333(.A(new_n251), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n231), .B1(new_n245), .B2(KEYINPUT80), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(KEYINPUT80), .B2(new_n245), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n522), .B2(new_n510), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n519), .B1(new_n523), .B2(new_n509), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n502), .A2(new_n504), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G101), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(KEYINPUT4), .A3(new_n506), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT4), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n528), .A3(G101), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n239), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n222), .ZN(new_n531));
  INV_X1    g345(.A(new_n509), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(KEYINPUT10), .A3(new_n252), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n524), .A2(new_n530), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n535), .B(new_n222), .C1(new_n515), .C2(new_n516), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n518), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G110), .B(G140), .ZN(new_n538));
  INV_X1    g352(.A(G227), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(G953), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n538), .B(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n541), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n524), .A2(new_n530), .A3(new_n533), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n222), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n545), .B2(new_n534), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n498), .B(new_n293), .C1(new_n542), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n537), .A2(new_n541), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n534), .A3(new_n543), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(G469), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(G469), .A2(G902), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G221), .B1(new_n382), .B2(G902), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n497), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G214), .B1(G237), .B2(G902), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G122), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n527), .A2(new_n529), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n206), .B2(new_n211), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n532), .A2(new_n209), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT5), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n191), .A3(G116), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G113), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n196), .A2(new_n198), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(KEYINPUT5), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n559), .B1(new_n561), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n560), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n267), .B2(new_n268), .ZN(new_n571));
  INV_X1    g385(.A(new_n568), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n558), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n573), .A3(KEYINPUT6), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n246), .A2(new_n251), .A3(new_n338), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n235), .A2(new_n238), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n232), .B(new_n233), .C1(new_n249), .C2(new_n250), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n338), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT81), .B(G224), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n364), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n246), .A2(new_n251), .A3(new_n338), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n583), .B(new_n581), .C1(new_n239), .C2(new_n338), .ZN(new_n584));
  AND3_X1   g398(.A1(new_n582), .A2(KEYINPUT82), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT82), .B1(new_n582), .B2(new_n584), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT6), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n588), .B(new_n559), .C1(new_n561), .C2(new_n568), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n574), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT85), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n579), .A2(new_n591), .A3(KEYINPUT7), .A4(new_n581), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT7), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT85), .B1(new_n584), .B2(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT84), .B(KEYINPUT7), .Z(new_n595));
  NAND2_X1  g409(.A1(new_n581), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n575), .B2(new_n578), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n592), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n568), .B1(new_n282), .B2(new_n570), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n598), .B1(new_n599), .B2(new_n558), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n558), .B(KEYINPUT8), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n194), .A2(new_n563), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n532), .B(new_n209), .C1(new_n565), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT83), .ZN(new_n604));
  INV_X1    g418(.A(new_n209), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n509), .B1(new_n605), .B2(new_n567), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n603), .A2(KEYINPUT83), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n601), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n600), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n590), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G210), .B1(G237), .B2(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n590), .A2(new_n610), .A3(new_n612), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n557), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n555), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n380), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n505), .ZN(G3));
  AND3_X1   g433(.A1(new_n590), .A2(new_n610), .A3(new_n612), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n612), .B1(new_n590), .B2(new_n610), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n556), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(G478), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n438), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT96), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT94), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n385), .A2(new_n386), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n213), .B1(new_n408), .B2(new_n409), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n431), .B(new_n627), .C1(new_n628), .C2(new_n402), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT33), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n627), .B1(new_n428), .B2(new_n431), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT95), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n424), .A2(new_n432), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n627), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n411), .B2(new_n423), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT33), .A4(new_n629), .ZN(new_n638));
  INV_X1    g452(.A(new_n293), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n623), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n632), .A2(new_n634), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT96), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n438), .A2(new_n642), .A3(new_n623), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n625), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n489), .A2(G475), .ZN(new_n645));
  INV_X1    g459(.A(new_n482), .ZN(new_n646));
  INV_X1    g460(.A(new_n475), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT87), .B1(new_n647), .B2(new_n358), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n446), .A2(new_n449), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n479), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n469), .ZN(new_n651));
  INV_X1    g465(.A(new_n460), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI211_X1 g467(.A(KEYINPUT20), .B(new_n646), .C1(new_n653), .C2(new_n470), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n645), .B1(new_n654), .B2(new_n483), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n644), .A2(new_n655), .A3(new_n496), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n622), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n374), .A2(new_n378), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n554), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n301), .A2(new_n293), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n660), .A2(G472), .B1(new_n302), .B2(new_n301), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n657), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT34), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  AND2_X1   g478(.A1(new_n440), .A2(new_n437), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n490), .B(new_n496), .C1(new_n665), .C2(new_n436), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n622), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n659), .A3(new_n661), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT35), .B(G107), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  OR2_X1    g484(.A1(new_n367), .A2(KEYINPUT36), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n362), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n377), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n372), .A2(new_n373), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(new_n313), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n555), .A2(new_n661), .A3(new_n616), .A4(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  NOR2_X1   g493(.A1(new_n554), .A2(new_n675), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n490), .B1(new_n665), .B2(new_n436), .ZN(new_n681));
  INV_X1    g495(.A(new_n492), .ZN(new_n682));
  INV_X1    g496(.A(new_n493), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n682), .B1(new_n683), .B2(G900), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT97), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n311), .A2(new_n616), .A3(new_n680), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  OAI21_X1  g503(.A(new_n655), .B1(new_n665), .B2(new_n436), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n301), .A2(new_n302), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n304), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n260), .A2(new_n261), .A3(new_n269), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n277), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n694), .B(new_n486), .C1(new_n285), .C2(new_n277), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n301), .A2(new_n305), .B1(G472), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n690), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n556), .A3(new_n675), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n620), .A2(new_n621), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT38), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n685), .B(KEYINPUT39), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n552), .A2(new_n553), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT40), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n698), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT98), .B(G143), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G45));
  NAND3_X1  g520(.A1(new_n644), .A2(new_n655), .A3(new_n685), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT99), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(new_n311), .A3(new_n616), .A4(new_n680), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  NOR2_X1   g524(.A1(new_n542), .A2(new_n546), .ZN(new_n711));
  OAI21_X1  g525(.A(G469), .B1(new_n711), .B2(new_n639), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n553), .A3(new_n547), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n658), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n657), .A2(new_n714), .A3(new_n311), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NAND3_X1  g531(.A1(new_n667), .A2(new_n714), .A3(new_n311), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NOR2_X1   g533(.A1(new_n622), .A2(new_n713), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n497), .A2(new_n675), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n311), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  INV_X1    g537(.A(new_n713), .ZN(new_n724));
  INV_X1    g538(.A(new_n690), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n616), .A2(new_n724), .A3(new_n725), .A4(new_n496), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT100), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n661), .A2(new_n727), .A3(new_n379), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n639), .B1(new_n308), .B2(new_n309), .ZN(new_n729));
  INV_X1    g543(.A(G472), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n379), .B(new_n691), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT100), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n726), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n396), .ZN(G24));
  AOI21_X1  g548(.A(new_n730), .B1(new_n301), .B2(new_n293), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n735), .A2(new_n675), .A3(new_n310), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n708), .A2(new_n736), .A3(new_n720), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  NAND2_X1  g552(.A1(new_n306), .A2(KEYINPUT102), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n301), .A2(new_n740), .A3(new_n305), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n692), .A2(new_n739), .A3(new_n295), .A4(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n614), .A2(new_n556), .A3(new_n615), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT101), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n548), .B2(new_n549), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT101), .B1(new_n537), .B2(new_n541), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n745), .A2(new_n498), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n547), .A2(new_n551), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n553), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n742), .A2(new_n379), .A3(new_n708), .A4(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n750), .A2(new_n311), .A3(new_n379), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n708), .A2(new_n753), .ZN(new_n754));
  AOI22_X1  g568(.A1(KEYINPUT42), .A2(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  NAND4_X1  g570(.A1(new_n750), .A2(new_n311), .A3(new_n379), .A4(new_n687), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  NAND2_X1  g572(.A1(new_n548), .A2(new_n549), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n498), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n745), .A2(new_n746), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n761), .B1(new_n762), .B2(new_n760), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n551), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n764), .A2(KEYINPUT103), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT46), .B1(new_n763), .B2(new_n551), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT104), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n764), .A2(KEYINPUT103), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n547), .B1(new_n766), .B2(KEYINPUT104), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n553), .B(new_n701), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n490), .A2(new_n644), .ZN(new_n772));
  AND2_X1   g586(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n773));
  NOR2_X1   g587(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n772), .B2(new_n774), .ZN(new_n776));
  INV_X1    g590(.A(new_n661), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n676), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n743), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n779), .B2(new_n778), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n771), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n215), .ZN(G39));
  NOR3_X1   g597(.A1(new_n311), .A2(new_n379), .A3(new_n743), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(new_n708), .ZN(new_n785));
  OAI211_X1 g599(.A(KEYINPUT47), .B(new_n553), .C1(new_n769), .C2(new_n770), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n770), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(new_n765), .A3(new_n767), .A4(new_n768), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT47), .B1(new_n789), .B2(new_n553), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n785), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  NAND2_X1  g606(.A1(new_n692), .A2(new_n696), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n658), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n712), .A2(new_n547), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT49), .ZN(new_n796));
  INV_X1    g610(.A(new_n553), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n772), .A2(new_n557), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n700), .A2(new_n794), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n685), .B(KEYINPUT107), .Z(new_n801));
  OAI21_X1  g615(.A(KEYINPUT108), .B1(new_n676), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n622), .A2(new_n749), .ZN(new_n803));
  OR4_X1    g617(.A1(KEYINPUT108), .A2(new_n374), .A3(new_n673), .A4(new_n801), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n697), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n709), .A3(new_n737), .A4(new_n688), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT52), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n715), .A2(new_n718), .A3(new_n722), .A4(new_n677), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n662), .B1(new_n380), .B2(new_n617), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT106), .B1(new_n622), .B2(new_n666), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT106), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n441), .A2(new_n495), .A3(new_n655), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n616), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n811), .A2(new_n814), .A3(new_n661), .A4(new_n659), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n733), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n708), .A2(new_n750), .A3(new_n736), .ZN(new_n818));
  INV_X1    g632(.A(new_n743), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n441), .A2(new_n490), .A3(new_n685), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n311), .A2(new_n819), .A3(new_n680), .A4(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n757), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n810), .A2(new_n755), .A3(new_n817), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n800), .B1(new_n807), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n755), .A2(new_n822), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n737), .A2(new_n688), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(KEYINPUT52), .A3(new_n709), .A4(new_n805), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n806), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n726), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n727), .B1(new_n661), .B2(new_n379), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n731), .A2(KEYINPUT100), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n815), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n835), .A2(new_n809), .A3(new_n808), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n825), .A2(new_n830), .A3(new_n836), .A4(KEYINPUT53), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n824), .A2(KEYINPUT110), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n823), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT110), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT53), .A4(new_n830), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g656(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n843));
  INV_X1    g657(.A(KEYINPUT109), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n837), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n839), .A2(KEYINPUT109), .A3(KEYINPUT53), .A4(new_n830), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n846), .A3(new_n824), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n842), .A2(new_n843), .B1(new_n847), .B2(KEYINPUT54), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n776), .A2(new_n492), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n819), .A2(new_n724), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR4_X1   g665(.A1(new_n850), .A2(new_n793), .A3(new_n658), .A4(new_n682), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n644), .A2(new_n655), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n736), .A2(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n724), .A2(new_n557), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n855), .A2(KEYINPUT114), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(KEYINPUT114), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n856), .A2(new_n700), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n849), .B1(new_n728), .B2(new_n732), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n858), .A2(KEYINPUT50), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT50), .B1(new_n858), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n854), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n553), .B1(new_n769), .B2(new_n770), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT47), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n795), .A2(KEYINPUT112), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n795), .A2(KEYINPUT112), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n797), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n786), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n859), .A2(new_n819), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n862), .A2(new_n863), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n864), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n742), .A2(new_n379), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n851), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT48), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n859), .A2(new_n720), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n644), .A2(new_n655), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n491), .B(G953), .C1(new_n852), .C2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n871), .A2(new_n873), .B1(new_n872), .B2(new_n877), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n862), .A2(KEYINPUT51), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n848), .A2(new_n878), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n799), .B1(new_n890), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n364), .A2(G952), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT116), .Z(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n842), .A2(new_n293), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n613), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n574), .A2(new_n589), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(new_n587), .Z(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n897), .A2(new_n898), .A3(new_n902), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n895), .B1(new_n904), .B2(new_n905), .ZN(G51));
  XOR2_X1   g720(.A(new_n711), .B(KEYINPUT117), .Z(new_n907));
  NAND2_X1  g721(.A1(new_n842), .A2(new_n843), .ZN(new_n908));
  INV_X1    g722(.A(new_n843), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n838), .A2(new_n841), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n551), .B(KEYINPUT57), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n907), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n763), .B(KEYINPUT118), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n896), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n893), .B1(new_n914), .B2(new_n916), .ZN(G54));
  AND2_X1   g731(.A1(KEYINPUT58), .A2(G475), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n838), .A2(new_n639), .A3(new_n841), .A4(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n481), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n893), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n920), .B2(new_n919), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT119), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n921), .B(new_n924), .C1(new_n920), .C2(new_n919), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(G60));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n847), .A2(KEYINPUT54), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n908), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n632), .A2(new_n634), .A3(new_n638), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n927), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(KEYINPUT120), .B(new_n932), .C1(new_n848), .C2(new_n929), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n932), .A2(new_n929), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n895), .B1(new_n911), .B2(new_n936), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT121), .Z(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n842), .A2(new_n672), .A3(new_n941), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n375), .B(KEYINPUT122), .Z(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n842), .B2(new_n941), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n894), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n942), .A2(KEYINPUT61), .A3(new_n894), .A4(new_n944), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n494), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n364), .B1(new_n950), .B2(new_n580), .ZN(new_n951));
  INV_X1    g765(.A(new_n836), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n364), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n900), .B1(G898), .B2(new_n364), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n953), .B(new_n954), .Z(G69));
  NAND2_X1  g769(.A1(new_n867), .A2(new_n786), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n782), .B1(new_n956), .B2(new_n785), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n826), .A2(new_n709), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  OR3_X1    g773(.A1(new_n958), .A2(new_n959), .A3(new_n704), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n958), .B2(new_n704), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n702), .B1(new_n883), .B2(new_n681), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n819), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT124), .B1(new_n963), .B2(new_n380), .ZN(new_n964));
  OR3_X1    g778(.A1(new_n963), .A2(new_n380), .A3(KEYINPUT124), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n960), .A2(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n957), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n265), .A2(new_n266), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT123), .Z(new_n969));
  NAND2_X1  g783(.A1(new_n473), .A2(new_n474), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n967), .A2(new_n364), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(G900), .ZN(new_n973));
  INV_X1    g787(.A(new_n771), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n974), .A2(new_n616), .A3(new_n725), .A4(new_n879), .ZN(new_n975));
  INV_X1    g789(.A(new_n782), .ZN(new_n976));
  AND4_X1   g790(.A1(new_n709), .A2(new_n755), .A3(new_n757), .A4(new_n826), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n791), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  MUX2_X1   g792(.A(new_n973), .B(new_n978), .S(new_n364), .Z(new_n979));
  OAI21_X1  g793(.A(new_n972), .B1(new_n979), .B2(new_n971), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n364), .B1(G227), .B2(G900), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT125), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n980), .B(new_n982), .ZN(G72));
  NAND3_X1  g797(.A1(new_n957), .A2(new_n966), .A3(new_n836), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  NAND3_X1  g800(.A1(new_n984), .A2(KEYINPUT126), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n694), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT126), .B1(new_n984), .B2(new_n986), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n986), .B1(new_n978), .B2(new_n952), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n693), .A2(new_n277), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n893), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n993), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n847), .A2(new_n694), .A3(new_n986), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT127), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n990), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n988), .A3(new_n987), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT127), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1000), .A2(new_n1001), .A3(new_n996), .A4(new_n994), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n998), .A2(new_n1002), .ZN(G57));
endmodule


