//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND3_X1  g0013(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n203), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G50), .B(G68), .Z(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G1698), .ZN(new_n246));
  AND2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT65), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT65), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI211_X1 g0055(.A(G226), .B(new_n246), .C1(new_n250), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT71), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G97), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n249), .B1(new_n247), .B2(new_n248), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n253), .A2(KEYINPUT65), .A3(new_n254), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n231), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n260), .B1(new_n263), .B2(G1698), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1698), .B1(new_n261), .B2(new_n262), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(KEYINPUT71), .A3(G226), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n258), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G1), .A2(G13), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(G33), .B2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n269), .A2(new_n273), .A3(KEYINPUT64), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT64), .ZN(new_n275));
  OAI211_X1 g0075(.A(G1), .B(G13), .C1(new_n252), .C2(new_n271), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(G238), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n276), .A2(G274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n273), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n270), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT13), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT13), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n270), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G200), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n286), .B1(new_n270), .B2(new_n283), .ZN(new_n290));
  AOI211_X1 g0090(.A(KEYINPUT13), .B(new_n282), .C1(new_n267), .C2(new_n269), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G190), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n208), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT67), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G77), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n297), .B1(new_n208), .B2(G68), .C1(new_n201), .C2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n268), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n300), .A2(KEYINPUT11), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(KEYINPUT11), .B1(new_n300), .B2(new_n302), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G68), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT12), .ZN(new_n307));
  INV_X1    g0107(.A(new_n305), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n302), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n203), .B1(new_n207), .B2(G20), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n303), .A2(new_n304), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n289), .A2(new_n293), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT14), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n288), .A2(KEYINPUT72), .A3(new_n316), .A4(G169), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(G169), .C1(new_n290), .C2(new_n291), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT72), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n292), .A2(G179), .ZN(new_n321));
  OAI21_X1  g0121(.A(G169), .B1(new_n290), .B2(new_n291), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT14), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n317), .A2(new_n320), .A3(new_n321), .A4(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n313), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n315), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n274), .A2(new_n278), .ZN(new_n327));
  INV_X1    g0127(.A(G226), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n281), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n265), .A2(G222), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n246), .B1(new_n261), .B2(new_n262), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G223), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n261), .A2(new_n262), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n330), .B(new_n332), .C1(new_n222), .C2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n329), .B1(new_n334), .B2(new_n269), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  OR3_X1    g0136(.A1(new_n335), .A2(KEYINPUT70), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n302), .ZN(new_n338));
  XOR2_X1   g0138(.A(KEYINPUT8), .B(G58), .Z(new_n339));
  INV_X1    g0139(.A(KEYINPUT66), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT8), .B(G58), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT66), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n296), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n298), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n338), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n207), .A2(G20), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n309), .A2(G50), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G50), .B2(new_n305), .ZN(new_n349));
  OR3_X1    g0149(.A1(new_n346), .A2(KEYINPUT9), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT9), .B1(new_n346), .B2(new_n349), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n350), .A2(new_n351), .B1(new_n335), .B2(G190), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT70), .B1(new_n335), .B2(new_n336), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n337), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT10), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT10), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n337), .A2(new_n352), .A3(new_n356), .A4(new_n353), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n342), .A2(new_n299), .B1(new_n208), .B2(new_n222), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n294), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n302), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n309), .A2(G77), .A3(new_n347), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n362), .B(new_n363), .C1(G77), .C2(new_n305), .ZN(new_n364));
  INV_X1    g0164(.A(new_n333), .ZN(new_n365));
  AOI22_X1  g0165(.A1(G107), .A2(new_n365), .B1(new_n263), .B2(new_n246), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n331), .A2(G238), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n269), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n281), .B1(new_n327), .B2(new_n223), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n364), .B1(new_n372), .B2(G200), .ZN(new_n373));
  INV_X1    g0173(.A(G190), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(new_n372), .ZN(new_n375));
  INV_X1    g0175(.A(G169), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G179), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n369), .A2(new_n378), .A3(new_n371), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n379), .A3(new_n364), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n335), .A2(new_n378), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n382), .A2(KEYINPUT69), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n346), .A2(new_n349), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n335), .B2(G169), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n385), .A2(KEYINPUT68), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(KEYINPUT68), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n382), .A2(KEYINPUT69), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n383), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n358), .A2(new_n381), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(KEYINPUT7), .A2(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n261), .A2(new_n262), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n254), .A2(new_n208), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT73), .B(G33), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n251), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n392), .B(G68), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(G58), .B(G68), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(G20), .B1(G159), .B2(new_n298), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g0200(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n208), .B(new_n253), .C1(new_n394), .C2(new_n251), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n403), .B2(KEYINPUT7), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n252), .A2(KEYINPUT73), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT73), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G33), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n248), .B1(new_n408), .B2(KEYINPUT3), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n396), .B1(new_n409), .B2(new_n208), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT16), .B(new_n399), .C1(new_n404), .C2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n402), .A2(new_n302), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n342), .B(new_n340), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n347), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT75), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n341), .A2(KEYINPUT75), .A3(new_n347), .A4(new_n343), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n417), .A2(new_n309), .ZN(new_n418));
  INV_X1    g0218(.A(new_n413), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n416), .A2(new_n418), .B1(new_n308), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n412), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n253), .B1(new_n394), .B2(new_n251), .ZN(new_n422));
  NOR2_X1   g0222(.A1(G223), .A2(G1698), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n328), .B2(G1698), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n422), .A2(new_n424), .B1(G33), .B2(G87), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT76), .B1(new_n425), .B2(new_n276), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G87), .ZN(new_n427));
  INV_X1    g0227(.A(new_n424), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n427), .B1(new_n409), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT76), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n269), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n276), .A2(G232), .A3(new_n277), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n281), .A2(new_n432), .A3(new_n378), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n426), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n425), .A2(new_n276), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n281), .A2(new_n432), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n376), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n421), .A2(new_n438), .A3(KEYINPUT18), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT77), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT77), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n421), .A2(new_n438), .A3(new_n441), .A4(KEYINPUT18), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n421), .A2(new_n438), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n440), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n436), .A2(G190), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(new_n426), .A3(new_n431), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n336), .B1(new_n435), .B2(new_n436), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n412), .A3(new_n420), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(KEYINPUT78), .A2(KEYINPUT17), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n450), .A2(new_n412), .A3(new_n420), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n446), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT79), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT79), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n446), .A2(new_n459), .A3(new_n456), .ZN(new_n460));
  AND4_X1   g0260(.A1(new_n326), .A2(new_n390), .A3(new_n458), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT88), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n305), .A2(G107), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n463), .B(KEYINPUT25), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n207), .A2(G33), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n338), .A2(new_n305), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT81), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n309), .A2(KEYINPUT81), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n464), .B1(new_n470), .B2(new_n224), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n251), .B1(new_n405), .B2(new_n407), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n208), .B(G87), .C1(new_n473), .C2(new_n248), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n218), .A2(KEYINPUT22), .A3(G20), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n474), .A2(KEYINPUT22), .B1(new_n333), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n394), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n208), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n224), .A2(G20), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT23), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n480), .B(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(KEYINPUT86), .B(new_n472), .C1(new_n476), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n302), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n474), .A2(KEYINPUT22), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n333), .A2(new_n475), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT86), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(new_n479), .A4(new_n482), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT86), .B1(new_n476), .B2(new_n483), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(KEYINPUT24), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n471), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(G250), .A2(G1698), .ZN(new_n495));
  INV_X1    g0295(.A(G257), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(G1698), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n422), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n408), .A2(G294), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n276), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g0300(.A(KEYINPUT5), .B(G41), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n272), .A2(G1), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(G264), .A3(new_n276), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n501), .A2(new_n276), .A3(G274), .A4(new_n502), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n500), .A2(new_n378), .A3(new_n506), .ZN(new_n507));
  OR2_X1    g0307(.A1(new_n500), .A2(KEYINPUT87), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n500), .A2(KEYINPUT87), .ZN(new_n509));
  INV_X1    g0309(.A(new_n506), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n507), .B1(new_n511), .B2(G169), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n462), .B1(new_n494), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n509), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n510), .B1(new_n500), .B2(KEYINPUT87), .ZN(new_n515));
  OAI21_X1  g0315(.A(G169), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n507), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n492), .A2(KEYINPUT24), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n485), .B1(new_n519), .B2(new_n491), .ZN(new_n520));
  OAI211_X1 g0320(.A(KEYINPUT88), .B(new_n518), .C1(new_n520), .C2(new_n471), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n500), .A2(new_n506), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n511), .A2(G190), .B1(G200), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n494), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n513), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n496), .A2(new_n246), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n225), .A2(G1698), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n526), .B(new_n527), .C1(new_n473), .C2(new_n248), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n261), .A2(new_n262), .A3(G303), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n276), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n269), .B1(new_n502), .B2(new_n501), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G270), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n505), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n301), .A2(new_n268), .B1(G20), .B2(new_n477), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G283), .ZN(new_n536));
  INV_X1    g0336(.A(G97), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n536), .B(new_n208), .C1(G33), .C2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n535), .A2(KEYINPUT20), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT20), .B1(new_n535), .B2(new_n538), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n308), .A2(new_n477), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n466), .B2(new_n477), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n534), .A2(KEYINPUT21), .A3(new_n545), .A4(G169), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  INV_X1    g0347(.A(new_n533), .ZN(new_n548));
  INV_X1    g0348(.A(new_n505), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n530), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(G169), .B1(new_n541), .B2(new_n543), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(G179), .A3(new_n545), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n546), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n534), .A2(G200), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n550), .A2(G190), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(new_n544), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT85), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n555), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT4), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n246), .A2(G244), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n563), .B1(new_n409), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n333), .A2(KEYINPUT4), .A3(G244), .A4(new_n246), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n333), .A2(G250), .A3(G1698), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n536), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n269), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n532), .A2(G257), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n505), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n376), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n571), .B1(new_n568), .B2(new_n269), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n378), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT6), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n537), .A2(new_n224), .ZN(new_n578));
  NOR2_X1   g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n224), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(G97), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT80), .ZN(new_n582));
  NAND2_X1  g0382(.A1(KEYINPUT6), .A2(G97), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n582), .B1(new_n583), .B2(G107), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n585), .A2(G20), .B1(G77), .B2(new_n298), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(new_n224), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n302), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n305), .A2(G97), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n470), .B2(new_n537), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n574), .A2(new_n576), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n280), .A2(new_n502), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n502), .A2(new_n219), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n276), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G238), .A2(G1698), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n223), .B2(G1698), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n478), .B1(new_n422), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n596), .B(new_n598), .C1(new_n601), .C2(new_n276), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(G179), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n376), .B2(new_n602), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT84), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n208), .B(G68), .C1(new_n473), .C2(new_n248), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n579), .A2(new_n218), .B1(new_n259), .B2(new_n208), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT19), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(G97), .ZN(new_n609));
  OAI22_X1  g0409(.A1(new_n607), .A2(new_n608), .B1(new_n294), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n302), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n360), .A2(new_n308), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(KEYINPUT82), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT82), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n338), .B1(new_n606), .B2(new_n610), .ZN(new_n616));
  INV_X1    g0416(.A(new_n613), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n360), .B(KEYINPUT83), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(new_n468), .A3(new_n469), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n605), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n621), .ZN(new_n623));
  AOI211_X1 g0423(.A(KEYINPUT84), .B(new_n623), .C1(new_n614), .C2(new_n618), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n604), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n575), .A2(G190), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n592), .B1(new_n302), .B2(new_n588), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n626), .B(new_n627), .C1(new_n336), .C2(new_n575), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT82), .B1(new_n612), .B2(new_n613), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n616), .A2(new_n615), .A3(new_n617), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n629), .A2(new_n630), .B1(new_n218), .B2(new_n470), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n602), .A2(G200), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n374), .B2(new_n602), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n595), .A2(new_n625), .A3(new_n628), .A4(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n461), .A2(new_n525), .A3(new_n562), .A4(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n389), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n445), .A2(new_n439), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n380), .A2(KEYINPUT89), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT89), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n377), .A2(new_n641), .A3(new_n379), .A4(new_n364), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n325), .A2(new_n324), .B1(new_n643), .B2(new_n314), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n453), .A2(new_n455), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n639), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n638), .B1(new_n646), .B2(new_n358), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n621), .B1(new_n629), .B2(new_n630), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT84), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n619), .A2(new_n605), .A3(new_n621), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n634), .B1(new_n651), .B2(new_n604), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n554), .B1(new_n494), .B2(new_n512), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n595), .A2(new_n628), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n652), .A2(new_n524), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n595), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT26), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n625), .A2(new_n656), .A3(new_n635), .A4(KEYINPUT26), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n625), .B(new_n655), .C1(new_n657), .C2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n461), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n647), .A2(new_n661), .ZN(G369));
  NAND3_X1  g0462(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n545), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n562), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n554), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G330), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n672), .B(KEYINPUT90), .Z(new_n673));
  NOR2_X1   g0473(.A1(new_n494), .A2(new_n512), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n668), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT92), .ZN(new_n676));
  INV_X1    g0476(.A(new_n668), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n494), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT91), .Z(new_n679));
  INV_X1    g0479(.A(new_n525), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n494), .A2(new_n512), .A3(new_n668), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n554), .A2(new_n668), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n683), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT93), .Z(G399));
  INV_X1    g0487(.A(new_n211), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G1), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n579), .A2(new_n218), .A3(new_n477), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n691), .A2(new_n692), .B1(new_n215), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  INV_X1    g0494(.A(G330), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n530), .A2(new_n548), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n598), .A2(new_n596), .ZN(new_n698));
  INV_X1    g0498(.A(new_n601), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n269), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n507), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n696), .B1(new_n701), .B2(new_n573), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT94), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n701), .A2(new_n573), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT30), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT94), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n706), .B(new_n696), .C1(new_n701), .C2(new_n573), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n700), .A2(new_n522), .A3(G179), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(new_n573), .A3(new_n534), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n703), .A2(new_n705), .A3(new_n707), .A4(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT31), .B1(new_n710), .B2(new_n668), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n705), .A2(new_n702), .A3(new_n709), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n668), .A2(KEYINPUT31), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n525), .A2(new_n636), .A3(new_n562), .A4(new_n677), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n695), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n660), .A2(new_n677), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n625), .A2(new_n656), .A3(new_n635), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT26), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(KEYINPUT95), .A3(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n513), .A2(new_n521), .A3(new_n554), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n652), .A2(new_n524), .A3(new_n654), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n722), .B(new_n625), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n720), .A2(new_n721), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT95), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n726), .A2(new_n727), .A3(new_n658), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT29), .B(new_n677), .C1(new_n725), .C2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n716), .B1(new_n719), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n694), .B1(new_n730), .B2(G1), .ZN(G364));
  INV_X1    g0531(.A(G13), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G45), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT96), .Z(new_n735));
  NAND3_X1  g0535(.A1(new_n690), .A2(G1), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT97), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT98), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n671), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(G20), .B1(KEYINPUT99), .B2(G169), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(KEYINPUT99), .B2(G169), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n268), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT100), .Z(new_n747));
  NOR2_X1   g0547(.A1(new_n208), .A2(new_n378), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n749), .A2(new_n374), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n749), .A2(new_n336), .A3(G190), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n202), .A2(new_n751), .B1(new_n753), .B2(new_n203), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n749), .A2(new_n374), .A3(new_n336), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G190), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n756), .A2(new_n201), .B1(new_n758), .B2(new_n222), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n374), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n208), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n537), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n208), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n757), .ZN(new_n765));
  INV_X1    g0565(.A(G159), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT32), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n763), .B(new_n769), .C1(G87), .C2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n764), .A2(new_n374), .A3(G200), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT101), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G107), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n365), .B1(new_n768), .B2(new_n767), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n760), .A2(new_n772), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n750), .A2(G322), .B1(new_n755), .B2(G326), .ZN(new_n778));
  INV_X1    g0578(.A(new_n758), .ZN(new_n779));
  INV_X1    g0579(.A(new_n765), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G311), .A2(new_n779), .B1(new_n780), .B2(G329), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G294), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n365), .B1(new_n783), .B2(new_n762), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G303), .B2(new_n771), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n774), .A2(G283), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT33), .B(G317), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT102), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(KEYINPUT102), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n789), .A2(new_n752), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n782), .A2(new_n785), .A3(new_n786), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n747), .B1(new_n777), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n747), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n741), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n365), .A2(new_n688), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n796), .A2(G355), .B1(new_n477), .B2(new_n688), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n688), .A2(new_n422), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n215), .A2(G45), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(new_n241), .C2(new_n272), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n793), .B1(new_n795), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n738), .B1(new_n743), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n672), .B(KEYINPUT90), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(G330), .B2(new_n671), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n803), .B1(new_n805), .B2(new_n738), .ZN(G396));
  NAND4_X1  g0606(.A1(new_n640), .A2(new_n364), .A3(new_n642), .A4(new_n668), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n364), .A2(new_n668), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n375), .A2(new_n380), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n660), .A2(new_n677), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n625), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n726), .B2(new_n658), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n668), .B1(new_n813), .B2(new_n655), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT106), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n807), .A2(KEYINPUT106), .A3(new_n809), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n811), .B1(new_n814), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n716), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT107), .Z(new_n822));
  AOI21_X1  g0622(.A(new_n737), .B1(new_n819), .B2(new_n820), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n747), .A2(new_n740), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT103), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n737), .B1(new_n826), .B2(G77), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT104), .B(G283), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n753), .A2(new_n828), .B1(new_n765), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G294), .B2(new_n750), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n774), .A2(G87), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n758), .A2(new_n477), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n333), .B(new_n833), .C1(G303), .C2(new_n755), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n763), .B1(G107), .B2(new_n771), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n831), .A2(new_n832), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n774), .A2(G68), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n201), .B2(new_n770), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT105), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n750), .A2(G143), .B1(new_n755), .B2(G137), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n752), .A2(G150), .B1(G159), .B2(new_n779), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n840), .A2(KEYINPUT34), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT34), .B1(new_n840), .B2(new_n841), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n422), .B1(new_n844), .B2(new_n765), .C1(new_n202), .C2(new_n762), .ZN(new_n845));
  OR3_X1    g0645(.A1(new_n842), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n836), .B1(new_n839), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n827), .B1(new_n847), .B2(new_n794), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n810), .B2(new_n740), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n824), .A2(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n733), .A2(new_n207), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT40), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n411), .A2(new_n302), .ZN(new_n853));
  INV_X1    g0653(.A(new_n401), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n409), .A2(new_n396), .A3(new_n208), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n403), .A2(KEYINPUT7), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(G68), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n854), .B1(new_n857), .B2(new_n399), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n420), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n666), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n457), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n859), .A2(new_n438), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n861), .A2(new_n864), .A3(new_n451), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT109), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n421), .B2(new_n860), .ZN(new_n868));
  AOI211_X1 g0668(.A(KEYINPUT109), .B(new_n666), .C1(new_n412), .C2(new_n420), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n451), .B(new_n443), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XOR2_X1   g0670(.A(KEYINPUT110), .B(KEYINPUT37), .Z(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n866), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n863), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(KEYINPUT38), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n861), .B1(new_n446), .B2(new_n456), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT111), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n443), .A2(new_n451), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n879), .B(new_n871), .C1(new_n869), .C2(new_n868), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n878), .B1(new_n880), .B2(new_n866), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT111), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n863), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n874), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n324), .A2(new_n325), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n325), .A2(new_n668), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n314), .A3(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n325), .B(new_n668), .C1(new_n324), .C2(new_n315), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n711), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n715), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n889), .A2(new_n810), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n852), .B1(new_n884), .B2(new_n893), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n868), .A2(new_n869), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(new_n879), .C1(KEYINPUT113), .C2(new_n871), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n456), .B2(new_n639), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT113), .B1(new_n868), .B2(new_n869), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n870), .A2(new_n872), .A3(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n878), .B(new_n896), .C1(new_n897), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n881), .A2(new_n863), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT40), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n894), .B1(new_n893), .B2(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT114), .Z(new_n905));
  NAND2_X1  g0705(.A1(new_n461), .A2(new_n892), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n695), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n905), .B2(new_n907), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n900), .A2(new_n901), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n884), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT112), .B1(new_n885), .B2(new_n668), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT112), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n324), .A2(new_n914), .A3(new_n325), .A4(new_n677), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n863), .A2(new_n873), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n878), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n875), .A2(KEYINPUT111), .A3(new_n876), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n882), .B1(new_n881), .B2(new_n863), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n380), .A2(new_n668), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n811), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(new_n889), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n445), .A2(new_n439), .A3(new_n666), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n917), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n719), .A2(new_n729), .A3(new_n461), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n647), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n928), .B(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n851), .B1(new_n909), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n931), .B2(new_n909), .ZN(new_n933));
  OAI21_X1  g0733(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n934), .A2(new_n215), .B1(G50), .B2(new_n203), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(G1), .A3(new_n732), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT108), .Z(new_n937));
  AOI211_X1 g0737(.A(new_n477), .B(new_n214), .C1(new_n585), .C2(KEYINPUT35), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(KEYINPUT35), .B2(new_n585), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT36), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n940), .B2(new_n939), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n933), .A2(new_n942), .ZN(G367));
  NAND2_X1  g0743(.A1(new_n681), .A2(new_n684), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n654), .B1(new_n627), .B2(new_n677), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n656), .A2(new_n668), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n944), .A2(KEYINPUT42), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n945), .B1(new_n513), .B2(new_n521), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n677), .B1(new_n950), .B2(new_n656), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT42), .B1(new_n944), .B2(new_n948), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n631), .A2(new_n668), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n652), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n625), .B2(new_n954), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT115), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n953), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(new_n953), .B2(new_n959), .ZN(new_n962));
  NOR4_X1   g0762(.A1(new_n961), .A2(new_n962), .A3(new_n682), .A4(new_n948), .ZN(new_n963));
  INV_X1    g0763(.A(new_n962), .ZN(new_n964));
  INV_X1    g0764(.A(new_n682), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n964), .A2(new_n960), .B1(new_n965), .B2(new_n947), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n689), .B(KEYINPUT41), .Z(new_n968));
  INV_X1    g0768(.A(KEYINPUT44), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n685), .A2(new_n969), .A3(new_n947), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n685), .B2(new_n947), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT116), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT116), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n973), .B(new_n969), .C1(new_n685), .C2(new_n947), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n685), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT45), .B1(new_n685), .B2(new_n947), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n965), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n681), .A2(new_n684), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n944), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n673), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n804), .A2(new_n944), .A3(new_n979), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n730), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n975), .A2(new_n976), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT116), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n986), .A2(new_n987), .A3(new_n682), .A4(new_n974), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n978), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n968), .B1(new_n989), .B2(new_n730), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n735), .A2(G1), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n967), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n795), .ZN(new_n993));
  INV_X1    g0793(.A(new_n798), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n994), .A2(new_n237), .B1(new_n211), .B2(new_n360), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n737), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n753), .A2(new_n766), .B1(new_n758), .B2(new_n201), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G143), .B2(new_n755), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n773), .A2(new_n222), .B1(new_n770), .B2(new_n202), .ZN(new_n999));
  INV_X1    g0799(.A(new_n762), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n999), .B1(G68), .B2(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n750), .A2(G150), .B1(G137), .B2(new_n780), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n998), .A2(new_n333), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n756), .A2(new_n829), .ZN(new_n1004));
  INV_X1    g0804(.A(G303), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n783), .A2(new_n753), .B1(new_n751), .B2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(G317), .C2(new_n780), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n773), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n422), .B1(G97), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n828), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1000), .A2(G107), .B1(new_n779), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1007), .B(new_n1009), .C1(KEYINPUT117), .C2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n771), .A2(G116), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT46), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1011), .A2(KEYINPUT117), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1003), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT47), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AND2_X1   g0819(.A1(new_n1019), .A2(new_n794), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n996), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n742), .B2(new_n956), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n992), .A2(new_n1023), .ZN(G387));
  NAND2_X1  g0824(.A1(new_n983), .A2(new_n991), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n750), .A2(G317), .B1(new_n755), .B2(G322), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n752), .A2(G311), .B1(G303), .B2(new_n779), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT48), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(KEYINPUT48), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1000), .A2(new_n1010), .B1(new_n771), .B2(G294), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n773), .A2(new_n477), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n422), .B(new_n1036), .C1(G326), .C2(new_n780), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G68), .A2(new_n779), .B1(new_n780), .B2(G150), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n756), .B2(new_n766), .C1(new_n201), .C2(new_n751), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n409), .B(new_n1040), .C1(G77), .C2(new_n771), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n774), .A2(G97), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n620), .A2(new_n1000), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n413), .A2(new_n752), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n747), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n234), .A2(new_n272), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1047), .A2(new_n798), .B1(new_n692), .B2(new_n796), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT50), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n339), .B2(new_n201), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n342), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n272), .B1(new_n203), .B2(new_n222), .ZN(new_n1052));
  NOR4_X1   g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n692), .A4(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1048), .A2(new_n1053), .B1(G107), .B2(new_n211), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n738), .B(new_n1046), .C1(new_n795), .C2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n681), .B2(new_n742), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n984), .A2(new_n689), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n983), .A2(new_n730), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1025), .B(new_n1056), .C1(new_n1057), .C2(new_n1058), .ZN(G393));
  NAND3_X1  g0859(.A1(new_n978), .A2(new_n988), .A3(new_n991), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n994), .A2(new_n244), .B1(new_n537), .B2(new_n211), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n737), .B1(new_n993), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n422), .B1(new_n203), .B2(new_n770), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n752), .A2(G50), .B1(G143), .B2(new_n780), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n342), .B2(new_n758), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(G77), .C2(new_n1000), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n750), .A2(G159), .B1(new_n755), .B2(G150), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G87), .B2(new_n774), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n750), .A2(G311), .B1(new_n755), .B2(G317), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT52), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G107), .B2(new_n774), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n365), .B1(new_n770), .B2(new_n828), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n752), .A2(G303), .B1(G322), .B2(new_n780), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n783), .B2(new_n758), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(G116), .C2(new_n1000), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1066), .A2(new_n1069), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1077), .A2(KEYINPUT118), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n747), .B1(new_n1077), .B2(KEYINPUT118), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1062), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n947), .B2(new_n742), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n989), .A2(new_n689), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n985), .B1(new_n978), .B2(new_n988), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1060), .B(new_n1081), .C1(new_n1082), .C2(new_n1083), .ZN(G390));
  AOI21_X1  g0884(.A(new_n916), .B1(new_n925), .B2(new_n889), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n889), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n677), .B(new_n810), .C1(new_n725), .C2(new_n728), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n924), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n916), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n902), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n912), .A2(new_n1085), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  AND4_X1   g0891(.A1(G330), .A2(new_n889), .A3(new_n810), .A4(new_n892), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n900), .A2(new_n901), .A3(new_n910), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n922), .B2(KEYINPUT39), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n923), .B1(new_n814), .B2(new_n810), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1089), .B1(new_n1096), .B2(new_n1086), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n916), .B1(new_n901), .B2(new_n900), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1087), .A2(new_n924), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n1086), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n716), .A2(new_n889), .A3(new_n810), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1093), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n461), .A2(G330), .A3(new_n892), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n929), .A2(new_n1105), .A3(new_n647), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n889), .B1(new_n716), .B2(new_n810), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n925), .B1(new_n1092), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n892), .A2(new_n818), .A3(G330), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1086), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1100), .A2(new_n1110), .A3(new_n1102), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1106), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1104), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1093), .A2(new_n1103), .A3(new_n1112), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n689), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1093), .A2(new_n1103), .A3(new_n991), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n758), .A2(new_n537), .B1(new_n765), .B2(new_n783), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n750), .A2(G116), .B1(new_n755), .B2(G283), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n224), .B2(new_n753), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1118), .B(new_n1120), .C1(G77), .C2(new_n1000), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n333), .B1(G87), .B2(new_n771), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT119), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n837), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n751), .A2(new_n844), .B1(new_n756), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1126), .A2(new_n365), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n780), .A2(G125), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  INV_X1    g0929(.A(G137), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1128), .B1(new_n758), .B2(new_n1129), .C1(new_n753), .C2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n771), .A2(G150), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT53), .Z(new_n1134));
  AOI22_X1  g0934(.A1(new_n1000), .A2(G159), .B1(new_n1008), .B2(G50), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1127), .A2(new_n1132), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n747), .B1(new_n1124), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n826), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n738), .B(new_n1137), .C1(new_n419), .C2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n912), .B2(new_n740), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1117), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1116), .A2(new_n1141), .ZN(G378));
  NAND2_X1  g0942(.A1(new_n358), .A2(new_n389), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n384), .A2(new_n860), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT124), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1143), .B(new_n1145), .ZN(new_n1146));
  XOR2_X1   g0946(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n740), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n737), .B1(G50), .B2(new_n825), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n409), .A2(new_n271), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1152), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n1153), .B(KEYINPUT120), .Z(new_n1154));
  OAI22_X1  g0954(.A1(new_n762), .A2(new_n203), .B1(new_n773), .B2(new_n202), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n750), .A2(G107), .B1(G283), .B2(new_n780), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n537), .B2(new_n753), .C1(new_n477), .C2(new_n756), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(new_n620), .C2(new_n779), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1152), .B1(G77), .B2(new_n771), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(KEYINPUT121), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1159), .A2(KEYINPUT121), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1158), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT58), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1154), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G125), .A2(new_n755), .B1(new_n1000), .B2(G150), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT123), .Z(new_n1166));
  AOI22_X1  g0966(.A1(new_n752), .A2(G132), .B1(G137), .B2(new_n779), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1125), .B2(new_n751), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT122), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n770), .A2(new_n1129), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1166), .B(new_n1171), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(KEYINPUT59), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1008), .A2(G159), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G33), .B(G41), .C1(new_n780), .C2(G124), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1164), .B1(new_n1163), .B2(new_n1162), .C1(new_n1173), .C2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1151), .B1(new_n1178), .B2(new_n794), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1150), .A2(new_n1179), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n889), .A2(new_n810), .A3(new_n892), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT40), .B1(new_n1181), .B2(new_n922), .ZN(new_n1182));
  OAI21_X1  g0982(.A(G330), .B1(new_n903), .B2(new_n893), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1147), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1146), .B(new_n1184), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n852), .B1(new_n900), .B2(new_n901), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n695), .B1(new_n1181), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1148), .B1(new_n1188), .B2(new_n894), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n928), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1185), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n894), .A3(new_n1148), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n926), .A2(new_n927), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n917), .A4(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1190), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1180), .B1(new_n1195), .B2(new_n991), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1106), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1115), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1190), .A2(KEYINPUT57), .A3(new_n1194), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n689), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1115), .A2(new_n1197), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1196), .B1(new_n1200), .B2(new_n1202), .ZN(G375));
  INV_X1    g1003(.A(new_n968), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1108), .A2(new_n1111), .A3(new_n1106), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1113), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1086), .A2(new_n1149), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n753), .A2(new_n477), .B1(new_n756), .B2(new_n783), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n333), .B(new_n1209), .C1(G97), .C2(new_n771), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n774), .A2(G77), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n750), .A2(G283), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1005), .B2(new_n765), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G107), .B2(new_n779), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1210), .A2(new_n1043), .A3(new_n1211), .A4(new_n1214), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n751), .A2(new_n1130), .B1(new_n756), .B2(new_n844), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G150), .B2(new_n779), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n422), .B1(new_n202), .B2(new_n773), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT125), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n753), .A2(new_n1129), .B1(new_n765), .B2(new_n1125), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G50), .B2(new_n1000), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n771), .A2(G159), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1217), .A2(new_n1219), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n747), .B1(new_n1215), .B2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n738), .B(new_n1224), .C1(new_n203), .C2(new_n1138), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1207), .A2(new_n991), .B1(new_n1208), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1206), .A2(new_n1226), .ZN(G381));
  OR2_X1    g1027(.A1(G393), .A2(G396), .ZN(new_n1228));
  OR4_X1    g1028(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1228), .ZN(new_n1229));
  OR4_X1    g1029(.A1(G387), .A2(new_n1229), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1030(.A(G378), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n667), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G407), .B(G213), .C1(G375), .C2(new_n1232), .ZN(G409));
  XOR2_X1   g1033(.A(G393), .B(G396), .Z(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n992), .A2(new_n1023), .A3(G390), .ZN(new_n1236));
  AOI21_X1  g1036(.A(G390), .B1(new_n992), .B2(new_n1023), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G390), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(G387), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n992), .A2(new_n1023), .A3(G390), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1234), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1238), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(G213), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(G343), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1190), .A2(new_n1204), .A3(new_n1194), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1198), .B2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1195), .A2(KEYINPUT126), .A3(new_n1201), .A4(new_n1204), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1196), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1231), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G378), .B(new_n1196), .C1(new_n1200), .C2(new_n1202), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1245), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT60), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1205), .B1(new_n1112), .B2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1108), .A2(new_n1111), .A3(new_n1106), .A4(KEYINPUT60), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n689), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1226), .ZN(new_n1258));
  INV_X1    g1058(.A(G384), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT62), .B1(new_n1253), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT127), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1245), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  AOI211_X1 g1069(.A(KEYINPUT127), .B(new_n1245), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1264), .A2(KEYINPUT62), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1265), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1245), .A2(G2897), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1263), .B(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1243), .B1(new_n1273), .B2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1271), .A2(KEYINPUT63), .A3(new_n1264), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1253), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(new_n1263), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1243), .A2(KEYINPUT61), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1275), .A2(new_n1282), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1280), .A2(new_n1283), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1279), .A2(new_n1286), .ZN(G405));
  NAND2_X1  g1087(.A1(G375), .A2(new_n1231), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1252), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1289), .B(new_n1264), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1243), .ZN(G402));
endmodule


