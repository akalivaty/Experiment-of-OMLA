//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n449, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n459), .A2(new_n461), .A3(G125), .ZN(new_n462));
  AND2_X1   g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(new_n460), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(KEYINPUT3), .A3(new_n467), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n471), .A2(G137), .A3(new_n472), .A4(new_n459), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n471), .A2(new_n459), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(new_n472), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(new_n459), .A2(new_n461), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n486), .A2(new_n472), .A3(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n472), .A2(G138), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n471), .A2(new_n459), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n488), .B1(new_n490), .B2(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n471), .A2(G126), .A3(G2105), .A4(new_n459), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G114), .C2(new_n472), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n491), .A2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(KEYINPUT6), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT69), .B(KEYINPUT6), .ZN(new_n500));
  OAI211_X1 g075(.A(G50), .B(new_n499), .C1(new_n500), .C2(new_n498), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n506));
  OAI21_X1  g081(.A(G651), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n507), .A2(new_n508), .A3(G50), .A4(new_n499), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n498), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n514), .A2(new_n515), .B1(new_n505), .B2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n514), .A2(new_n515), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n517), .A2(G88), .B1(new_n521), .B2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n510), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  OR2_X1    g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n507), .A2(new_n499), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  OAI221_X1 g108(.A(new_n528), .B1(new_n530), .B2(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n517), .A2(G89), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n517), .A2(G90), .ZN(new_n538));
  INV_X1    g113(.A(new_n499), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n513), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n519), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n538), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n547), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(G171));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  INV_X1    g126(.A(G68), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n519), .A2(new_n551), .B1(new_n552), .B2(new_n497), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI221_X1 g130(.A(KEYINPUT72), .B1(new_n552), .B2(new_n497), .C1(new_n519), .C2(new_n551), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n555), .A2(G651), .A3(new_n556), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(KEYINPUT73), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(KEYINPUT73), .ZN(new_n559));
  AOI22_X1  g134(.A1(G81), .A2(new_n517), .B1(new_n540), .B2(G43), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n563));
  XOR2_X1   g138(.A(new_n563), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  AOI22_X1  g142(.A1(new_n525), .A2(new_n526), .B1(KEYINPUT6), .B2(new_n498), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n507), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  OR3_X1    g145(.A1(new_n569), .A2(KEYINPUT77), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT77), .B1(new_n569), .B2(new_n570), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n519), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n571), .A2(new_n572), .B1(G651), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI211_X1 g152(.A(KEYINPUT75), .B(KEYINPUT9), .C1(new_n532), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n540), .A2(G53), .A3(new_n579), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n578), .A2(KEYINPUT76), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT76), .B1(new_n578), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n576), .B1(new_n581), .B2(new_n582), .ZN(G299));
  AND2_X1   g158(.A1(new_n548), .A2(new_n549), .ZN(G301));
  NAND3_X1  g159(.A1(new_n507), .A2(new_n568), .A3(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n586));
  OAI211_X1 g161(.A(G49), .B(new_n499), .C1(new_n500), .C2(new_n498), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n519), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n507), .A2(new_n568), .A3(G86), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n507), .A2(G48), .A3(new_n499), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n517), .A2(G85), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  XNOR2_X1  g172(.A(KEYINPUT78), .B(G47), .ZN(new_n598));
  OAI221_X1 g173(.A(new_n596), .B1(new_n498), .B2(new_n597), .C1(new_n532), .C2(new_n598), .ZN(G290));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(G301), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n517), .A2(G92), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT10), .Z(new_n603));
  AOI22_X1  g178(.A1(new_n527), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(new_n498), .ZN(new_n605));
  INV_X1    g180(.A(G54), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n606), .B1(new_n532), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n540), .A2(KEYINPUT79), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(KEYINPUT80), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n603), .A2(new_n610), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n601), .B1(new_n616), .B2(new_n600), .ZN(G284));
  AOI21_X1  g192(.A(new_n601), .B1(new_n616), .B2(new_n600), .ZN(G321));
  NAND2_X1  g193(.A1(G299), .A2(new_n600), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n600), .B2(G168), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(new_n600), .B2(G168), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n616), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND3_X1  g198(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n616), .A2(new_n622), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT81), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n625), .B1(new_n627), .B2(G868), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g204(.A1(new_n468), .A2(new_n459), .A3(new_n461), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT82), .B(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n477), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n479), .A2(G123), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n638));
  INV_X1    g213(.A(G111), .ZN(new_n639));
  AOI22_X1  g214(.A1(new_n637), .A2(new_n638), .B1(new_n639), .B2(G2105), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n638), .B2(new_n637), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n635), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n642), .A2(G2096), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(G2096), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n634), .A2(new_n643), .A3(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT86), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT85), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT15), .B(G2435), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2438), .ZN(new_n655));
  XOR2_X1   g230(.A(G2427), .B(G2430), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT84), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n653), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(KEYINPUT88), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(new_n669), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n673));
  OAI221_X1 g248(.A(new_n666), .B1(new_n668), .B2(new_n669), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n666), .A2(new_n667), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n683), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n683), .B2(new_n689), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G229));
  MUX2_X1   g273(.A(G21), .B(G286), .S(G16), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT100), .ZN(new_n700));
  INV_X1    g275(.A(G1966), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  MUX2_X1   g278(.A(G5), .B(G301), .S(G16), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G1961), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT27), .B(G1996), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G29), .A2(G32), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n479), .A2(G129), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT98), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n477), .A2(G141), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT26), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G105), .B2(new_n468), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n711), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT99), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n709), .B1(new_n717), .B2(G29), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n702), .B(new_n706), .C1(new_n708), .C2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G33), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n477), .A2(G139), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n723));
  NAND3_X1  g298(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT97), .ZN(new_n727));
  NAND2_X1  g302(.A1(G115), .A2(G2104), .ZN(new_n728));
  INV_X1    g303(.A(G127), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n485), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n727), .B1(G2105), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n721), .B1(new_n731), .B2(new_n720), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2072), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n720), .A2(G35), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G162), .B2(new_n720), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT29), .B(G2090), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G34), .ZN(new_n738));
  AOI21_X1  g313(.A(G29), .B1(new_n738), .B2(KEYINPUT24), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(KEYINPUT24), .B2(new_n738), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n474), .B2(new_n720), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT30), .B(G28), .ZN(new_n745));
  OR2_X1    g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  NAND2_X1  g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n745), .A2(new_n720), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n642), .B2(new_n720), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n737), .A2(new_n743), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n477), .A2(G140), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n479), .A2(G128), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n472), .A2(G116), .ZN(new_n754));
  OAI21_X1  g329(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n752), .B(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n720), .A2(G26), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT28), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2067), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n704), .A2(G1961), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n733), .A2(new_n751), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n616), .ZN(new_n764));
  MUX2_X1   g339(.A(G4), .B(new_n764), .S(G16), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G1348), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n720), .A2(G27), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G164), .B2(new_n720), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT102), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT101), .B(G2078), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n719), .A2(new_n763), .A3(new_n766), .A4(new_n771), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT90), .B(G16), .Z(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(G19), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n561), .B2(new_n774), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT95), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G1341), .Z(new_n778));
  OR2_X1    g353(.A1(new_n718), .A2(new_n708), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n765), .A2(G1348), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n773), .A2(G20), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT23), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1956), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n778), .A2(new_n779), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n772), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G6), .B(G305), .S(G16), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT91), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT32), .B(G1981), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT92), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n789), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n774), .A2(G22), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n774), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT93), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n587), .A2(new_n586), .ZN(new_n798));
  INV_X1    g373(.A(G87), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n513), .A2(new_n516), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n797), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n585), .A2(KEYINPUT93), .A3(new_n586), .A4(new_n587), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  MUX2_X1   g378(.A(G23), .B(new_n803), .S(G16), .Z(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT33), .B(G1976), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n792), .A2(new_n796), .A3(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT94), .Z(new_n808));
  INV_X1    g383(.A(KEYINPUT34), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n720), .A2(G25), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n477), .A2(G131), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n479), .A2(G119), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n472), .A2(G107), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n812), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT89), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n811), .B1(new_n817), .B2(new_n720), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G1991), .Z(new_n819));
  XOR2_X1   g394(.A(new_n818), .B(new_n819), .Z(new_n820));
  MUX2_X1   g395(.A(G24), .B(G290), .S(new_n774), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1986), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n808), .B2(new_n809), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n810), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT36), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n810), .A2(new_n827), .A3(new_n824), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n787), .B1(new_n826), .B2(new_n828), .ZN(G311));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(new_n786), .ZN(G150));
  AOI22_X1  g406(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(new_n498), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT103), .B(G93), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n517), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n540), .A2(G55), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n616), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n624), .A2(new_n837), .ZN(new_n842));
  INV_X1    g417(.A(new_n837), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n559), .A2(new_n560), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n844), .B2(new_n558), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n841), .B(new_n846), .Z(new_n847));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(G860), .B1(new_n847), .B2(new_n848), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n849), .A2(KEYINPUT104), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(KEYINPUT104), .B1(new_n849), .B2(new_n850), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n839), .B1(new_n851), .B2(new_n852), .ZN(G145));
  NOR2_X1   g428(.A1(new_n731), .A2(new_n716), .ZN(new_n854));
  INV_X1    g429(.A(new_n717), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(new_n731), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n477), .A2(G142), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n479), .A2(G130), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n472), .A2(G118), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n631), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n816), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(G164), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n756), .B(KEYINPUT105), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(G164), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n856), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n864), .A2(new_n866), .ZN(new_n871));
  INV_X1    g446(.A(new_n865), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n856), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n642), .B(new_n474), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n483), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  INV_X1    g455(.A(new_n878), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n870), .A2(new_n875), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  AND2_X1   g459(.A1(new_n627), .A2(new_n846), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n627), .A2(new_n846), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n611), .A2(G299), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n611), .A2(G299), .A3(KEYINPUT106), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT107), .B1(new_n611), .B2(G299), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n581), .A2(new_n582), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n894), .A2(new_n613), .A3(new_n895), .A4(new_n576), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT41), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n897), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n890), .A2(new_n891), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n887), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n900), .B(new_n899), .C1(new_n885), .C2(new_n886), .ZN(new_n905));
  XNOR2_X1  g480(.A(G305), .B(KEYINPUT108), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(G166), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n803), .B(G290), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT109), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(KEYINPUT42), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n911), .B(new_n912), .Z(new_n913));
  AND3_X1   g488(.A1(new_n904), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n904), .B2(new_n905), .ZN(new_n915));
  OAI21_X1  g490(.A(G868), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(G868), .B2(new_n843), .ZN(G295));
  OAI21_X1  g492(.A(new_n916), .B1(G868), .B2(new_n843), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT111), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n548), .A2(KEYINPUT110), .A3(new_n549), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT110), .B1(new_n548), .B2(new_n549), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n845), .B2(new_n842), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n561), .A2(new_n843), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n624), .A2(new_n837), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n928), .B(new_n929), .C1(new_n924), .C2(new_n925), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(G286), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n899), .A2(new_n900), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n927), .A2(new_n930), .A3(G168), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n927), .A2(new_n930), .A3(G168), .ZN(new_n936));
  AOI21_X1  g511(.A(G168), .B1(new_n927), .B2(new_n930), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n935), .B1(new_n903), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n909), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n909), .B(new_n935), .C1(new_n903), .C2(new_n938), .ZN(new_n942));
  AND4_X1   g517(.A1(new_n923), .A2(new_n941), .A3(new_n880), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n939), .B2(new_n940), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n923), .B1(new_n944), .B2(new_n942), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n921), .B(new_n922), .C1(new_n943), .C2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n941), .A2(new_n880), .A3(new_n942), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n923), .A3(new_n942), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n919), .A4(new_n920), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n946), .A2(new_n950), .ZN(G397));
  NAND3_X1  g526(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT113), .ZN(new_n953));
  NAND2_X1  g528(.A1(G303), .A2(G8), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n957));
  NAND4_X1  g532(.A1(G303), .A2(new_n957), .A3(KEYINPUT55), .A4(G8), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n953), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n961));
  INV_X1    g536(.A(new_n488), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n492), .A2(new_n494), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n464), .A2(G40), .A3(new_n473), .A4(new_n469), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n491), .B2(new_n495), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT115), .B1(new_n967), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G2090), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n966), .B1(new_n491), .B2(new_n495), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT50), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n976), .A2(new_n977), .A3(new_n969), .A4(new_n971), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n973), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n968), .B1(new_n975), .B2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(KEYINPUT45), .B(new_n966), .C1(new_n491), .C2(new_n495), .ZN(new_n982));
  AOI21_X1  g557(.A(G1971), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n959), .B1(new_n985), .B2(G8), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n967), .A2(new_n972), .A3(G2090), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n959), .B(G8), .C1(new_n983), .C2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G8), .ZN(new_n989));
  AOI21_X1  g564(.A(G1384), .B1(new_n963), .B2(new_n964), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n990), .B2(new_n969), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n801), .A2(G1976), .A3(new_n802), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT114), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n801), .A2(new_n994), .A3(G1976), .A4(new_n802), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(G288), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n991), .A2(new_n993), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT49), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n540), .A2(G48), .B1(new_n591), .B2(G651), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(new_n593), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G305), .A2(G1981), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1000), .A3(new_n593), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G305), .A2(G1981), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(KEYINPUT49), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n1007), .A3(new_n991), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n998), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n991), .A2(new_n993), .A3(new_n995), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT52), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n988), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT122), .B1(new_n986), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n959), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n969), .B(new_n971), .C1(new_n990), .C2(new_n960), .ZN(new_n1015));
  AOI21_X1  g590(.A(G2090), .B1(new_n1015), .B2(KEYINPUT115), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n983), .B1(new_n1016), .B2(new_n978), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n1017), .B2(new_n989), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT122), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1011), .A2(new_n998), .A3(new_n1008), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1018), .A2(new_n1019), .A3(new_n988), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1013), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n975), .A2(new_n980), .ZN(new_n1023));
  INV_X1    g598(.A(G2078), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n969), .A4(new_n982), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n980), .A2(G1384), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n968), .B1(new_n965), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n975), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1029), .A2(KEYINPUT53), .A3(new_n1024), .A4(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT120), .B(G1961), .Z(new_n1033));
  NAND2_X1  g608(.A1(new_n1015), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1027), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1035), .A2(new_n1036), .A3(G171), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n1035), .B2(G171), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1022), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT45), .B1(new_n965), .B2(new_n966), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1028), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n969), .B1(G164), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n701), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n976), .A2(new_n742), .A3(new_n969), .A4(new_n971), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1044), .A2(KEYINPUT117), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT117), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G286), .A2(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1051), .B(G8), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1049), .B(KEYINPUT119), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n967), .A2(new_n972), .A3(G2084), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1966), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1044), .A2(KEYINPUT117), .A3(new_n1045), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n989), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(new_n1051), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT51), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1065), .A3(new_n1049), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1050), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1040), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1050), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1053), .B1(new_n1061), .B2(new_n1051), .ZN(new_n1071));
  OAI21_X1  g646(.A(G8), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT118), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1065), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1066), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1068), .B(new_n1070), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT124), .B1(new_n1069), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1035), .A2(G171), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT121), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1035), .A2(new_n1036), .A3(G171), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1023), .A2(new_n969), .A3(new_n982), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(KEYINPUT53), .A3(new_n1024), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1083), .A2(G301), .A3(new_n1027), .A4(new_n1034), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1027), .A3(new_n1034), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G171), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1089), .B(KEYINPUT54), .C1(G171), .C2(new_n1035), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1087), .A2(new_n1013), .A3(new_n1021), .A4(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT123), .B1(new_n1067), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1013), .A2(new_n1021), .A3(new_n1090), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT54), .B1(new_n1039), .B2(new_n1084), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1070), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT56), .B(G2072), .ZN(new_n1099));
  INV_X1    g674(.A(G1956), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1082), .A2(new_n1099), .B1(new_n1015), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(new_n578), .B2(new_n580), .ZN(new_n1102));
  AOI22_X1  g677(.A1(G299), .A2(KEYINPUT57), .B1(new_n576), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1015), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n990), .A2(new_n969), .ZN(new_n1106));
  OAI22_X1  g681(.A1(new_n1105), .A2(G1348), .B1(G2067), .B2(new_n1106), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n616), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1104), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1996), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT58), .B(G1341), .Z(new_n1112));
  AOI22_X1  g687(.A1(new_n1082), .A2(new_n1111), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(new_n624), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1114), .B(KEYINPUT59), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n1104), .A2(KEYINPUT61), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1104), .A2(KEYINPUT61), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1107), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT116), .B1(new_n612), .B2(new_n615), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n764), .A2(KEYINPUT116), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1122), .A2(new_n1123), .B1(new_n1119), .B2(new_n1107), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1110), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1092), .A2(new_n1098), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1020), .ZN(new_n1127));
  INV_X1    g702(.A(new_n991), .ZN(new_n1128));
  NOR2_X1   g703(.A1(G288), .A2(G1976), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1003), .B1(new_n1008), .B2(new_n1129), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1127), .A2(new_n988), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1012), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1018), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1064), .A2(G286), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1135), .A2(new_n1132), .ZN(new_n1137));
  INV_X1    g712(.A(new_n987), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n989), .B1(new_n1138), .B2(new_n984), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1137), .B(new_n1133), .C1(new_n959), .C2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1131), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1096), .A2(KEYINPUT62), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(new_n1076), .A4(new_n1040), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1078), .A2(new_n1126), .A3(new_n1141), .A4(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1023), .A2(new_n968), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n717), .A2(new_n1111), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n756), .B(G2067), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n716), .B2(G1996), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n816), .B(new_n819), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(G290), .B(G1986), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1146), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1145), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n817), .A2(new_n819), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT125), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1155), .A2(new_n1157), .B1(G2067), .B2(new_n756), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1151), .A2(new_n1146), .ZN(new_n1159));
  NOR2_X1   g734(.A1(G290), .A2(G1986), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1146), .A2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT48), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1158), .A2(new_n1146), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1146), .A2(new_n1111), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT46), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1146), .B1(new_n1148), .B2(new_n716), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT47), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT126), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n1154), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g746(.A(G401), .ZN(new_n1173));
  NAND3_X1  g747(.A1(new_n1173), .A2(G319), .A3(new_n680), .ZN(new_n1174));
  NOR2_X1   g748(.A1(G229), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g749(.A(new_n883), .B(new_n1175), .C1(new_n945), .C2(new_n943), .ZN(G225));
  INV_X1    g750(.A(G225), .ZN(G308));
endmodule


