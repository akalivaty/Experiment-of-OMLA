

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U322 ( .A(n348), .B(n347), .Z(n552) );
  XOR2_X1 U323 ( .A(n342), .B(n341), .Z(n290) );
  XNOR2_X1 U324 ( .A(n331), .B(KEYINPUT107), .ZN(n332) );
  XNOR2_X1 U325 ( .A(n333), .B(n332), .ZN(n364) );
  AND2_X1 U326 ( .A1(n364), .A2(n363), .ZN(n365) );
  XNOR2_X1 U327 ( .A(n297), .B(KEYINPUT32), .ZN(n298) );
  INV_X1 U328 ( .A(KEYINPUT110), .ZN(n373) );
  XNOR2_X1 U329 ( .A(n335), .B(n298), .ZN(n300) );
  XNOR2_X1 U330 ( .A(n373), .B(KEYINPUT48), .ZN(n374) );
  XNOR2_X1 U331 ( .A(n375), .B(n374), .ZN(n541) );
  XNOR2_X1 U332 ( .A(G8GAT), .B(G183GAT), .ZN(n336) );
  NOR2_X1 U333 ( .A1(n412), .A2(n511), .ZN(n568) );
  XNOR2_X1 U334 ( .A(n445), .B(G176GAT), .ZN(n446) );
  XNOR2_X1 U335 ( .A(n447), .B(n446), .ZN(G1349GAT) );
  INV_X1 U336 ( .A(KEYINPUT13), .ZN(n291) );
  NAND2_X1 U337 ( .A1(n291), .A2(G57GAT), .ZN(n294) );
  INV_X1 U338 ( .A(G57GAT), .ZN(n292) );
  NAND2_X1 U339 ( .A1(n292), .A2(KEYINPUT13), .ZN(n293) );
  NAND2_X1 U340 ( .A1(n294), .A2(n293), .ZN(n296) );
  XNOR2_X1 U341 ( .A(G71GAT), .B(G78GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n335) );
  AND2_X1 U343 ( .A1(G230GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U344 ( .A(G176GAT), .B(G92GAT), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n299), .B(G64GAT), .ZN(n383) );
  XOR2_X1 U346 ( .A(n300), .B(n383), .Z(n303) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n301), .B(KEYINPUT71), .ZN(n349) );
  XNOR2_X1 U349 ( .A(G120GAT), .B(n349), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n303), .B(n302), .ZN(n312) );
  XOR2_X1 U351 ( .A(G204GAT), .B(G106GAT), .Z(n305) );
  XNOR2_X1 U352 ( .A(KEYINPUT70), .B(G148GAT), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U354 ( .A(KEYINPUT69), .B(n306), .Z(n427) );
  INV_X1 U355 ( .A(n427), .ZN(n310) );
  XOR2_X1 U356 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n308) );
  XNOR2_X1 U357 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U359 ( .A(n310), .B(n309), .Z(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n367) );
  XOR2_X1 U361 ( .A(n367), .B(KEYINPUT41), .Z(n498) );
  XOR2_X1 U362 ( .A(G29GAT), .B(G36GAT), .Z(n314) );
  XNOR2_X1 U363 ( .A(G50GAT), .B(G43GAT), .ZN(n313) );
  XNOR2_X1 U364 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U365 ( .A(KEYINPUT7), .B(KEYINPUT67), .Z(n316) );
  XNOR2_X1 U366 ( .A(KEYINPUT66), .B(KEYINPUT8), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n362) );
  XOR2_X1 U369 ( .A(G113GAT), .B(G197GAT), .Z(n320) );
  XNOR2_X1 U370 ( .A(G169GAT), .B(G141GAT), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U372 ( .A(KEYINPUT64), .B(KEYINPUT30), .Z(n322) );
  XNOR2_X1 U373 ( .A(KEYINPUT29), .B(KEYINPUT65), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n329) );
  XNOR2_X1 U376 ( .A(G22GAT), .B(G15GAT), .ZN(n325) );
  XOR2_X1 U377 ( .A(n325), .B(G1GAT), .Z(n334) );
  XNOR2_X1 U378 ( .A(n334), .B(G8GAT), .ZN(n327) );
  NAND2_X1 U379 ( .A1(G229GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U382 ( .A(n362), .B(n330), .Z(n569) );
  OR2_X1 U383 ( .A1(n569), .A2(n498), .ZN(n333) );
  XOR2_X1 U384 ( .A(KEYINPUT46), .B(KEYINPUT108), .Z(n331) );
  XNOR2_X1 U385 ( .A(n335), .B(n334), .ZN(n348) );
  XOR2_X1 U386 ( .A(n336), .B(G211GAT), .Z(n380) );
  XNOR2_X1 U387 ( .A(n380), .B(KEYINPUT79), .ZN(n338) );
  XOR2_X1 U388 ( .A(G127GAT), .B(G155GAT), .Z(n395) );
  XNOR2_X1 U389 ( .A(n395), .B(G64GAT), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U391 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n340) );
  NAND2_X1 U392 ( .A1(G231GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U394 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n344) );
  XNOR2_X1 U395 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U397 ( .A(n345), .B(KEYINPUT78), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n290), .B(n346), .ZN(n347) );
  XOR2_X1 U399 ( .A(KEYINPUT106), .B(n552), .Z(n557) );
  XOR2_X1 U400 ( .A(KEYINPUT10), .B(n349), .Z(n351) );
  NAND2_X1 U401 ( .A1(G232GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U403 ( .A(G92GAT), .B(G162GAT), .Z(n353) );
  XNOR2_X1 U404 ( .A(G134GAT), .B(G106GAT), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U406 ( .A(n355), .B(n354), .ZN(n360) );
  XOR2_X1 U407 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n357) );
  XNOR2_X1 U408 ( .A(G190GAT), .B(KEYINPUT74), .ZN(n356) );
  XNOR2_X1 U409 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U410 ( .A(G218GAT), .B(n358), .Z(n359) );
  XNOR2_X1 U411 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U412 ( .A(n362), .B(n361), .ZN(n554) );
  INV_X1 U413 ( .A(n554), .ZN(n562) );
  AND2_X1 U414 ( .A1(n557), .A2(n562), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n365), .B(KEYINPUT47), .ZN(n372) );
  XOR2_X1 U416 ( .A(KEYINPUT36), .B(n554), .Z(n582) );
  INV_X1 U417 ( .A(n552), .ZN(n575) );
  NOR2_X1 U418 ( .A1(n582), .A2(n575), .ZN(n366) );
  XNOR2_X1 U419 ( .A(KEYINPUT45), .B(n366), .ZN(n368) );
  NAND2_X1 U420 ( .A1(n368), .A2(n367), .ZN(n369) );
  XNOR2_X1 U421 ( .A(KEYINPUT109), .B(n369), .ZN(n370) );
  INV_X1 U422 ( .A(n569), .ZN(n544) );
  XOR2_X1 U423 ( .A(KEYINPUT68), .B(n544), .Z(n452) );
  NAND2_X1 U424 ( .A1(n370), .A2(n452), .ZN(n371) );
  NAND2_X1 U425 ( .A1(n372), .A2(n371), .ZN(n375) );
  XNOR2_X1 U426 ( .A(KEYINPUT82), .B(KEYINPUT18), .ZN(n376) );
  XNOR2_X1 U427 ( .A(n376), .B(KEYINPUT19), .ZN(n377) );
  XOR2_X1 U428 ( .A(n377), .B(KEYINPUT17), .Z(n379) );
  XNOR2_X1 U429 ( .A(G169GAT), .B(G190GAT), .ZN(n378) );
  XNOR2_X1 U430 ( .A(n379), .B(n378), .ZN(n441) );
  XNOR2_X1 U431 ( .A(n441), .B(n380), .ZN(n390) );
  XOR2_X1 U432 ( .A(G204GAT), .B(KEYINPUT89), .Z(n382) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U435 ( .A(n384), .B(n383), .Z(n388) );
  XOR2_X1 U436 ( .A(KEYINPUT83), .B(KEYINPUT21), .Z(n386) );
  XNOR2_X1 U437 ( .A(G197GAT), .B(G218GAT), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n386), .B(n385), .ZN(n417) );
  XNOR2_X1 U439 ( .A(G36GAT), .B(n417), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U441 ( .A(n390), .B(n389), .Z(n514) );
  INV_X1 U442 ( .A(n514), .ZN(n455) );
  NOR2_X1 U443 ( .A1(n541), .A2(n455), .ZN(n391) );
  XOR2_X1 U444 ( .A(KEYINPUT54), .B(n391), .Z(n412) );
  XOR2_X1 U445 ( .A(G57GAT), .B(G85GAT), .Z(n393) );
  XNOR2_X1 U446 ( .A(G29GAT), .B(G148GAT), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U448 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U449 ( .A1(G225GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n397), .B(n396), .ZN(n411) );
  XOR2_X1 U451 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n399) );
  XNOR2_X1 U452 ( .A(G1GAT), .B(KEYINPUT87), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U454 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n401) );
  XNOR2_X1 U455 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U457 ( .A(n403), .B(n402), .Z(n409) );
  XOR2_X1 U458 ( .A(G120GAT), .B(KEYINPUT0), .Z(n405) );
  XNOR2_X1 U459 ( .A(G113GAT), .B(G134GAT), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n431) );
  XOR2_X1 U461 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n407) );
  XNOR2_X1 U462 ( .A(G141GAT), .B(G162GAT), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n418) );
  XNOR2_X1 U464 ( .A(n431), .B(n418), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n467) );
  INV_X1 U467 ( .A(n467), .ZN(n511) );
  XOR2_X1 U468 ( .A(KEYINPUT84), .B(KEYINPUT22), .Z(n414) );
  XNOR2_X1 U469 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U471 ( .A(G50GAT), .B(G22GAT), .Z(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n424) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U474 ( .A(G78GAT), .B(G155GAT), .Z(n420) );
  XNOR2_X1 U475 ( .A(KEYINPUT85), .B(G211GAT), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U477 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n426) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U481 ( .A(n428), .B(n427), .Z(n461) );
  NAND2_X1 U482 ( .A1(n568), .A2(n461), .ZN(n430) );
  XOR2_X1 U483 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n444) );
  XOR2_X1 U485 ( .A(n431), .B(G127GAT), .Z(n433) );
  NAND2_X1 U486 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U488 ( .A(G176GAT), .B(G183GAT), .Z(n435) );
  XNOR2_X1 U489 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U491 ( .A(n437), .B(n436), .Z(n443) );
  XOR2_X1 U492 ( .A(KEYINPUT81), .B(G71GAT), .Z(n439) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(G99GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U496 ( .A(n443), .B(n442), .Z(n524) );
  INV_X1 U497 ( .A(n524), .ZN(n517) );
  NAND2_X1 U498 ( .A1(n444), .A2(n517), .ZN(n448) );
  NOR2_X1 U499 ( .A1(n498), .A2(n448), .ZN(n447) );
  XNOR2_X1 U500 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n445) );
  NOR2_X1 U501 ( .A1(n452), .A2(n448), .ZN(n451) );
  INV_X1 U502 ( .A(KEYINPUT118), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n449), .B(G169GAT), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(G1348GAT) );
  XOR2_X1 U505 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n475) );
  INV_X1 U506 ( .A(n452), .ZN(n528) );
  NAND2_X1 U507 ( .A1(n367), .A2(n528), .ZN(n487) );
  XOR2_X1 U508 ( .A(n461), .B(KEYINPUT28), .Z(n520) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(n514), .ZN(n463) );
  NAND2_X1 U510 ( .A1(n511), .A2(n463), .ZN(n540) );
  NOR2_X1 U511 ( .A1(n520), .A2(n540), .ZN(n526) );
  XOR2_X1 U512 ( .A(n526), .B(KEYINPUT90), .Z(n453) );
  NOR2_X1 U513 ( .A1(n517), .A2(n453), .ZN(n454) );
  XNOR2_X1 U514 ( .A(KEYINPUT91), .B(n454), .ZN(n469) );
  NOR2_X1 U515 ( .A1(n524), .A2(n455), .ZN(n456) );
  XOR2_X1 U516 ( .A(KEYINPUT92), .B(n456), .Z(n457) );
  NAND2_X1 U517 ( .A1(n457), .A2(n461), .ZN(n460) );
  XNOR2_X1 U518 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n458), .B(KEYINPUT25), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n460), .B(n459), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n461), .A2(n517), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT26), .ZN(n567) );
  NAND2_X1 U523 ( .A1(n567), .A2(n463), .ZN(n464) );
  NAND2_X1 U524 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n484) );
  XOR2_X1 U527 ( .A(KEYINPUT16), .B(KEYINPUT80), .Z(n471) );
  NAND2_X1 U528 ( .A1(n552), .A2(n562), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n484), .A2(n472), .ZN(n473) );
  XOR2_X1 U531 ( .A(KEYINPUT95), .B(n473), .Z(n499) );
  NOR2_X1 U532 ( .A1(n487), .A2(n499), .ZN(n482) );
  NAND2_X1 U533 ( .A1(n482), .A2(n511), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U535 ( .A(G1GAT), .B(n476), .Z(G1324GAT) );
  NAND2_X1 U536 ( .A1(n482), .A2(n514), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT35), .B(KEYINPUT98), .Z(n479) );
  NAND2_X1 U539 ( .A1(n482), .A2(n517), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n479), .B(n478), .ZN(n481) );
  XOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT97), .Z(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NAND2_X1 U543 ( .A1(n482), .A2(n520), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT39), .Z(n490) );
  NAND2_X1 U546 ( .A1(n575), .A2(n484), .ZN(n485) );
  NOR2_X1 U547 ( .A1(n485), .A2(n582), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n486), .B(KEYINPUT37), .ZN(n510) );
  NOR2_X1 U549 ( .A1(n510), .A2(n487), .ZN(n488) );
  XNOR2_X1 U550 ( .A(KEYINPUT38), .B(n488), .ZN(n496) );
  NAND2_X1 U551 ( .A1(n511), .A2(n496), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U553 ( .A1(n514), .A2(n496), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G36GAT), .B(n491), .ZN(G1329GAT) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n495) );
  XOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n493) );
  NAND2_X1 U557 ( .A1(n517), .A2(n496), .ZN(n492) );
  XNOR2_X1 U558 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n496), .A2(n520), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n497), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT101), .B(KEYINPUT42), .Z(n501) );
  INV_X1 U563 ( .A(n498), .ZN(n547) );
  NAND2_X1 U564 ( .A1(n569), .A2(n547), .ZN(n509) );
  NOR2_X1 U565 ( .A1(n499), .A2(n509), .ZN(n506) );
  NAND2_X1 U566 ( .A1(n506), .A2(n511), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n506), .A2(n514), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n503), .B(KEYINPUT102), .ZN(n504) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n504), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n506), .A2(n517), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n505), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .Z(n508) );
  NAND2_X1 U575 ( .A1(n506), .A2(n520), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  XOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT103), .Z(n513) );
  NOR2_X1 U578 ( .A1(n510), .A2(n509), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n521), .A2(n511), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n521), .A2(n514), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(KEYINPUT104), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(n516), .ZN(G1337GAT) );
  XOR2_X1 U584 ( .A(G99GAT), .B(KEYINPUT105), .Z(n519) );
  NAND2_X1 U585 ( .A1(n521), .A2(n517), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n541), .ZN(n525) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U592 ( .A(KEYINPUT111), .B(n527), .Z(n533) );
  INV_X1 U593 ( .A(n533), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n528), .A2(n537), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n529), .B(KEYINPUT112), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U598 ( .A1(n537), .A2(n547), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U600 ( .A1(n557), .A2(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(KEYINPUT113), .B(KEYINPUT50), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U605 ( .A1(n537), .A2(n554), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  XOR2_X1 U607 ( .A(G141GAT), .B(KEYINPUT115), .Z(n546) );
  NOR2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U609 ( .A1(n567), .A2(n542), .ZN(n543) );
  XOR2_X1 U610 ( .A(KEYINPUT114), .B(n543), .Z(n555) );
  NAND2_X1 U611 ( .A1(n544), .A2(n555), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1344GAT) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n551) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U615 ( .A1(n555), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n552), .A2(n555), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(n553), .ZN(G1346GAT) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U622 ( .A1(n557), .A2(n448), .ZN(n559) );
  XNOR2_X1 U623 ( .A(G183GAT), .B(KEYINPUT119), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1350GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT120), .B(KEYINPUT58), .Z(n561) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n564) );
  NOR2_X1 U628 ( .A1(n562), .A2(n448), .ZN(n563) );
  XOR2_X1 U629 ( .A(n564), .B(n563), .Z(G1351GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n566) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n581) );
  NOR2_X1 U634 ( .A1(n569), .A2(n581), .ZN(n570) );
  XOR2_X1 U635 ( .A(n571), .B(n570), .Z(G1352GAT) );
  NOR2_X1 U636 ( .A1(n367), .A2(n581), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT123), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G204GAT), .B(n574), .Z(G1353GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n581), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n580) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(n584), .B(n583), .Z(G1355GAT) );
endmodule

