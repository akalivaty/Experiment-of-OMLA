

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593;

  OR2_X1 U323 ( .A1(n485), .A2(n474), .ZN(n475) );
  XNOR2_X1 U324 ( .A(n378), .B(n377), .ZN(n379) );
  NOR2_X1 U325 ( .A1(n455), .A2(n454), .ZN(n456) );
  XNOR2_X1 U326 ( .A(n432), .B(n379), .ZN(n381) );
  XNOR2_X1 U327 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U328 ( .A(n387), .B(n386), .ZN(n391) );
  NOR2_X1 U329 ( .A1(n534), .A2(n447), .ZN(n573) );
  INV_X1 U330 ( .A(G183GAT), .ZN(n449) );
  XNOR2_X1 U331 ( .A(n449), .B(KEYINPUT124), .ZN(n450) );
  XNOR2_X1 U332 ( .A(n478), .B(KEYINPUT44), .ZN(n479) );
  XNOR2_X1 U333 ( .A(n451), .B(n450), .ZN(G1350GAT) );
  XOR2_X1 U334 ( .A(G15GAT), .B(G127GAT), .Z(n312) );
  XOR2_X1 U335 ( .A(G8GAT), .B(G211GAT), .Z(n331) );
  XOR2_X1 U336 ( .A(G22GAT), .B(G155GAT), .Z(n440) );
  XOR2_X1 U337 ( .A(n331), .B(n440), .Z(n292) );
  NAND2_X1 U338 ( .A1(G231GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U339 ( .A(n292), .B(n291), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n312), .B(n293), .ZN(n304) );
  XOR2_X1 U341 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n299) );
  XNOR2_X1 U342 ( .A(G71GAT), .B(G57GAT), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n294), .B(KEYINPUT13), .ZN(n388) );
  XOR2_X1 U344 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n296) );
  XNOR2_X1 U345 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n388), .B(n297), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U349 ( .A(n300), .B(G78GAT), .Z(n302) );
  XOR2_X1 U350 ( .A(KEYINPUT69), .B(G1GAT), .Z(n359) );
  XNOR2_X1 U351 ( .A(n359), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U353 ( .A(n304), .B(n303), .Z(n588) );
  XOR2_X1 U354 ( .A(n588), .B(KEYINPUT112), .Z(n545) );
  XNOR2_X1 U355 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n305), .B(G120GAT), .ZN(n423) );
  XOR2_X1 U357 ( .A(KEYINPUT83), .B(n423), .Z(n307) );
  NAND2_X1 U358 ( .A1(G227GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U360 ( .A(G71GAT), .B(KEYINPUT20), .Z(n309) );
  XNOR2_X1 U361 ( .A(G99GAT), .B(KEYINPUT80), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U363 ( .A(n311), .B(n310), .Z(n314) );
  XOR2_X1 U364 ( .A(G43GAT), .B(G134GAT), .Z(n348) );
  XNOR2_X1 U365 ( .A(n348), .B(n312), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n322) );
  XOR2_X1 U367 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n316) );
  XNOR2_X1 U368 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U370 ( .A(n317), .B(G183GAT), .Z(n319) );
  XNOR2_X1 U371 ( .A(G190GAT), .B(KEYINPUT81), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n321) );
  XOR2_X1 U373 ( .A(G169GAT), .B(G176GAT), .Z(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n338) );
  XNOR2_X1 U375 ( .A(n322), .B(n338), .ZN(n534) );
  INV_X1 U376 ( .A(n331), .ZN(n330) );
  XOR2_X1 U377 ( .A(G64GAT), .B(KEYINPUT73), .Z(n324) );
  XNOR2_X1 U378 ( .A(G204GAT), .B(G92GAT), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n389) );
  XOR2_X1 U380 ( .A(n389), .B(KEYINPUT95), .Z(n329) );
  XOR2_X1 U381 ( .A(KEYINPUT21), .B(G218GAT), .Z(n326) );
  XNOR2_X1 U382 ( .A(KEYINPUT86), .B(KEYINPUT85), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U384 ( .A(n327), .B(G197GAT), .Z(n445) );
  XNOR2_X1 U385 ( .A(G36GAT), .B(n445), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n332) );
  OR2_X1 U387 ( .A1(n330), .A2(n332), .ZN(n334) );
  NAND2_X1 U388 ( .A1(n330), .A2(n332), .ZN(n333) );
  NAND2_X1 U389 ( .A1(n334), .A2(n333), .ZN(n336) );
  NAND2_X1 U390 ( .A1(G226GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X2 U392 ( .A(n338), .B(n337), .ZN(n527) );
  XOR2_X1 U393 ( .A(G99GAT), .B(G85GAT), .Z(n380) );
  XOR2_X1 U394 ( .A(G50GAT), .B(G162GAT), .Z(n441) );
  XOR2_X1 U395 ( .A(n380), .B(n441), .Z(n340) );
  NAND2_X1 U396 ( .A1(G232GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U398 ( .A(KEYINPUT64), .B(KEYINPUT9), .Z(n342) );
  XNOR2_X1 U399 ( .A(G190GAT), .B(KEYINPUT75), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U401 ( .A(n344), .B(n343), .Z(n350) );
  XOR2_X1 U402 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n346) );
  XNOR2_X1 U403 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U407 ( .A(n351), .B(G92GAT), .Z(n355) );
  XOR2_X1 U408 ( .A(G29GAT), .B(G36GAT), .Z(n353) );
  XNOR2_X1 U409 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n362) );
  XNOR2_X1 U411 ( .A(n362), .B(G106GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n572) );
  INV_X1 U413 ( .A(KEYINPUT46), .ZN(n393) );
  XOR2_X1 U414 ( .A(G15GAT), .B(G113GAT), .Z(n357) );
  XNOR2_X1 U415 ( .A(G50GAT), .B(G43GAT), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U417 ( .A(n358), .B(G22GAT), .Z(n361) );
  XNOR2_X1 U418 ( .A(G169GAT), .B(n359), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n366) );
  XOR2_X1 U420 ( .A(n362), .B(KEYINPUT65), .Z(n364) );
  NAND2_X1 U421 ( .A1(G229GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U423 ( .A(n366), .B(n365), .Z(n374) );
  XOR2_X1 U424 ( .A(KEYINPUT68), .B(G8GAT), .Z(n368) );
  XNOR2_X1 U425 ( .A(G141GAT), .B(G197GAT), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U427 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n370) );
  XNOR2_X1 U428 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n578) );
  XOR2_X1 U432 ( .A(G78GAT), .B(G148GAT), .Z(n376) );
  XNOR2_X1 U433 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n432) );
  NAND2_X1 U435 ( .A1(G230GAT), .A2(G233GAT), .ZN(n378) );
  INV_X1 U436 ( .A(KEYINPUT31), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n387) );
  XOR2_X1 U438 ( .A(KEYINPUT70), .B(KEYINPUT32), .Z(n383) );
  XNOR2_X1 U439 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n382) );
  XOR2_X1 U440 ( .A(n383), .B(n382), .Z(n385) );
  XOR2_X1 U441 ( .A(G176GAT), .B(G120GAT), .Z(n384) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n391), .B(n390), .ZN(n583) );
  XOR2_X1 U444 ( .A(n583), .B(KEYINPUT41), .Z(n541) );
  INV_X1 U445 ( .A(n541), .ZN(n567) );
  NAND2_X1 U446 ( .A1(n578), .A2(n567), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n394) );
  NOR2_X1 U448 ( .A1(n572), .A2(n394), .ZN(n395) );
  NAND2_X1 U449 ( .A1(n395), .A2(n545), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n396), .B(KEYINPUT47), .ZN(n402) );
  XNOR2_X1 U451 ( .A(KEYINPUT36), .B(n572), .ZN(n591) );
  NAND2_X1 U452 ( .A1(n588), .A2(n591), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n397), .B(KEYINPUT113), .ZN(n398) );
  XNOR2_X1 U454 ( .A(KEYINPUT45), .B(n398), .ZN(n399) );
  NAND2_X1 U455 ( .A1(n399), .A2(n583), .ZN(n400) );
  NOR2_X1 U456 ( .A1(n400), .A2(n578), .ZN(n401) );
  NOR2_X1 U457 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U458 ( .A(KEYINPUT48), .B(n403), .ZN(n531) );
  NOR2_X1 U459 ( .A1(n527), .A2(n531), .ZN(n404) );
  XNOR2_X1 U460 ( .A(KEYINPUT54), .B(n404), .ZN(n428) );
  XOR2_X1 U461 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n406) );
  XNOR2_X1 U462 ( .A(G1GAT), .B(KEYINPUT92), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U464 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n408) );
  XNOR2_X1 U465 ( .A(KEYINPUT89), .B(KEYINPUT5), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U467 ( .A(n410), .B(n409), .Z(n415) );
  XOR2_X1 U468 ( .A(KEYINPUT1), .B(KEYINPUT94), .Z(n412) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U471 ( .A(KEYINPUT6), .B(n413), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n427) );
  XOR2_X1 U473 ( .A(G85GAT), .B(G162GAT), .Z(n417) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(G134GAT), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U476 ( .A(G57GAT), .B(G155GAT), .Z(n419) );
  XNOR2_X1 U477 ( .A(G127GAT), .B(G148GAT), .ZN(n418) );
  XNOR2_X1 U478 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U479 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U480 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n422), .B(KEYINPUT2), .ZN(n433) );
  XNOR2_X1 U482 ( .A(n423), .B(n433), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U484 ( .A(n427), .B(n426), .Z(n524) );
  NAND2_X1 U485 ( .A1(n428), .A2(n524), .ZN(n576) );
  XOR2_X1 U486 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n430) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U489 ( .A(n431), .B(KEYINPUT87), .Z(n435) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U492 ( .A(G204GAT), .B(G211GAT), .Z(n437) );
  XNOR2_X1 U493 ( .A(KEYINPUT88), .B(KEYINPUT23), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U495 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U498 ( .A(n445), .B(n444), .Z(n464) );
  NOR2_X1 U499 ( .A1(n576), .A2(n464), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n446), .B(KEYINPUT55), .ZN(n447) );
  INV_X1 U501 ( .A(n573), .ZN(n448) );
  NOR2_X1 U502 ( .A1(n545), .A2(n448), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n464), .B(KEYINPUT28), .ZN(n455) );
  INV_X1 U504 ( .A(n455), .ZN(n536) );
  XNOR2_X1 U505 ( .A(n534), .B(KEYINPUT84), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n527), .B(KEYINPUT96), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n452), .B(KEYINPUT27), .ZN(n462) );
  NOR2_X1 U508 ( .A1(n524), .A2(n462), .ZN(n532) );
  NAND2_X1 U509 ( .A1(n453), .A2(n532), .ZN(n454) );
  NAND2_X1 U510 ( .A1(KEYINPUT97), .A2(n456), .ZN(n460) );
  INV_X1 U511 ( .A(KEYINPUT97), .ZN(n458) );
  INV_X1 U512 ( .A(n456), .ZN(n457) );
  NAND2_X1 U513 ( .A1(n458), .A2(n457), .ZN(n459) );
  NAND2_X1 U514 ( .A1(n460), .A2(n459), .ZN(n471) );
  NAND2_X1 U515 ( .A1(n464), .A2(n534), .ZN(n461) );
  XNOR2_X1 U516 ( .A(KEYINPUT26), .B(n461), .ZN(n577) );
  OR2_X1 U517 ( .A1(n462), .A2(n577), .ZN(n468) );
  NOR2_X1 U518 ( .A1(n534), .A2(n527), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n465), .B(KEYINPUT25), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n466), .B(KEYINPUT98), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U523 ( .A1(n469), .A2(n524), .ZN(n470) );
  NAND2_X1 U524 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U525 ( .A(n472), .B(KEYINPUT99), .ZN(n485) );
  INV_X1 U526 ( .A(n588), .ZN(n473) );
  NAND2_X1 U527 ( .A1(n591), .A2(n473), .ZN(n474) );
  XOR2_X1 U528 ( .A(KEYINPUT37), .B(n475), .Z(n498) );
  INV_X1 U529 ( .A(n578), .ZN(n538) );
  NAND2_X1 U530 ( .A1(n567), .A2(n538), .ZN(n476) );
  XOR2_X1 U531 ( .A(KEYINPUT107), .B(n476), .Z(n512) );
  NOR2_X1 U532 ( .A1(n498), .A2(n512), .ZN(n477) );
  XOR2_X1 U533 ( .A(KEYINPUT110), .B(n477), .Z(n529) );
  NOR2_X1 U534 ( .A1(n536), .A2(n529), .ZN(n480) );
  INV_X1 U535 ( .A(G106GAT), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n480), .B(n479), .ZN(G1339GAT) );
  NAND2_X1 U537 ( .A1(n578), .A2(n583), .ZN(n497) );
  INV_X1 U538 ( .A(n497), .ZN(n486) );
  XOR2_X1 U539 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n482) );
  INV_X1 U540 ( .A(n572), .ZN(n548) );
  NAND2_X1 U541 ( .A1(n588), .A2(n548), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n483), .B(KEYINPUT16), .ZN(n484) );
  NOR2_X1 U544 ( .A1(n485), .A2(n484), .ZN(n513) );
  NAND2_X1 U545 ( .A1(n486), .A2(n513), .ZN(n494) );
  NOR2_X1 U546 ( .A1(n524), .A2(n494), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U549 ( .A(G1GAT), .B(n489), .Z(G1324GAT) );
  NOR2_X1 U550 ( .A1(n527), .A2(n494), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(G1325GAT) );
  NOR2_X1 U553 ( .A1(n534), .A2(n494), .ZN(n493) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  NOR2_X1 U556 ( .A1(n536), .A2(n494), .ZN(n495) );
  XOR2_X1 U557 ( .A(KEYINPUT102), .B(n495), .Z(n496) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(n496), .ZN(G1327GAT) );
  INV_X1 U559 ( .A(KEYINPUT38), .ZN(n500) );
  NOR2_X1 U560 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n509) );
  NOR2_X1 U562 ( .A1(n524), .A2(n509), .ZN(n503) );
  XOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT103), .Z(n501) );
  XNOR2_X1 U564 ( .A(KEYINPUT39), .B(n501), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U566 ( .A1(n527), .A2(n509), .ZN(n504) );
  XOR2_X1 U567 ( .A(KEYINPUT104), .B(n504), .Z(n505) );
  XNOR2_X1 U568 ( .A(G36GAT), .B(n505), .ZN(G1329GAT) );
  XNOR2_X1 U569 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n507) );
  NOR2_X1 U570 ( .A1(n534), .A2(n509), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NOR2_X1 U573 ( .A1(n536), .A2(n509), .ZN(n510) );
  XOR2_X1 U574 ( .A(G50GAT), .B(n510), .Z(n511) );
  XNOR2_X1 U575 ( .A(KEYINPUT106), .B(n511), .ZN(G1331GAT) );
  INV_X1 U576 ( .A(n512), .ZN(n514) );
  NAND2_X1 U577 ( .A1(n514), .A2(n513), .ZN(n520) );
  NOR2_X1 U578 ( .A1(n524), .A2(n520), .ZN(n515) );
  XOR2_X1 U579 ( .A(n515), .B(KEYINPUT42), .Z(n516) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(n516), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n527), .A2(n520), .ZN(n517) );
  XOR2_X1 U582 ( .A(G64GAT), .B(n517), .Z(G1333GAT) );
  NOR2_X1 U583 ( .A1(n534), .A2(n520), .ZN(n518) );
  XOR2_X1 U584 ( .A(KEYINPUT108), .B(n518), .Z(n519) );
  XNOR2_X1 U585 ( .A(G71GAT), .B(n519), .ZN(G1334GAT) );
  NOR2_X1 U586 ( .A1(n536), .A2(n520), .ZN(n522) );
  XNOR2_X1 U587 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U589 ( .A(G78GAT), .B(n523), .Z(G1335GAT) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n526) );
  NOR2_X1 U591 ( .A1(n524), .A2(n529), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1336GAT) );
  NOR2_X1 U593 ( .A1(n527), .A2(n529), .ZN(n528) );
  XOR2_X1 U594 ( .A(G92GAT), .B(n528), .Z(G1337GAT) );
  NOR2_X1 U595 ( .A1(n534), .A2(n529), .ZN(n530) );
  XOR2_X1 U596 ( .A(G99GAT), .B(n530), .Z(G1338GAT) );
  INV_X1 U597 ( .A(n531), .ZN(n533) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n553) );
  NOR2_X1 U599 ( .A1(n534), .A2(n553), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U601 ( .A(KEYINPUT114), .B(n537), .ZN(n549) );
  NOR2_X1 U602 ( .A1(n549), .A2(n538), .ZN(n540) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(G1340GAT) );
  XNOR2_X1 U605 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n543) );
  NOR2_X1 U606 ( .A1(n541), .A2(n549), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U609 ( .A1(n549), .A2(n545), .ZN(n546) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(n546), .Z(n547) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  NOR2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U613 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U615 ( .A(G134GAT), .B(n552), .Z(G1343GAT) );
  NOR2_X1 U616 ( .A1(n553), .A2(n577), .ZN(n554) );
  XNOR2_X1 U617 ( .A(n554), .B(KEYINPUT118), .ZN(n562) );
  NAND2_X1 U618 ( .A1(n578), .A2(n562), .ZN(n555) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U621 ( .A1(n562), .A2(n567), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n560) );
  NAND2_X1 U625 ( .A1(n562), .A2(n588), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n561), .ZN(G1346GAT) );
  XOR2_X1 U628 ( .A(G162GAT), .B(KEYINPUT121), .Z(n564) );
  NAND2_X1 U629 ( .A1(n572), .A2(n562), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n573), .A2(n578), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(n566), .ZN(G1348GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n569) );
  NAND2_X1 U635 ( .A1(n573), .A2(n567), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT56), .Z(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT58), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G190GAT), .B(n575), .ZN(G1351GAT) );
  XOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT60), .Z(n580) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n590) );
  NAND2_X1 U644 ( .A1(n590), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n586) );
  INV_X1 U649 ( .A(n583), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n590), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(n587), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n590), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n592), .B(KEYINPUT62), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

