

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742;

  XNOR2_X1 U368 ( .A(n437), .B(n436), .ZN(n671) );
  INV_X1 U369 ( .A(G953), .ZN(n735) );
  AND2_X1 U370 ( .A1(n367), .A2(n368), .ZN(n354) );
  AND2_X1 U371 ( .A1(n516), .A2(n382), .ZN(n381) );
  XNOR2_X2 U372 ( .A(G128), .B(G143), .ZN(n430) );
  XNOR2_X1 U373 ( .A(n553), .B(KEYINPUT45), .ZN(n708) );
  NAND2_X1 U374 ( .A1(n354), .A2(n365), .ZN(n364) );
  NAND2_X1 U375 ( .A1(n399), .A2(n398), .ZN(n390) );
  AND2_X1 U376 ( .A1(n399), .A2(n395), .ZN(n375) );
  XNOR2_X1 U377 ( .A(n621), .B(n620), .ZN(n622) );
  OR2_X1 U378 ( .A1(n610), .A2(n350), .ZN(n396) );
  XNOR2_X1 U379 ( .A(n411), .B(n410), .ZN(n531) );
  XNOR2_X1 U380 ( .A(n378), .B(n442), .ZN(n610) );
  AND2_X1 U381 ( .A1(n398), .A2(n503), .ZN(n395) );
  XNOR2_X1 U382 ( .A(n393), .B(n716), .ZN(n442) );
  XNOR2_X1 U383 ( .A(n425), .B(n414), .ZN(n717) );
  XNOR2_X1 U384 ( .A(n348), .B(n413), .ZN(n425) );
  XNOR2_X1 U385 ( .A(KEYINPUT16), .B(G122), .ZN(n414) );
  XNOR2_X1 U386 ( .A(KEYINPUT93), .B(KEYINPUT18), .ZN(n417) );
  BUF_X1 U387 ( .A(n619), .Z(n345) );
  XNOR2_X1 U388 ( .A(n608), .B(KEYINPUT2), .ZN(n346) );
  XNOR2_X1 U389 ( .A(n364), .B(n389), .ZN(n619) );
  XNOR2_X1 U390 ( .A(n608), .B(KEYINPUT2), .ZN(n650) );
  NAND2_X1 U391 ( .A1(n708), .A2(n733), .ZN(n608) );
  XNOR2_X1 U392 ( .A(KEYINPUT13), .B(G475), .ZN(n410) );
  OR2_X1 U393 ( .A1(n699), .A2(G902), .ZN(n411) );
  XNOR2_X1 U394 ( .A(G119), .B(KEYINPUT3), .ZN(n413) );
  XNOR2_X1 U395 ( .A(n427), .B(n422), .ZN(n393) );
  XNOR2_X1 U396 ( .A(n575), .B(n387), .ZN(n407) );
  INV_X1 U397 ( .A(KEYINPUT83), .ZN(n387) );
  XNOR2_X1 U398 ( .A(n363), .B(KEYINPUT73), .ZN(n362) );
  AND2_X1 U399 ( .A1(n643), .A2(n645), .ZN(n657) );
  XNOR2_X1 U400 ( .A(KEYINPUT4), .B(KEYINPUT65), .ZN(n724) );
  XNOR2_X1 U401 ( .A(n360), .B(n358), .ZN(n489) );
  XNOR2_X1 U402 ( .A(KEYINPUT8), .B(KEYINPUT66), .ZN(n360) );
  NOR2_X1 U403 ( .A1(n359), .A2(G953), .ZN(n358) );
  NOR2_X1 U404 ( .A1(G953), .A2(G237), .ZN(n479) );
  XNOR2_X1 U405 ( .A(n426), .B(G131), .ZN(n388) );
  XNOR2_X1 U406 ( .A(G101), .B(n724), .ZN(n427) );
  XNOR2_X1 U407 ( .A(G116), .B(G107), .ZN(n493) );
  INV_X1 U408 ( .A(KEYINPUT9), .ZN(n357) );
  XOR2_X1 U409 ( .A(G122), .B(KEYINPUT7), .Z(n491) );
  INV_X1 U410 ( .A(KEYINPUT80), .ZN(n402) );
  XNOR2_X1 U411 ( .A(n483), .B(n403), .ZN(n723) );
  INV_X1 U412 ( .A(KEYINPUT96), .ZN(n403) );
  AND2_X1 U413 ( .A1(n374), .A2(n372), .ZN(n371) );
  NOR2_X1 U414 ( .A1(n535), .A2(n529), .ZN(n386) );
  XNOR2_X1 U415 ( .A(n580), .B(KEYINPUT19), .ZN(n565) );
  NOR2_X1 U416 ( .A1(n704), .A2(G902), .ZN(n495) );
  XNOR2_X1 U417 ( .A(n488), .B(n487), .ZN(n699) );
  XNOR2_X1 U418 ( .A(n486), .B(n347), .ZN(n487) );
  AND2_X1 U419 ( .A1(n614), .A2(G953), .ZN(n707) );
  NAND2_X1 U420 ( .A1(n406), .A2(n361), .ZN(n405) );
  XNOR2_X1 U421 ( .A(n657), .B(n408), .ZN(n555) );
  INV_X1 U422 ( .A(KEYINPUT84), .ZN(n408) );
  NAND2_X1 U423 ( .A1(G234), .A2(G237), .ZN(n466) );
  INV_X1 U424 ( .A(KEYINPUT107), .ZN(n525) );
  NAND2_X1 U425 ( .A1(n349), .A2(n609), .ZN(n398) );
  NAND2_X1 U426 ( .A1(n373), .A2(n351), .ZN(n372) );
  INV_X1 U427 ( .A(n396), .ZN(n373) );
  AND2_X1 U428 ( .A1(n390), .A2(n351), .ZN(n370) );
  BUF_X1 U429 ( .A(n513), .Z(n562) );
  XNOR2_X1 U430 ( .A(G119), .B(G140), .ZN(n453) );
  XNOR2_X1 U431 ( .A(G137), .B(G128), .ZN(n446) );
  XOR2_X1 U432 ( .A(G122), .B(G104), .Z(n485) );
  XNOR2_X1 U433 ( .A(G143), .B(G113), .ZN(n484) );
  XNOR2_X1 U434 ( .A(n457), .B(KEYINPUT15), .ZN(n609) );
  INV_X1 U435 ( .A(KEYINPUT0), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n391), .B(n462), .ZN(n559) );
  XNOR2_X1 U437 ( .A(n392), .B(n461), .ZN(n391) );
  XNOR2_X1 U438 ( .A(n671), .B(n512), .ZN(n578) );
  XNOR2_X1 U439 ( .A(n425), .B(n388), .ZN(n429) );
  XNOR2_X1 U440 ( .A(n492), .B(n355), .ZN(n704) );
  XNOR2_X1 U441 ( .A(n494), .B(n356), .ZN(n355) );
  XNOR2_X1 U442 ( .A(n493), .B(n357), .ZN(n356) );
  XNOR2_X1 U443 ( .A(n441), .B(n400), .ZN(n394) );
  XNOR2_X1 U444 ( .A(n723), .B(n401), .ZN(n400) );
  XNOR2_X1 U445 ( .A(n443), .B(n402), .ZN(n401) );
  XNOR2_X1 U446 ( .A(n610), .B(n611), .ZN(n612) );
  INV_X1 U447 ( .A(KEYINPUT35), .ZN(n389) );
  AND2_X1 U448 ( .A1(n572), .A2(n571), .ZN(n639) );
  AND2_X1 U449 ( .A1(n498), .A2(n530), .ZN(n499) );
  NOR2_X1 U450 ( .A1(n701), .A2(n707), .ZN(n702) );
  XNOR2_X1 U451 ( .A(n409), .B(n700), .ZN(n701) );
  XOR2_X1 U452 ( .A(n485), .B(n484), .Z(n347) );
  XOR2_X1 U453 ( .A(G113), .B(G116), .Z(n348) );
  XOR2_X1 U454 ( .A(n423), .B(KEYINPUT82), .Z(n349) );
  OR2_X1 U455 ( .A1(n349), .A2(n609), .ZN(n350) );
  NAND2_X1 U456 ( .A1(n371), .A2(n369), .ZN(n580) );
  XNOR2_X1 U457 ( .A(n384), .B(KEYINPUT22), .ZN(n520) );
  AND2_X1 U458 ( .A1(n653), .A2(KEYINPUT91), .ZN(n351) );
  INV_X1 U459 ( .A(G234), .ZN(n359) );
  NOR2_X1 U460 ( .A1(n653), .A2(KEYINPUT91), .ZN(n352) );
  XOR2_X1 U461 ( .A(KEYINPUT81), .B(KEYINPUT34), .Z(n529) );
  XNOR2_X1 U462 ( .A(n394), .B(n442), .ZN(n694) );
  AND2_X1 U463 ( .A1(n609), .A2(G475), .ZN(n353) );
  NAND2_X1 U464 ( .A1(n366), .A2(n386), .ZN(n365) );
  NAND2_X1 U465 ( .A1(n362), .A2(n566), .ZN(n361) );
  NAND2_X1 U466 ( .A1(n555), .A2(n554), .ZN(n363) );
  INV_X1 U467 ( .A(n651), .ZN(n366) );
  NAND2_X1 U468 ( .A1(n651), .A2(n529), .ZN(n367) );
  AND2_X1 U469 ( .A1(n385), .A2(n570), .ZN(n368) );
  NOR2_X1 U470 ( .A1(n370), .A2(n352), .ZN(n369) );
  NAND2_X1 U471 ( .A1(n375), .A2(n396), .ZN(n374) );
  INV_X1 U472 ( .A(n377), .ZN(n535) );
  NAND2_X1 U473 ( .A1(n377), .A2(n510), .ZN(n384) );
  XNOR2_X2 U474 ( .A(n508), .B(n376), .ZN(n377) );
  NAND2_X1 U475 ( .A1(n377), .A2(n539), .ZN(n631) );
  XNOR2_X1 U476 ( .A(n379), .B(n717), .ZN(n378) );
  XNOR2_X1 U477 ( .A(n380), .B(n419), .ZN(n379) );
  XNOR2_X1 U478 ( .A(n418), .B(n431), .ZN(n380) );
  NOR2_X1 U479 ( .A1(n520), .A2(n578), .ZN(n517) );
  NAND2_X1 U480 ( .A1(n383), .A2(n381), .ZN(n519) );
  INV_X1 U481 ( .A(n578), .ZN(n382) );
  INV_X1 U482 ( .A(n520), .ZN(n383) );
  NAND2_X1 U483 ( .A1(n535), .A2(n529), .ZN(n385) );
  XNOR2_X2 U484 ( .A(n528), .B(n527), .ZN(n651) );
  INV_X1 U485 ( .A(n390), .ZN(n397) );
  INV_X1 U486 ( .A(n559), .ZN(n666) );
  NAND2_X1 U487 ( .A1(n463), .A2(G217), .ZN(n392) );
  INV_X1 U488 ( .A(n430), .ZN(n431) );
  NAND2_X1 U489 ( .A1(n431), .A2(n432), .ZN(n433) );
  XNOR2_X2 U490 ( .A(n729), .B(G146), .ZN(n441) );
  XNOR2_X2 U491 ( .A(n494), .B(G137), .ZN(n729) );
  NAND2_X2 U492 ( .A1(n433), .A2(n434), .ZN(n494) );
  XNOR2_X2 U493 ( .A(G146), .B(G125), .ZN(n451) );
  NAND2_X1 U494 ( .A1(n397), .A2(n396), .ZN(n602) );
  NAND2_X1 U495 ( .A1(n610), .A2(n349), .ZN(n399) );
  NAND2_X1 U496 ( .A1(n404), .A2(n594), .ZN(n596) );
  XNOR2_X1 U497 ( .A(n405), .B(KEYINPUT67), .ZN(n404) );
  NOR2_X1 U498 ( .A1(n585), .A2(n407), .ZN(n406) );
  XNOR2_X2 U499 ( .A(n499), .B(KEYINPUT105), .ZN(n643) );
  AND2_X2 U500 ( .A1(n650), .A2(n609), .ZN(n703) );
  NAND2_X1 U501 ( .A1(n346), .A2(n353), .ZN(n409) );
  XNOR2_X1 U502 ( .A(n513), .B(KEYINPUT1), .ZN(n523) );
  NOR2_X2 U503 ( .A1(n694), .A2(G902), .ZN(n445) );
  AND2_X1 U504 ( .A1(n479), .A2(G210), .ZN(n412) );
  BUF_X1 U505 ( .A(n651), .Z(n683) );
  XNOR2_X1 U506 ( .A(n427), .B(n412), .ZN(n428) );
  XNOR2_X1 U507 ( .A(n429), .B(n428), .ZN(n435) );
  INV_X1 U508 ( .A(n643), .ZN(n500) );
  XNOR2_X1 U509 ( .A(n694), .B(n695), .ZN(n696) );
  BUF_X1 U510 ( .A(n523), .Z(n663) );
  XOR2_X1 U511 ( .A(KEYINPUT94), .B(KEYINPUT17), .Z(n416) );
  NAND2_X1 U512 ( .A1(G224), .A2(n735), .ZN(n415) );
  XNOR2_X1 U513 ( .A(n416), .B(n415), .ZN(n419) );
  XNOR2_X1 U514 ( .A(n451), .B(n417), .ZN(n418) );
  XOR2_X1 U515 ( .A(G104), .B(G107), .Z(n421) );
  XNOR2_X1 U516 ( .A(KEYINPUT92), .B(G110), .ZN(n420) );
  XNOR2_X1 U517 ( .A(n421), .B(n420), .ZN(n716) );
  XOR2_X1 U518 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n422) );
  OR2_X1 U519 ( .A1(G237), .A2(G902), .ZN(n424) );
  NAND2_X1 U520 ( .A1(G210), .A2(n424), .ZN(n423) );
  XOR2_X1 U521 ( .A(KEYINPUT38), .B(n602), .Z(n652) );
  INV_X1 U522 ( .A(n652), .ZN(n440) );
  NAND2_X1 U523 ( .A1(G214), .A2(n424), .ZN(n653) );
  XOR2_X1 U524 ( .A(KEYINPUT5), .B(KEYINPUT76), .Z(n426) );
  NAND2_X1 U525 ( .A1(G134), .A2(n430), .ZN(n434) );
  INV_X1 U526 ( .A(G134), .ZN(n432) );
  XNOR2_X1 U527 ( .A(n441), .B(n435), .ZN(n621) );
  NOR2_X1 U528 ( .A1(G902), .A2(n621), .ZN(n437) );
  XNOR2_X1 U529 ( .A(G472), .B(KEYINPUT99), .ZN(n436) );
  NAND2_X1 U530 ( .A1(n653), .A2(n671), .ZN(n439) );
  XNOR2_X1 U531 ( .A(KEYINPUT112), .B(KEYINPUT30), .ZN(n438) );
  XNOR2_X1 U532 ( .A(n439), .B(n438), .ZN(n568) );
  NOR2_X1 U533 ( .A1(n440), .A2(n568), .ZN(n475) );
  XOR2_X1 U534 ( .A(G131), .B(G140), .Z(n483) );
  NAND2_X1 U535 ( .A1(G227), .A2(n735), .ZN(n443) );
  INV_X1 U536 ( .A(G469), .ZN(n444) );
  XNOR2_X2 U537 ( .A(n445), .B(n444), .ZN(n513) );
  NAND2_X1 U538 ( .A1(n489), .A2(G221), .ZN(n450) );
  XNOR2_X1 U539 ( .A(n446), .B(KEYINPUT23), .ZN(n448) );
  XNOR2_X1 U540 ( .A(KEYINPUT68), .B(KEYINPUT79), .ZN(n447) );
  XNOR2_X1 U541 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U542 ( .A(n450), .B(n449), .ZN(n456) );
  XNOR2_X1 U543 ( .A(n451), .B(KEYINPUT10), .ZN(n725) );
  XNOR2_X1 U544 ( .A(G110), .B(KEYINPUT24), .ZN(n452) );
  XNOR2_X1 U545 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U546 ( .A(n725), .B(n454), .ZN(n455) );
  XNOR2_X1 U547 ( .A(n456), .B(n455), .ZN(n628) );
  INV_X1 U548 ( .A(G902), .ZN(n457) );
  NAND2_X1 U549 ( .A1(n628), .A2(n457), .ZN(n462) );
  OR2_X1 U550 ( .A1(n609), .A2(n359), .ZN(n459) );
  XOR2_X1 U551 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n458) );
  XNOR2_X1 U552 ( .A(n459), .B(n458), .ZN(n463) );
  XNOR2_X1 U553 ( .A(KEYINPUT78), .B(KEYINPUT98), .ZN(n460) );
  XNOR2_X1 U554 ( .A(n460), .B(KEYINPUT25), .ZN(n461) );
  NAND2_X1 U555 ( .A1(n463), .A2(G221), .ZN(n465) );
  INV_X1 U556 ( .A(KEYINPUT21), .ZN(n464) );
  XNOR2_X1 U557 ( .A(n465), .B(n464), .ZN(n665) );
  AND2_X1 U558 ( .A1(n666), .A2(n665), .ZN(n662) );
  NAND2_X1 U559 ( .A1(n562), .A2(n662), .ZN(n538) );
  XNOR2_X1 U560 ( .A(n466), .B(KEYINPUT14), .ZN(n467) );
  XNOR2_X1 U561 ( .A(KEYINPUT74), .B(n467), .ZN(n471) );
  NAND2_X1 U562 ( .A1(G952), .A2(n471), .ZN(n681) );
  NOR2_X1 U563 ( .A1(G953), .A2(n681), .ZN(n469) );
  INV_X1 U564 ( .A(KEYINPUT95), .ZN(n468) );
  XNOR2_X1 U565 ( .A(n469), .B(n468), .ZN(n506) );
  AND2_X1 U566 ( .A1(G953), .A2(G902), .ZN(n470) );
  NAND2_X1 U567 ( .A1(n471), .A2(n470), .ZN(n504) );
  XOR2_X1 U568 ( .A(n504), .B(KEYINPUT109), .Z(n472) );
  NOR2_X1 U569 ( .A1(n472), .A2(G900), .ZN(n473) );
  NOR2_X1 U570 ( .A1(n506), .A2(n473), .ZN(n557) );
  OR2_X1 U571 ( .A1(n538), .A2(n557), .ZN(n474) );
  XNOR2_X1 U572 ( .A(n474), .B(KEYINPUT77), .ZN(n571) );
  NAND2_X1 U573 ( .A1(n475), .A2(n571), .ZN(n476) );
  XNOR2_X1 U574 ( .A(n476), .B(KEYINPUT39), .ZN(n501) );
  XOR2_X1 U575 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n478) );
  XNOR2_X1 U576 ( .A(KEYINPUT12), .B(KEYINPUT101), .ZN(n477) );
  XNOR2_X1 U577 ( .A(n478), .B(n477), .ZN(n481) );
  NAND2_X1 U578 ( .A1(G214), .A2(n479), .ZN(n480) );
  XNOR2_X1 U579 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U580 ( .A(n482), .B(n725), .Z(n488) );
  XNOR2_X1 U581 ( .A(n483), .B(KEYINPUT11), .ZN(n486) );
  XOR2_X1 U582 ( .A(KEYINPUT104), .B(n531), .Z(n498) );
  INV_X1 U583 ( .A(n498), .ZN(n497) );
  NAND2_X1 U584 ( .A1(G217), .A2(n489), .ZN(n490) );
  XNOR2_X1 U585 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U586 ( .A(G478), .B(n495), .ZN(n530) );
  INV_X1 U587 ( .A(n530), .ZN(n496) );
  NAND2_X1 U588 ( .A1(n497), .A2(n496), .ZN(n645) );
  INV_X1 U589 ( .A(n645), .ZN(n540) );
  NAND2_X1 U590 ( .A1(n501), .A2(n540), .ZN(n605) );
  XNOR2_X1 U591 ( .A(n605), .B(G134), .ZN(G36) );
  NAND2_X1 U592 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U593 ( .A(n502), .B(KEYINPUT40), .ZN(n591) );
  XNOR2_X1 U594 ( .A(n591), .B(G131), .ZN(G33) );
  INV_X1 U595 ( .A(KEYINPUT91), .ZN(n503) );
  NOR2_X1 U596 ( .A1(G898), .A2(n504), .ZN(n505) );
  OR2_X1 U597 ( .A1(n506), .A2(n505), .ZN(n507) );
  NAND2_X1 U598 ( .A1(n565), .A2(n507), .ZN(n508) );
  NAND2_X1 U599 ( .A1(n531), .A2(n530), .ZN(n655) );
  INV_X1 U600 ( .A(n655), .ZN(n509) );
  AND2_X1 U601 ( .A1(n665), .A2(n509), .ZN(n510) );
  INV_X1 U602 ( .A(KEYINPUT106), .ZN(n511) );
  XNOR2_X1 U603 ( .A(n511), .B(KEYINPUT6), .ZN(n512) );
  XNOR2_X1 U604 ( .A(n517), .B(KEYINPUT88), .ZN(n515) );
  NOR2_X1 U605 ( .A1(n663), .A2(n559), .ZN(n514) );
  NAND2_X1 U606 ( .A1(n515), .A2(n514), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(G101), .ZN(G3) );
  AND2_X1 U608 ( .A1(n663), .A2(n559), .ZN(n516) );
  XOR2_X1 U609 ( .A(KEYINPUT64), .B(KEYINPUT32), .Z(n518) );
  XNOR2_X1 U610 ( .A(n519), .B(n518), .ZN(n740) );
  NOR2_X1 U611 ( .A1(n671), .A2(n666), .ZN(n521) );
  NAND2_X1 U612 ( .A1(n383), .A2(n521), .ZN(n522) );
  NOR2_X1 U613 ( .A1(n522), .A2(n663), .ZN(n635) );
  NOR2_X1 U614 ( .A1(n740), .A2(n635), .ZN(n533) );
  NAND2_X1 U615 ( .A1(n523), .A2(n662), .ZN(n524) );
  XNOR2_X2 U616 ( .A(n524), .B(KEYINPUT75), .ZN(n534) );
  XNOR2_X1 U617 ( .A(n534), .B(n525), .ZN(n526) );
  NAND2_X1 U618 ( .A1(n526), .A2(n578), .ZN(n528) );
  XNOR2_X1 U619 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n527) );
  NOR2_X1 U620 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U621 ( .A(n532), .B(KEYINPUT108), .ZN(n570) );
  NAND2_X1 U622 ( .A1(n533), .A2(n619), .ZN(n547) );
  NAND2_X1 U623 ( .A1(n547), .A2(KEYINPUT44), .ZN(n545) );
  NAND2_X1 U624 ( .A1(n534), .A2(n671), .ZN(n674) );
  NOR2_X1 U625 ( .A1(n535), .A2(n674), .ZN(n537) );
  XNOR2_X1 U626 ( .A(KEYINPUT100), .B(KEYINPUT31), .ZN(n536) );
  XNOR2_X1 U627 ( .A(n537), .B(n536), .ZN(n646) );
  NOR2_X1 U628 ( .A1(n538), .A2(n671), .ZN(n539) );
  NAND2_X1 U629 ( .A1(n646), .A2(n631), .ZN(n541) );
  NAND2_X1 U630 ( .A1(n541), .A2(n555), .ZN(n543) );
  AND2_X1 U631 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U632 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U633 ( .A(n546), .B(KEYINPUT89), .ZN(n552) );
  INV_X1 U634 ( .A(n547), .ZN(n549) );
  INV_X1 U635 ( .A(KEYINPUT44), .ZN(n548) );
  NAND2_X1 U636 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U637 ( .A(n550), .B(KEYINPUT72), .ZN(n551) );
  NAND2_X1 U638 ( .A1(n552), .A2(n551), .ZN(n553) );
  INV_X1 U639 ( .A(KEYINPUT47), .ZN(n554) );
  XNOR2_X1 U640 ( .A(KEYINPUT28), .B(KEYINPUT113), .ZN(n561) );
  INV_X1 U641 ( .A(n665), .ZN(n556) );
  NOR2_X1 U642 ( .A1(n557), .A2(n556), .ZN(n558) );
  AND2_X1 U643 ( .A1(n559), .A2(n558), .ZN(n576) );
  NAND2_X1 U644 ( .A1(n671), .A2(n576), .ZN(n560) );
  XOR2_X1 U645 ( .A(n561), .B(n560), .Z(n564) );
  INV_X1 U646 ( .A(n562), .ZN(n563) );
  NOR2_X1 U647 ( .A1(n564), .A2(n563), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n587), .A2(n565), .ZN(n641) );
  INV_X1 U649 ( .A(n641), .ZN(n566) );
  INV_X1 U650 ( .A(n602), .ZN(n567) );
  NOR2_X1 U651 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U652 ( .A1(n570), .A2(n569), .ZN(n572) );
  XNOR2_X1 U653 ( .A(n639), .B(KEYINPUT85), .ZN(n574) );
  NAND2_X1 U654 ( .A1(n657), .A2(KEYINPUT47), .ZN(n573) );
  NAND2_X1 U655 ( .A1(n574), .A2(n573), .ZN(n575) );
  INV_X1 U656 ( .A(n576), .ZN(n577) );
  NOR2_X1 U657 ( .A1(n643), .A2(n577), .ZN(n579) );
  NAND2_X1 U658 ( .A1(n579), .A2(n578), .ZN(n597) );
  NOR2_X1 U659 ( .A1(n597), .A2(n580), .ZN(n582) );
  XNOR2_X1 U660 ( .A(KEYINPUT36), .B(KEYINPUT90), .ZN(n581) );
  XNOR2_X1 U661 ( .A(n582), .B(n581), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n583), .A2(n663), .ZN(n649) );
  NAND2_X1 U663 ( .A1(KEYINPUT47), .A2(n641), .ZN(n584) );
  NAND2_X1 U664 ( .A1(n649), .A2(n584), .ZN(n585) );
  NAND2_X1 U665 ( .A1(n653), .A2(n652), .ZN(n658) );
  NOR2_X1 U666 ( .A1(n655), .A2(n658), .ZN(n586) );
  XNOR2_X1 U667 ( .A(KEYINPUT41), .B(n586), .ZN(n682) );
  INV_X1 U668 ( .A(n682), .ZN(n588) );
  NAND2_X1 U669 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U670 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n589) );
  XNOR2_X1 U671 ( .A(n590), .B(n589), .ZN(n739) );
  NAND2_X1 U672 ( .A1(n739), .A2(n591), .ZN(n593) );
  XNOR2_X1 U673 ( .A(KEYINPUT87), .B(KEYINPUT46), .ZN(n592) );
  XNOR2_X1 U674 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U675 ( .A(KEYINPUT86), .B(KEYINPUT48), .ZN(n595) );
  XNOR2_X1 U676 ( .A(n596), .B(n595), .ZN(n607) );
  INV_X1 U677 ( .A(n597), .ZN(n598) );
  NAND2_X1 U678 ( .A1(n598), .A2(n653), .ZN(n599) );
  XNOR2_X1 U679 ( .A(KEYINPUT110), .B(n599), .ZN(n600) );
  NOR2_X1 U680 ( .A1(n663), .A2(n600), .ZN(n601) );
  XNOR2_X1 U681 ( .A(n601), .B(KEYINPUT43), .ZN(n603) );
  NOR2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U683 ( .A(n604), .B(KEYINPUT111), .ZN(n741) );
  NAND2_X1 U684 ( .A1(n741), .A2(n605), .ZN(n606) );
  NOR2_X2 U685 ( .A1(n607), .A2(n606), .ZN(n733) );
  NAND2_X1 U686 ( .A1(n703), .A2(G210), .ZN(n613) );
  XNOR2_X1 U687 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n613), .B(n612), .ZN(n615) );
  INV_X1 U689 ( .A(G952), .ZN(n614) );
  INV_X1 U690 ( .A(n707), .ZN(n624) );
  NAND2_X1 U691 ( .A1(n615), .A2(n624), .ZN(n617) );
  INV_X1 U692 ( .A(KEYINPUT56), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n617), .B(n616), .ZN(G51) );
  XOR2_X1 U694 ( .A(G122), .B(KEYINPUT127), .Z(n618) );
  XNOR2_X1 U695 ( .A(n345), .B(n618), .ZN(G24) );
  NAND2_X1 U696 ( .A1(n703), .A2(G472), .ZN(n623) );
  XNOR2_X1 U697 ( .A(KEYINPUT115), .B(KEYINPUT62), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n623), .B(n622), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n626), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U701 ( .A1(n703), .A2(G217), .ZN(n627) );
  XOR2_X1 U702 ( .A(n628), .B(n627), .Z(n629) );
  NOR2_X1 U703 ( .A1(n629), .A2(n707), .ZN(G66) );
  NOR2_X1 U704 ( .A1(n643), .A2(n631), .ZN(n630) );
  XOR2_X1 U705 ( .A(G104), .B(n630), .Z(G6) );
  NOR2_X1 U706 ( .A1(n645), .A2(n631), .ZN(n633) );
  XNOR2_X1 U707 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U709 ( .A(G107), .B(n634), .ZN(G9) );
  XOR2_X1 U710 ( .A(G110), .B(n635), .Z(G12) );
  NOR2_X1 U711 ( .A1(n645), .A2(n641), .ZN(n637) );
  XNOR2_X1 U712 ( .A(KEYINPUT29), .B(KEYINPUT116), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U714 ( .A(G128), .B(n638), .ZN(G30) );
  XNOR2_X1 U715 ( .A(n639), .B(G143), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n640), .B(KEYINPUT117), .ZN(G45) );
  NOR2_X1 U717 ( .A1(n643), .A2(n641), .ZN(n642) );
  XOR2_X1 U718 ( .A(G146), .B(n642), .Z(G48) );
  NOR2_X1 U719 ( .A1(n646), .A2(n643), .ZN(n644) );
  XOR2_X1 U720 ( .A(G113), .B(n644), .Z(G15) );
  NOR2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U722 ( .A(G116), .B(n647), .Z(G18) );
  XOR2_X1 U723 ( .A(G125), .B(KEYINPUT37), .Z(n648) );
  XNOR2_X1 U724 ( .A(n649), .B(n648), .ZN(G27) );
  INV_X1 U725 ( .A(n346), .ZN(n689) );
  NOR2_X1 U726 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U727 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n656), .B(KEYINPUT120), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U731 ( .A1(n683), .A2(n661), .ZN(n678) );
  NOR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U733 ( .A(KEYINPUT50), .B(n664), .Z(n669) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n667), .B(KEYINPUT49), .ZN(n668) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(KEYINPUT119), .ZN(n673) );
  NAND2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U740 ( .A(KEYINPUT51), .B(n675), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n682), .A2(n676), .ZN(n677) );
  NOR2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U743 ( .A(n679), .B(KEYINPUT52), .ZN(n680) );
  NOR2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n686) );
  NOR2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U746 ( .A(KEYINPUT121), .B(n684), .Z(n685) );
  NOR2_X1 U747 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U748 ( .A(n687), .B(KEYINPUT122), .ZN(n688) );
  NAND2_X1 U749 ( .A1(n689), .A2(n688), .ZN(n691) );
  INV_X1 U750 ( .A(KEYINPUT123), .ZN(n690) );
  XNOR2_X1 U751 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U752 ( .A1(G953), .A2(n692), .ZN(n693) );
  XNOR2_X1 U753 ( .A(KEYINPUT53), .B(n693), .ZN(G75) );
  NAND2_X1 U754 ( .A1(n703), .A2(G469), .ZN(n697) );
  XOR2_X1 U755 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n695) );
  XNOR2_X1 U756 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U757 ( .A1(n707), .A2(n698), .ZN(G54) );
  XOR2_X1 U758 ( .A(n699), .B(KEYINPUT59), .Z(n700) );
  XNOR2_X1 U759 ( .A(n702), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U760 ( .A1(n703), .A2(G478), .ZN(n705) );
  XNOR2_X1 U761 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U762 ( .A1(n707), .A2(n706), .ZN(G63) );
  INV_X1 U763 ( .A(n708), .ZN(n709) );
  NOR2_X1 U764 ( .A1(n709), .A2(G953), .ZN(n715) );
  XOR2_X1 U765 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n711) );
  NAND2_X1 U766 ( .A1(G224), .A2(G953), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n711), .B(n710), .ZN(n713) );
  INV_X1 U768 ( .A(G898), .ZN(n712) );
  NOR2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U770 ( .A1(n715), .A2(n714), .ZN(n722) );
  XNOR2_X1 U771 ( .A(G101), .B(n716), .ZN(n718) );
  XNOR2_X1 U772 ( .A(n718), .B(n717), .ZN(n720) );
  NOR2_X1 U773 ( .A1(G898), .A2(n735), .ZN(n719) );
  NOR2_X1 U774 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U775 ( .A(n722), .B(n721), .Z(G69) );
  XNOR2_X1 U776 ( .A(G227), .B(KEYINPUT126), .ZN(n730) );
  XNOR2_X1 U777 ( .A(n724), .B(n723), .ZN(n727) );
  XOR2_X1 U778 ( .A(KEYINPUT125), .B(n725), .Z(n726) );
  XNOR2_X1 U779 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n729), .B(n728), .ZN(n734) );
  XNOR2_X1 U781 ( .A(n730), .B(n734), .ZN(n731) );
  NAND2_X1 U782 ( .A1(n731), .A2(G900), .ZN(n732) );
  NAND2_X1 U783 ( .A1(n732), .A2(G953), .ZN(n738) );
  XOR2_X1 U784 ( .A(n734), .B(n733), .Z(n736) );
  NAND2_X1 U785 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U786 ( .A1(n738), .A2(n737), .ZN(G72) );
  XNOR2_X1 U787 ( .A(G137), .B(n739), .ZN(G39) );
  XOR2_X1 U788 ( .A(n740), .B(G119), .Z(G21) );
  XNOR2_X1 U789 ( .A(G140), .B(KEYINPUT118), .ZN(n742) );
  XNOR2_X1 U790 ( .A(n742), .B(n741), .ZN(G42) );
endmodule

