//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT74), .B(G902), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT84), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  OR2_X1    g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT64), .A2(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT64), .A2(G146), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n193), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n198), .A2(G143), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n195), .A2(new_n196), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G143), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n202), .B1(new_n205), .B2(new_n191), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n198), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT64), .A2(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(G143), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n203), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n210), .A2(new_n202), .A3(new_n211), .A4(new_n191), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n201), .B1(new_n206), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  INV_X1    g031(.A(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT83), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(KEYINPUT4), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n222), .B1(new_n221), .B2(new_n224), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n221), .A2(G101), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n216), .A2(new_n219), .A3(new_n223), .A4(new_n220), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT4), .ZN(new_n229));
  OAI22_X1  g043(.A1(new_n225), .A2(new_n226), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n190), .B1(new_n214), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n210), .A2(new_n211), .A3(new_n191), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n200), .B1(new_n233), .B2(new_n212), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n221), .A2(new_n224), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT83), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n221), .A2(G101), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT4), .A3(new_n228), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n234), .A2(KEYINPUT84), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n231), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n243));
  INV_X1    g057(.A(G137), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(G134), .ZN(new_n245));
  INV_X1    g059(.A(G134), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT67), .A3(G137), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(KEYINPUT66), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G137), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT11), .A2(G134), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n246), .B2(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G131), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n248), .A2(new_n253), .A3(new_n258), .A4(new_n255), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(KEYINPUT1), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n210), .A2(new_n211), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n197), .A2(new_n199), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n262), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n215), .A2(G107), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n218), .A2(G104), .ZN(new_n270));
  OAI21_X1  g084(.A(G101), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n228), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n268), .A2(KEYINPUT10), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT10), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n262), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n264), .B1(new_n205), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n277), .A2(new_n278), .A3(new_n273), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n278), .B1(new_n277), .B2(new_n273), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n275), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n242), .A2(new_n261), .A3(new_n274), .A4(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT69), .B(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G227), .ZN(new_n284));
  XOR2_X1   g098(.A(G110), .B(G140), .Z(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n264), .B(new_n272), .C1(new_n266), .C2(new_n267), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n279), .B2(new_n280), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n290), .A2(KEYINPUT12), .A3(new_n260), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT12), .B1(new_n290), .B2(new_n260), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n231), .A2(new_n241), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n281), .A2(new_n274), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n260), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n287), .B1(new_n297), .B2(new_n282), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n187), .B(new_n189), .C1(new_n294), .C2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n282), .B1(new_n291), .B2(new_n292), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n286), .B(KEYINPUT82), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n282), .A2(new_n303), .A3(new_n287), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n297), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n303), .B1(new_n282), .B2(new_n287), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n302), .B(G469), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(G469), .A2(G902), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n299), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT9), .B(G234), .Z(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT81), .ZN(new_n311));
  OAI21_X1  g125(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G214), .B1(G237), .B2(G902), .ZN(new_n314));
  OAI21_X1  g128(.A(G210), .B1(G237), .B2(G902), .ZN(new_n315));
  XOR2_X1   g129(.A(G116), .B(G119), .Z(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT2), .B(G113), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n318), .B(new_n240), .C1(new_n225), .C2(new_n226), .ZN(new_n319));
  OR2_X1    g133(.A1(new_n316), .A2(new_n317), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT5), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT87), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT87), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT5), .ZN(new_n324));
  INV_X1    g138(.A(G119), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n322), .A2(new_n324), .A3(G116), .A4(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT87), .B(KEYINPUT5), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(G113), .C1(new_n316), .C2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n273), .A2(new_n320), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n319), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(G110), .B(G122), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n319), .A2(new_n331), .A3(new_n329), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(KEYINPUT6), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT88), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT76), .B(G125), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n338), .B(new_n264), .C1(new_n266), .C2(new_n267), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n336), .B(new_n339), .C1(new_n234), .C2(new_n338), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n214), .A2(KEYINPUT88), .A3(new_n337), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G953), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G224), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n344), .B(KEYINPUT89), .Z(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n340), .A2(new_n341), .A3(new_n345), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n330), .A2(new_n349), .A3(new_n332), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n335), .A2(new_n347), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT90), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n340), .A2(new_n341), .A3(new_n345), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n345), .B1(new_n340), .B2(new_n341), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT90), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n355), .A2(new_n356), .A3(new_n350), .A4(new_n335), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G902), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n345), .A2(KEYINPUT7), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n340), .A2(new_n341), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n331), .B(KEYINPUT8), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n326), .B(G113), .C1(new_n316), .C2(new_n321), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n273), .A2(new_n363), .A3(new_n320), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n328), .A2(new_n320), .B1(new_n228), .B2(new_n271), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT91), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n328), .A2(new_n320), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n368), .A2(new_n366), .A3(new_n272), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n362), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n361), .A2(new_n370), .A3(new_n334), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n360), .B1(new_n340), .B2(new_n341), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n359), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n315), .B1(new_n358), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n315), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n376), .B(new_n373), .C1(new_n352), .C2(new_n357), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n314), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(G116), .B(G122), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT97), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n218), .ZN(new_n381));
  INV_X1    g195(.A(G116), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT14), .A3(G122), .ZN(new_n383));
  INV_X1    g197(.A(new_n379), .ZN(new_n384));
  OAI211_X1 g198(.A(G107), .B(new_n383), .C1(new_n384), .C2(KEYINPUT14), .ZN(new_n385));
  XNOR2_X1  g199(.A(G128), .B(G143), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(new_n246), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT98), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n381), .A2(KEYINPUT98), .A3(new_n385), .A4(new_n387), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n380), .B(new_n218), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT13), .B1(new_n262), .B2(G143), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(new_n246), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n386), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G217), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n311), .A2(new_n398), .A3(G953), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n392), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n399), .B1(new_n392), .B2(new_n397), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n189), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G478), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT15), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n343), .A2(G952), .ZN(new_n406));
  INV_X1    g220(.A(G234), .ZN(new_n407));
  INV_X1    g221(.A(G237), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n283), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n411), .B(new_n188), .C1(new_n407), .C2(new_n408), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(KEYINPUT99), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT21), .B(G898), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  OAI221_X1 g230(.A(new_n189), .B1(KEYINPUT15), .B2(new_n403), .C1(new_n400), .C2(new_n401), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n405), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT20), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n343), .A2(KEYINPUT69), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT69), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G953), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n420), .A2(new_n422), .A3(G214), .A4(new_n408), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n194), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n283), .A2(G143), .A3(G214), .A4(new_n408), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(KEYINPUT18), .A2(G131), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G125), .B(G140), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n204), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT77), .ZN(new_n431));
  INV_X1    g245(.A(G140), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(G125), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n337), .B2(new_n432), .ZN(new_n434));
  OR2_X1    g248(.A1(KEYINPUT76), .A2(G125), .ZN(new_n435));
  NAND2_X1  g249(.A1(KEYINPUT76), .A2(G125), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n435), .A2(new_n431), .A3(G140), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n430), .B1(new_n438), .B2(new_n198), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n426), .A2(new_n427), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n428), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(KEYINPUT16), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n338), .A2(KEYINPUT16), .A3(G140), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(G146), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n204), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n434), .A2(KEYINPUT19), .A3(new_n437), .ZN(new_n447));
  INV_X1    g261(.A(new_n429), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(KEYINPUT19), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n445), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n426), .A2(G131), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n424), .A2(new_n425), .A3(new_n258), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n441), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G113), .B(G122), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(G104), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(KEYINPUT92), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT17), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n451), .A2(new_n459), .A3(new_n452), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT16), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(new_n434), .B2(new_n437), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n198), .B1(new_n462), .B2(new_n443), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n445), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n426), .A2(KEYINPUT17), .A3(G131), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT93), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n426), .A2(KEYINPUT93), .A3(KEYINPUT17), .A4(G131), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n441), .B(new_n458), .C1(new_n464), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n457), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(G475), .A2(G902), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n419), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n419), .A3(new_n472), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n470), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n441), .B1(new_n464), .B2(new_n469), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT95), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT95), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n480), .B(new_n441), .C1(new_n464), .C2(new_n469), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n456), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT96), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n477), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n479), .A2(KEYINPUT96), .A3(new_n456), .A4(new_n481), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(KEYINPUT94), .B(G475), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n418), .B(new_n476), .C1(new_n486), .C2(new_n488), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n313), .A2(new_n378), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT22), .B(G137), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT78), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n493), .B(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT23), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n325), .B2(G128), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n262), .A2(KEYINPUT23), .A3(G119), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n325), .A2(G128), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n500), .A2(KEYINPUT75), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(KEYINPUT75), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n502), .A3(G110), .ZN(new_n503));
  XOR2_X1   g317(.A(KEYINPUT24), .B(G110), .Z(new_n504));
  XNOR2_X1  g318(.A(G119), .B(G128), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n445), .B2(new_n463), .ZN(new_n508));
  OAI22_X1  g322(.A1(new_n500), .A2(G110), .B1(new_n504), .B2(new_n505), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n509), .A2(new_n430), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n445), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n495), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n445), .A2(new_n463), .ZN(new_n513));
  INV_X1    g327(.A(new_n507), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n445), .A2(new_n430), .A3(new_n509), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n493), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n517), .A3(new_n189), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT79), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT25), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n398), .B1(new_n189), .B2(G234), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n518), .A2(new_n520), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n512), .A2(new_n517), .A3(KEYINPUT25), .A4(new_n189), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(KEYINPUT79), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n512), .A2(new_n517), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n522), .A2(G902), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT80), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n531), .A2(KEYINPUT80), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n535));
  AOI21_X1  g349(.A(G134), .B1(new_n249), .B2(new_n251), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n246), .A2(G137), .ZN(new_n537));
  OAI21_X1  g351(.A(G131), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n259), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT68), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n259), .A3(KEYINPUT68), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n268), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n318), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n234), .A2(new_n260), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n283), .A2(G210), .A3(new_n408), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT71), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT26), .B(G101), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n550), .B(new_n553), .Z(new_n554));
  NAND3_X1  g368(.A1(new_n268), .A2(new_n259), .A3(new_n538), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n545), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n318), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n543), .A2(KEYINPUT28), .A3(new_n545), .A4(new_n544), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n548), .A2(new_n554), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n546), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT30), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n545), .A2(new_n561), .A3(new_n555), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n543), .A2(new_n545), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n562), .B1(new_n563), .B2(new_n561), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n564), .B2(new_n318), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n535), .B(new_n559), .C1(new_n565), .C2(new_n554), .ZN(new_n566));
  INV_X1    g380(.A(new_n554), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(new_n535), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT28), .B1(new_n560), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT73), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n546), .A2(new_n572), .A3(new_n547), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n568), .A2(new_n570), .A3(new_n571), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n566), .A2(new_n189), .A3(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n545), .A2(new_n561), .A3(new_n555), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n561), .B1(new_n543), .B2(new_n545), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n318), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n546), .A3(new_n554), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT31), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT31), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n578), .A2(new_n581), .A3(new_n546), .A4(new_n554), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n548), .A2(new_n557), .A3(new_n558), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n583), .A2(KEYINPUT72), .A3(new_n567), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT72), .B1(new_n583), .B2(new_n567), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n580), .B(new_n582), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT32), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n587), .A2(G472), .A3(G902), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n575), .A2(G472), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(G472), .A2(G902), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n587), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n534), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n490), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  INV_X1    g409(.A(G472), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n586), .B2(new_n189), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(KEYINPUT100), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n599));
  AOI211_X1 g413(.A(new_n599), .B(new_n596), .C1(new_n586), .C2(new_n189), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n586), .A2(new_n590), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n476), .B1(new_n486), .B2(new_n488), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n606), .B(new_n607), .C1(new_n400), .C2(new_n401), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n392), .A2(new_n397), .ZN(new_n609));
  INV_X1    g423(.A(new_n399), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n392), .A2(new_n397), .A3(new_n399), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n611), .A2(new_n604), .A3(new_n605), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n188), .A2(new_n403), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT102), .B(G478), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n402), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n617), .B1(new_n402), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n616), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n603), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n314), .B(new_n416), .C1(new_n375), .C2(new_n377), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n313), .A2(new_n534), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n602), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT34), .B(G104), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT104), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n627), .B(new_n629), .ZN(G6));
  NAND2_X1  g444(.A1(new_n405), .A2(new_n417), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n631), .B(new_n476), .C1(new_n486), .C2(new_n488), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n597), .A2(KEYINPUT100), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n601), .B1(KEYINPUT100), .B2(new_n597), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n633), .A2(new_n626), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NAND2_X1  g452(.A1(new_n515), .A2(new_n516), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n495), .A2(KEYINPUT36), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n523), .A2(new_n526), .B1(new_n530), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n602), .A2(new_n490), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G12));
  AOI21_X1  g460(.A(new_n642), .B1(new_n589), .B2(new_n592), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n313), .A2(new_n378), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT105), .B(G900), .Z(new_n649));
  AOI21_X1  g463(.A(new_n410), .B1(new_n413), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n632), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n647), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  AND2_X1   g467(.A1(new_n309), .A2(new_n312), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n650), .B(KEYINPUT39), .Z(new_n656));
  NAND3_X1  g470(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n655), .B1(new_n654), .B2(new_n656), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT40), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n659), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n662), .A3(new_n657), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n586), .A2(new_n588), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n565), .A2(new_n567), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n560), .A2(new_n569), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n359), .B1(new_n666), .B2(new_n554), .ZN(new_n667));
  OAI21_X1  g481(.A(G472), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n592), .A2(new_n664), .A3(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n642), .A2(new_n314), .A3(new_n631), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n603), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n375), .A2(new_n377), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT38), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n660), .A2(new_n663), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  INV_X1    g490(.A(new_n650), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n482), .A2(new_n483), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(new_n470), .A3(new_n485), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n488), .B1(new_n679), .B2(new_n359), .ZN(new_n680));
  INV_X1    g494(.A(new_n475), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n473), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n622), .B(new_n677), .C1(new_n680), .C2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n648), .A2(new_n647), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  INV_X1    g500(.A(new_n312), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n189), .B1(new_n294), .B2(new_n298), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G469), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(KEYINPUT107), .A3(new_n299), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n688), .A2(new_n691), .A3(G469), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n687), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n625), .A2(new_n593), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NAND3_X1  g510(.A1(new_n633), .A2(new_n593), .A3(new_n693), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  INV_X1    g512(.A(new_n378), .ZN(new_n699));
  INV_X1    g513(.A(new_n489), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n647), .A2(new_n693), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  OAI211_X1 g516(.A(new_n314), .B(new_n631), .C1(new_n375), .C2(new_n377), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n679), .A2(new_n359), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n682), .B1(new_n704), .B2(new_n487), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n590), .B(KEYINPUT108), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n580), .A2(new_n582), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT109), .A4(new_n573), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n567), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n707), .B1(new_n708), .B2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n534), .A2(new_n714), .A3(new_n597), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n706), .A2(new_n715), .A3(new_n693), .A4(new_n416), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G122), .ZN(G24));
  NOR3_X1   g531(.A1(new_n714), .A2(new_n597), .A3(new_n642), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n684), .A2(new_n693), .A3(new_n718), .A4(new_n699), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NAND2_X1  g534(.A1(new_n358), .A2(new_n374), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n376), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n358), .A2(new_n315), .A3(new_n374), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n314), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n313), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n593), .A3(new_n684), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n725), .A2(new_n593), .A3(new_n684), .A4(KEYINPUT42), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT110), .B(G131), .Z(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G33));
  NAND3_X1  g546(.A1(new_n725), .A2(new_n593), .A3(new_n651), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  NAND2_X1  g548(.A1(new_n635), .A2(new_n634), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n643), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n705), .A2(new_n622), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT43), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n705), .A2(new_n739), .A3(new_n622), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n724), .B1(new_n742), .B2(KEYINPUT44), .ZN(new_n743));
  INV_X1    g557(.A(new_n299), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n187), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n748));
  OAI22_X1  g562(.A1(new_n747), .A2(new_n748), .B1(new_n746), .B2(new_n745), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n308), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n744), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n749), .A2(new_n750), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n308), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n687), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n736), .B2(new_n741), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n743), .A2(new_n656), .A3(new_n756), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  INV_X1    g574(.A(new_n314), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n375), .A2(new_n377), .A3(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n762), .A2(new_n592), .A3(new_n589), .A4(new_n534), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n683), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n756), .A2(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n756), .A2(KEYINPUT47), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n432), .ZN(G42));
  NAND2_X1  g583(.A1(new_n690), .A2(new_n692), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT49), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n669), .A2(new_n761), .A3(new_n687), .A4(new_n534), .ZN(new_n772));
  INV_X1    g586(.A(new_n737), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n673), .A4(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n719), .A2(new_n652), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n299), .A2(new_n307), .A3(new_n308), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n641), .A2(new_n530), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n312), .B1(new_n677), .B2(KEYINPUT113), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(KEYINPUT113), .B2(new_n677), .ZN(new_n779));
  INV_X1    g593(.A(new_n526), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n521), .A2(new_n522), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n777), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT114), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n309), .A2(new_n642), .A3(new_n784), .A4(new_n779), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n706), .A2(new_n669), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n786), .A2(new_n685), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n775), .A2(new_n787), .A3(KEYINPUT115), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n719), .A2(new_n786), .A3(new_n685), .A4(new_n652), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n594), .A2(new_n644), .A3(new_n627), .A4(new_n636), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n694), .A2(new_n716), .A3(new_n701), .A4(new_n697), .ZN(new_n794));
  INV_X1    g608(.A(new_n733), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n728), .B2(new_n729), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n603), .A2(new_n631), .A3(new_n650), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n725), .A2(new_n647), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n725), .A2(new_n684), .A3(new_n718), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n725), .A2(new_n684), .A3(new_n718), .A4(KEYINPUT112), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n793), .A2(new_n794), .A3(new_n796), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n792), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n788), .A2(KEYINPUT52), .A3(new_n791), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(KEYINPUT53), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n789), .A2(KEYINPUT52), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n792), .A2(new_n804), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n807), .B1(KEYINPUT53), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT54), .ZN(new_n812));
  INV_X1    g626(.A(new_n804), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n788), .A2(new_n791), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n813), .A2(new_n816), .A3(KEYINPUT53), .A4(new_n808), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n818));
  INV_X1    g632(.A(new_n806), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n792), .A3(new_n804), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n817), .B(new_n818), .C1(new_n820), .C2(KEYINPUT53), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n812), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n715), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n741), .B2(new_n409), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n738), .A2(KEYINPUT116), .A3(new_n410), .A4(new_n740), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n673), .A2(new_n761), .A3(new_n693), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(KEYINPUT50), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n829), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n693), .A2(new_n762), .ZN(new_n833));
  OR4_X1    g647(.A1(new_n409), .A2(new_n833), .A3(new_n534), .A4(new_n669), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n834), .A2(new_n603), .A3(new_n622), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n833), .B1(new_n825), .B2(new_n826), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n835), .B1(new_n836), .B2(new_n718), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n770), .A2(new_n687), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n766), .A2(new_n767), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n762), .A3(new_n827), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT51), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n832), .A3(KEYINPUT51), .A4(new_n837), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n827), .A2(new_n699), .A3(new_n693), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n844), .B(new_n406), .C1(new_n623), .C2(new_n834), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n836), .A2(new_n593), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n846), .A2(KEYINPUT48), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(KEYINPUT48), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n822), .A2(new_n842), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(G952), .A2(G953), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n774), .B1(new_n851), .B2(new_n852), .ZN(G75));
  NOR2_X1   g667(.A1(new_n283), .A2(G952), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n813), .A2(new_n816), .A3(new_n806), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n189), .B1(new_n858), .B2(new_n817), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT56), .B1(new_n859), .B2(new_n376), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n335), .A2(new_n350), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(new_n355), .ZN(new_n862));
  XNOR2_X1  g676(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n855), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT53), .B1(new_n805), .B2(new_n806), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n792), .A2(new_n804), .A3(new_n857), .A4(new_n809), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n188), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT119), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n870), .B(new_n188), .C1(new_n866), .C2(new_n867), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n376), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT56), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n865), .B1(new_n872), .B2(new_n874), .ZN(G51));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n866), .B2(new_n867), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(KEYINPUT120), .A3(new_n821), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n878), .B(KEYINPUT54), .C1(new_n866), .C2(new_n867), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n308), .B(KEYINPUT57), .Z(new_n880));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n294), .A2(new_n298), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n754), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n869), .A2(new_n884), .A3(new_n871), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n854), .B1(new_n883), .B2(new_n885), .ZN(G54));
  AND2_X1   g700(.A1(KEYINPUT58), .A2(G475), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n869), .A2(new_n871), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n471), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n869), .A2(new_n471), .A3(new_n871), .A4(new_n887), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n890), .A2(new_n855), .A3(new_n891), .ZN(G60));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT59), .Z(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n812), .B2(new_n821), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n855), .B1(new_n895), .B2(new_n614), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n894), .B1(new_n608), .B2(new_n613), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n877), .A2(new_n879), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(new_n898), .ZN(G63));
  XNOR2_X1  g713(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n398), .A2(new_n359), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n900), .B(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n858), .B2(new_n817), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n641), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n905), .B(new_n855), .C1(new_n529), .C2(new_n904), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n904), .A2(new_n529), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(KEYINPUT61), .A3(new_n855), .A4(new_n905), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(G66));
  NAND2_X1  g725(.A1(new_n793), .A2(new_n794), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n283), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT122), .Z(new_n914));
  INV_X1    g728(.A(G224), .ZN(new_n915));
  OAI21_X1  g729(.A(G953), .B1(new_n414), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n861), .B1(G898), .B2(new_n283), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(G69));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n658), .A2(new_n659), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n623), .A2(new_n632), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(KEYINPUT124), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n593), .A2(new_n762), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n623), .A2(KEYINPUT124), .A3(new_n632), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n921), .A2(new_n923), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n719), .A2(new_n652), .A3(new_n685), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n675), .A2(KEYINPUT62), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT62), .B1(new_n675), .B2(new_n927), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n759), .B(new_n926), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n283), .B1(new_n930), .B2(new_n768), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n564), .B(KEYINPUT123), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(new_n449), .Z(new_n933));
  AOI21_X1  g747(.A(new_n920), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n283), .B1(G227), .B2(G900), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n796), .A2(new_n927), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n756), .A2(new_n656), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n706), .A2(new_n593), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n759), .B(new_n936), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n283), .B1(new_n939), .B2(new_n768), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n283), .A2(G900), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(KEYINPUT126), .A3(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n933), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT126), .B1(new_n940), .B2(new_n942), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n934), .B(new_n935), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n940), .A2(new_n942), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n944), .A3(new_n943), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n935), .B1(new_n952), .B2(new_n934), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n948), .A2(new_n953), .ZN(G72));
  AND2_X1   g768(.A1(new_n565), .A2(new_n567), .ZN(new_n955));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT63), .Z(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n955), .A2(new_n665), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n811), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT127), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n930), .A2(new_n768), .A3(new_n912), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n665), .B1(new_n962), .B2(new_n958), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n939), .A2(new_n768), .A3(new_n912), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n955), .B1(new_n964), .B2(new_n958), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n963), .A2(new_n965), .A3(new_n855), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n961), .A2(new_n966), .ZN(G57));
endmodule


