//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1226, new_n1227, new_n1228, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(new_n203), .A2(G50), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  AND2_X1   g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n213), .B1(new_n214), .B2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G13), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n216), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT0), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n212), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(new_n220), .B2(new_n219), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT65), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n214), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n223), .A2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  OR2_X1    g0048(.A1(KEYINPUT67), .A2(G1), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT67), .A2(G1), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n249), .A2(G13), .A3(G20), .A4(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G97), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g0057(.A1(KEYINPUT68), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n257), .A2(new_n209), .A3(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT67), .A2(G1), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT67), .A2(G1), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n259), .A2(new_n251), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n254), .B1(new_n264), .B2(new_n253), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT79), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n257), .A2(new_n209), .A3(new_n258), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT6), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n269), .A2(G97), .A3(G107), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n253), .A2(KEYINPUT6), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT78), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G107), .ZN(new_n273));
  INV_X1    g0073(.A(G107), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(KEYINPUT78), .ZN(new_n275));
  OAI22_X1  g0075(.A1(new_n270), .A2(new_n271), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G97), .A2(G107), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT6), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n269), .A2(G97), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n274), .A2(KEYINPUT78), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n272), .A2(G107), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n278), .A2(new_n279), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n276), .A2(G20), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G77), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT7), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT3), .B(G33), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(G20), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n274), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n267), .B(new_n268), .C1(new_n286), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n288), .A2(new_n287), .A3(G20), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT7), .B1(new_n292), .B2(new_n210), .ZN(new_n298));
  OAI21_X1  g0098(.A(G107), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(new_n285), .A3(new_n283), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n267), .B1(new_n300), .B2(new_n268), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n266), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G41), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G1), .A3(G13), .ZN(new_n305));
  INV_X1    g0105(.A(G1698), .ZN(new_n306));
  OAI211_X1 g0106(.A(G244), .B(new_n306), .C1(new_n290), .C2(new_n291), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT4), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT4), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n288), .A2(new_n309), .A3(G244), .A4(new_n306), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(KEYINPUT3), .A2(G33), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n306), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n314), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT80), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT80), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n311), .A2(new_n318), .A3(new_n315), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n305), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n249), .A2(G45), .A3(new_n250), .ZN(new_n321));
  INV_X1    g0121(.A(G41), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT5), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT5), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G41), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(G257), .B(new_n305), .C1(new_n321), .C2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G274), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n208), .B2(new_n304), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT5), .B(G41), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n329), .A2(new_n262), .A3(new_n330), .A4(G45), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n303), .B1(new_n320), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n305), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n311), .A2(new_n318), .A3(new_n315), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n318), .B1(new_n311), .B2(new_n315), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n332), .A2(KEYINPUT81), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT81), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n327), .A2(new_n339), .A3(new_n331), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G179), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n337), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n302), .A2(new_n333), .A3(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(G200), .B1(new_n320), .B2(new_n341), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n268), .B1(new_n286), .B2(new_n294), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT79), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n265), .B1(new_n348), .B2(new_n295), .ZN(new_n349));
  INV_X1    g0149(.A(new_n332), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n337), .A2(G190), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n346), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT12), .B1(new_n252), .B2(new_n202), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n252), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n249), .A2(new_n250), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(new_n210), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n268), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n354), .B(new_n355), .C1(G68), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n210), .A2(G33), .ZN(new_n360));
  INV_X1    g0160(.A(G77), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n360), .A2(new_n361), .B1(new_n210), .B2(G68), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT72), .ZN(new_n363));
  INV_X1    g0163(.A(G50), .ZN(new_n364));
  INV_X1    g0164(.A(new_n284), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n362), .A2(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n362), .A2(new_n363), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n268), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT11), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n368), .A2(new_n369), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n359), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(G226), .A2(G1698), .ZN(new_n374));
  INV_X1    g0174(.A(G232), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(G1698), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n288), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G97), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(KEYINPUT71), .A3(new_n334), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT71), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n376), .A2(new_n288), .B1(G33), .B2(G97), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n305), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT13), .ZN(new_n385));
  INV_X1    g0185(.A(G1), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G41), .A2(G45), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n329), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n262), .A2(new_n388), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n305), .ZN(new_n391));
  INV_X1    g0191(.A(G238), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n384), .A2(new_n385), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n385), .B1(new_n384), .B2(new_n394), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT73), .B(G169), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n396), .A2(new_n397), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n398), .A2(KEYINPUT14), .B1(new_n399), .B2(G179), .ZN(new_n400));
  NAND2_X1  g0200(.A1(KEYINPUT73), .A2(G169), .ZN(new_n401));
  INV_X1    g0201(.A(new_n397), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n401), .B1(new_n402), .B2(new_n395), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT14), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n373), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n399), .A2(G190), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(new_n395), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G200), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(new_n409), .A3(new_n373), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n406), .A2(new_n411), .A3(KEYINPUT74), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT74), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n403), .A2(new_n404), .B1(new_n408), .B2(new_n343), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n398), .A2(KEYINPUT14), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n372), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n413), .B1(new_n416), .B2(new_n410), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n252), .A2(new_n361), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT70), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n358), .A2(G77), .ZN(new_n420));
  XNOR2_X1  g0220(.A(KEYINPUT8), .B(G58), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n421), .A2(new_n365), .B1(new_n210), .B2(new_n361), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT15), .B(G87), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n423), .A2(new_n360), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n268), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n419), .A2(new_n420), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n314), .A2(G238), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n288), .A2(new_n306), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n427), .B1(new_n274), .B2(new_n288), .C1(new_n375), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n334), .ZN(new_n430));
  INV_X1    g0230(.A(new_n391), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G244), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n389), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n426), .B1(G200), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G190), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(new_n433), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n303), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n430), .A2(new_n343), .A3(new_n389), .A4(new_n432), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(new_n426), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G226), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n389), .B1(new_n391), .B2(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n314), .A2(G223), .B1(new_n292), .B2(G77), .ZN(new_n443));
  INV_X1    g0243(.A(G222), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(new_n428), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n442), .B1(new_n445), .B2(new_n334), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n343), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(G169), .B2(new_n446), .ZN(new_n448));
  INV_X1    g0248(.A(G150), .ZN(new_n449));
  OAI22_X1  g0249(.A1(new_n421), .A2(new_n360), .B1(new_n449), .B2(new_n365), .ZN(new_n450));
  INV_X1    g0250(.A(new_n203), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n210), .B1(new_n451), .B2(new_n364), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n268), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(G50), .B1(new_n357), .B2(new_n268), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n251), .A2(new_n364), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n454), .A2(KEYINPUT69), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT69), .B1(new_n454), .B2(new_n455), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n453), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n448), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n458), .B(KEYINPUT9), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT10), .ZN(new_n463));
  INV_X1    g0263(.A(G200), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n446), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(G190), .B2(new_n446), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n463), .B1(new_n462), .B2(new_n466), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n440), .B(new_n461), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n412), .A2(new_n417), .A3(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n259), .A2(G116), .A3(new_n251), .A4(new_n263), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n252), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(G20), .B1(G33), .B2(G283), .ZN(new_n475));
  INV_X1    g0275(.A(G33), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G97), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n475), .A2(new_n477), .B1(G20), .B2(new_n473), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n268), .A2(KEYINPUT20), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT20), .B1(new_n268), .B2(new_n478), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n472), .B(new_n474), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n288), .A2(G264), .A3(G1698), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n288), .A2(G257), .A3(new_n306), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n292), .A2(G303), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n262), .A2(new_n330), .A3(G45), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n485), .A2(new_n334), .B1(new_n487), .B2(new_n329), .ZN(new_n488));
  OAI211_X1 g0288(.A(G270), .B(new_n305), .C1(new_n321), .C2(new_n326), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n486), .A2(new_n491), .A3(G270), .A4(new_n305), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n481), .B1(new_n494), .B2(G200), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n435), .B2(new_n494), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(G169), .A3(new_n481), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT21), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n494), .A2(new_n343), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n481), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n494), .A2(new_n481), .A3(KEYINPUT21), .A4(G169), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n496), .A2(new_n499), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT19), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n210), .B1(new_n378), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(G87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n277), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n210), .B(G68), .C1(new_n290), .C2(new_n291), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n504), .B1(new_n360), .B2(new_n253), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n268), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n252), .A2(new_n423), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n264), .A2(new_n423), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n321), .A2(G250), .A3(new_n305), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n329), .A2(G45), .A3(new_n262), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G244), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n519));
  OAI211_X1 g0319(.A(G238), .B(new_n306), .C1(new_n290), .C2(new_n291), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G116), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n518), .B1(new_n334), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n514), .A2(new_n515), .B1(new_n523), .B2(new_n343), .ZN(new_n524));
  INV_X1    g0324(.A(new_n518), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n522), .A2(new_n334), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n303), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n259), .A2(G87), .A3(new_n251), .A4(new_n263), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n512), .A2(new_n529), .A3(new_n513), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(G190), .B2(new_n523), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(G200), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n524), .A2(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT23), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n521), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n534), .A2(KEYINPUT84), .B1(new_n536), .B2(new_n210), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n274), .A3(G20), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT84), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n538), .A2(new_n539), .B1(KEYINPUT23), .B2(G107), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT22), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(KEYINPUT83), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n288), .A2(new_n210), .A3(G87), .A4(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n210), .B(G87), .C1(new_n290), .C2(new_n291), .ZN(new_n546));
  XNOR2_X1  g0346(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n541), .A2(new_n542), .A3(new_n545), .A4(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n548), .A2(new_n545), .A3(new_n537), .A4(new_n540), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT24), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n259), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g0352(.A(KEYINPUT85), .B(KEYINPUT25), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n252), .A2(new_n274), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT85), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n555), .B(KEYINPUT25), .C1(new_n251), .C2(G107), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n554), .B(new_n556), .C1(new_n264), .C2(new_n274), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G257), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n559));
  OAI211_X1 g0359(.A(G250), .B(new_n306), .C1(new_n290), .C2(new_n291), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G294), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT86), .B1(new_n562), .B2(new_n334), .ZN(new_n563));
  OAI211_X1 g0363(.A(G264), .B(new_n305), .C1(new_n321), .C2(new_n326), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n331), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(KEYINPUT86), .A3(new_n334), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n435), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n562), .A2(new_n334), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n331), .A3(new_n564), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n464), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n558), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n303), .B1(new_n566), .B2(new_n567), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n570), .A2(new_n343), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n574), .A2(new_n575), .B1(new_n552), .B2(new_n557), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n533), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n503), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G68), .B1(new_n297), .B2(new_n298), .ZN(new_n579));
  XNOR2_X1  g0379(.A(G58), .B(G68), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(G20), .B1(G159), .B2(new_n284), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT16), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n579), .A2(KEYINPUT16), .A3(new_n581), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n268), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n421), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(new_n251), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n358), .B2(new_n587), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G232), .B(new_n305), .C1(new_n356), .C2(new_n387), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT75), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G223), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n306), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n441), .A2(G1698), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(new_n290), .C2(new_n291), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G87), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n334), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n390), .A2(KEYINPUT75), .A3(G232), .A4(new_n305), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n594), .A2(new_n601), .A3(new_n602), .A4(new_n389), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT76), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n386), .A2(new_n305), .A3(G274), .A4(new_n388), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n334), .B2(new_n600), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT76), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n602), .A4(new_n594), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n464), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n603), .A2(G190), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT77), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(G200), .B1(new_n604), .B2(new_n608), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT77), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n614), .A2(new_n615), .A3(new_n611), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n591), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT17), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n603), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n609), .A2(new_n303), .B1(new_n343), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT18), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n621), .A2(new_n622), .A3(new_n590), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(new_n621), .B2(new_n590), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n610), .A2(KEYINPUT77), .A3(new_n612), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n615), .B1(new_n614), .B2(new_n611), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n590), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT17), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n619), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n353), .A2(new_n471), .A3(new_n578), .A4(new_n631), .ZN(G372));
  NAND2_X1  g0432(.A1(new_n626), .A2(new_n627), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT17), .B1(new_n633), .B2(new_n591), .ZN(new_n634));
  AOI211_X1 g0434(.A(new_n618), .B(new_n590), .C1(new_n626), .C2(new_n627), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n439), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n410), .B1(new_n406), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n625), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n468), .A2(new_n469), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n460), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n471), .A2(new_n631), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n576), .A2(new_n499), .A3(new_n501), .A4(new_n502), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT87), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n522), .A2(new_n645), .A3(new_n334), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n645), .B1(new_n522), .B2(new_n334), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n525), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G200), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n558), .A2(new_n572), .B1(new_n531), .B2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n644), .A2(new_n345), .A3(new_n352), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n303), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n524), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n317), .A2(new_n319), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n341), .B1(new_n655), .B2(new_n334), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n337), .A2(new_n350), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n343), .A2(new_n656), .B1(new_n657), .B2(new_n303), .ZN(new_n658));
  XNOR2_X1  g0458(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n658), .A2(new_n302), .A3(new_n533), .A4(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n524), .A2(new_n652), .B1(new_n649), .B2(new_n531), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n663), .A2(new_n302), .A3(new_n344), .A4(new_n333), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n661), .A2(KEYINPUT89), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n302), .A2(new_n333), .A3(new_n344), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT89), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n533), .A4(new_n660), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n654), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n642), .B1(new_n643), .B2(new_n669), .ZN(G369));
  AND2_X1   g0470(.A1(new_n501), .A2(new_n502), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n499), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n216), .A2(G20), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n262), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n679), .A2(new_n481), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n672), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n503), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n573), .A2(new_n576), .ZN(new_n685));
  INV_X1    g0485(.A(new_n679), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n558), .A2(new_n686), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n685), .A2(new_n687), .B1(new_n576), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  AOI211_X1 g0489(.A(new_n679), .B(new_n685), .C1(new_n499), .C2(new_n671), .ZN(new_n690));
  INV_X1    g0490(.A(new_n576), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n686), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n218), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n694), .A2(KEYINPUT91), .A3(G41), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT91), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n218), .B2(new_n322), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n507), .A2(G116), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT90), .Z(new_n700));
  NOR3_X1   g0500(.A1(new_n698), .A2(new_n700), .A3(new_n386), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(new_n207), .B2(new_n698), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT28), .Z(new_n703));
  XNOR2_X1  g0503(.A(KEYINPUT94), .B(KEYINPUT30), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n523), .A2(new_n569), .A3(new_n564), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n500), .A2(new_n706), .A3(new_n337), .A4(new_n350), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT93), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n320), .A2(new_n332), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(KEYINPUT93), .A3(new_n500), .A4(new_n706), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n705), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  AND4_X1   g0512(.A1(new_n343), .A2(new_n648), .A3(new_n494), .A4(new_n570), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n337), .A2(new_n342), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n707), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n679), .B1(new_n712), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n578), .A2(new_n353), .A3(new_n686), .ZN(new_n721));
  XNOR2_X1  g0521(.A(KEYINPUT92), .B(KEYINPUT31), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n679), .B(new_n723), .C1(new_n712), .C2(new_n717), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n720), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT95), .B1(new_n669), .B2(new_n679), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT95), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n533), .A2(new_n302), .A3(new_n344), .A4(new_n333), .ZN(new_n729));
  OAI21_X1  g0529(.A(KEYINPUT89), .B1(new_n729), .B2(new_n659), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n664), .A2(new_n662), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n730), .A2(new_n668), .A3(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n728), .B(new_n686), .C1(new_n732), .C2(new_n654), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT29), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n664), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n736), .A2(KEYINPUT26), .B1(new_n729), .B2(new_n659), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT29), .B(new_n686), .C1(new_n737), .C2(new_n654), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n726), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n703), .B1(new_n739), .B2(G1), .ZN(G364));
  AOI21_X1  g0540(.A(new_n386), .B1(new_n673), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n698), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n684), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G330), .B2(new_n682), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n218), .A2(G355), .A3(new_n288), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G116), .B2(new_n218), .ZN(new_n747));
  INV_X1    g0547(.A(G45), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n244), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n218), .A2(new_n292), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n748), .B2(new_n207), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n747), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT96), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n209), .B1(G20), .B2(new_n303), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n743), .B1(new_n752), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(G20), .A2(G179), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT97), .Z(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G190), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n464), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n761), .A2(new_n435), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G200), .ZN(new_n765));
  AOI22_X1  g0565(.A1(G50), .A2(new_n763), .B1(new_n765), .B2(G77), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n762), .A2(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n764), .A2(new_n464), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n766), .B1(new_n201), .B2(new_n768), .C1(new_n202), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n210), .A2(G179), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(new_n435), .A3(new_n464), .ZN(new_n773));
  INV_X1    g0573(.A(G159), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT32), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n772), .A2(G190), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n292), .B1(new_n778), .B2(G87), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n435), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n210), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n772), .A2(new_n435), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n782), .A2(G97), .B1(new_n784), .B2(G107), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n776), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G311), .A2(new_n765), .B1(new_n763), .B2(G326), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n770), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G303), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n292), .B1(new_n777), .B2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT98), .Z(new_n792));
  NAND2_X1  g0592(.A1(new_n767), .A2(G322), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n784), .A2(G283), .ZN(new_n794));
  INV_X1    g0594(.A(new_n773), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n782), .A2(G294), .B1(new_n795), .B2(G329), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n792), .A2(new_n793), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n771), .A2(new_n786), .B1(new_n789), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n759), .B1(new_n798), .B2(new_n756), .ZN(new_n799));
  INV_X1    g0599(.A(new_n755), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n682), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n745), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n727), .A2(new_n733), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n426), .A2(new_n679), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n436), .A2(new_n439), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n437), .A2(new_n438), .A3(new_n426), .A4(new_n679), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT100), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT102), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n806), .B(KEYINPUT102), .C1(new_n810), .C2(new_n811), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n804), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n730), .A2(new_n668), .A3(new_n731), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n817), .A2(new_n653), .A3(new_n651), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n812), .A2(new_n686), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n726), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n743), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n816), .A2(new_n726), .A3(new_n821), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n756), .A2(new_n753), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n743), .B1(G77), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n769), .A2(KEYINPUT99), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n769), .A2(KEYINPUT99), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G283), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n763), .A2(G303), .ZN(new_n833));
  INV_X1    g0633(.A(G311), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n292), .B1(new_n773), .B2(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n506), .A2(new_n783), .B1(new_n777), .B2(new_n274), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(G97), .C2(new_n782), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G116), .A2(new_n765), .B1(new_n767), .B2(G294), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n832), .A2(new_n833), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G143), .A2(new_n767), .B1(new_n765), .B2(G159), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  INV_X1    g0641(.A(new_n763), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n840), .B1(new_n841), .B2(new_n842), .C1(new_n449), .C2(new_n770), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT34), .Z(new_n844));
  AOI22_X1  g0644(.A1(new_n782), .A2(G58), .B1(new_n778), .B2(G50), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n292), .B1(new_n795), .B2(G132), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(new_n202), .C2(new_n783), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n839), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n827), .B1(new_n848), .B2(new_n756), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n754), .B2(new_n812), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT101), .Z(new_n851));
  NAND2_X1  g0651(.A1(new_n825), .A2(new_n851), .ZN(G384));
  NOR2_X1   g0652(.A1(new_n262), .A2(new_n673), .ZN(new_n853));
  INV_X1    g0653(.A(G330), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  INV_X1    g0655(.A(new_n677), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n590), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n636), .B2(new_n625), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n621), .A2(new_n590), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n857), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n628), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n590), .B1(new_n621), .B2(new_n856), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n617), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n855), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n857), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n630), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n812), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n372), .B(new_n679), .C1(new_n406), .C2(new_n411), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n372), .A2(new_n679), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n416), .A2(new_n410), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n872), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n718), .A2(new_n722), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n877), .B(new_n721), .C1(new_n719), .C2(new_n718), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT40), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n871), .A2(new_n879), .A3(KEYINPUT40), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT103), .Z(new_n885));
  AND3_X1   g0685(.A1(new_n471), .A2(new_n631), .A3(new_n878), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n854), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n886), .B2(new_n885), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT104), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n873), .A2(new_n875), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n439), .A2(new_n679), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n669), .B2(new_n819), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n871), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n625), .B2(new_n856), .ZN(new_n896));
  AOI221_X4 g0696(.A(new_n855), .B1(new_n861), .B2(new_n864), .C1(new_n630), .C2(new_n868), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n869), .B2(new_n865), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT39), .B1(new_n867), .B2(new_n870), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n406), .A2(new_n686), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n896), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n471), .A2(new_n631), .A3(new_n738), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n734), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n640), .A2(new_n641), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n907), .A2(new_n460), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n905), .B(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n853), .B1(new_n890), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n890), .B2(new_n910), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n276), .A2(new_n282), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT35), .ZN(new_n914));
  OAI211_X1 g0714(.A(G116), .B(new_n211), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n914), .B2(new_n913), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n916), .B(KEYINPUT36), .Z(new_n917));
  OAI21_X1  g0717(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n206), .A2(new_n918), .B1(G50), .B2(new_n202), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n216), .A3(new_n356), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n912), .A2(new_n917), .A3(new_n920), .ZN(G367));
  INV_X1    g0721(.A(new_n739), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n353), .B1(new_n349), .B2(new_n686), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n345), .B2(new_n686), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n692), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT107), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT107), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n692), .A2(new_n927), .A3(new_n924), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT45), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n692), .A2(new_n924), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT44), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n926), .A2(KEYINPUT45), .A3(new_n928), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT108), .ZN(new_n936));
  INV_X1    g0736(.A(new_n689), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n936), .B1(new_n935), .B2(new_n937), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n935), .A2(new_n937), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n690), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n679), .B1(new_n671), .B2(new_n499), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n942), .B1(new_n688), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(new_n684), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n922), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n698), .B(KEYINPUT41), .Z(new_n947));
  OAI21_X1  g0747(.A(new_n741), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n924), .A2(new_n690), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT42), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n345), .B1(new_n923), .B2(new_n576), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n686), .B1(new_n951), .B2(KEYINPUT106), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(KEYINPUT106), .B2(new_n951), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT43), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n679), .A2(new_n530), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n663), .A2(new_n955), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n956), .A2(KEYINPUT105), .B1(new_n653), .B2(new_n955), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(KEYINPUT105), .B2(new_n956), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n950), .A2(new_n953), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n954), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n937), .A2(new_n924), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n958), .A2(new_n755), .ZN(new_n964));
  INV_X1    g0764(.A(new_n743), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT109), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n757), .B1(new_n218), .B2(new_n423), .C1(new_n240), .C2(new_n750), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n966), .B2(new_n967), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n783), .A2(new_n253), .ZN(new_n970));
  INV_X1    g0770(.A(G317), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n292), .B1(new_n773), .B2(new_n971), .C1(new_n781), .C2(new_n274), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n778), .A2(KEYINPUT46), .A3(G116), .ZN(new_n973));
  AOI21_X1  g0773(.A(KEYINPUT46), .B1(new_n778), .B2(G116), .ZN(new_n974));
  OR4_X1    g0774(.A1(new_n970), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G283), .A2(new_n765), .B1(new_n763), .B2(G311), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n790), .B2(new_n768), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n975), .B(new_n977), .C1(G294), .C2(new_n831), .ZN(new_n978));
  INV_X1    g0778(.A(new_n765), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n830), .A2(new_n774), .B1(new_n364), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT110), .Z(new_n981));
  OAI22_X1  g0781(.A1(new_n773), .A2(new_n841), .B1(new_n777), .B2(new_n201), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT112), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n982), .A2(new_n983), .B1(G68), .B2(new_n782), .ZN(new_n984));
  INV_X1    g0784(.A(G143), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n984), .B1(new_n983), .B2(new_n982), .C1(new_n842), .C2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n288), .B1(new_n783), .B2(new_n361), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n767), .A2(G150), .B1(KEYINPUT111), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(KEYINPUT111), .B2(new_n987), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n978), .B1(new_n981), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n969), .B1(new_n993), .B2(new_n756), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n948), .A2(new_n963), .B1(new_n964), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(G387));
  NOR2_X1   g0796(.A1(new_n739), .A2(new_n945), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT115), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n739), .A2(new_n945), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(KEYINPUT115), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n998), .A2(new_n698), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n688), .A2(new_n800), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n237), .A2(new_n748), .A3(new_n288), .ZN(new_n1003));
  OR3_X1    g0803(.A1(new_n421), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT50), .B1(new_n421), .B2(G50), .ZN(new_n1005));
  AOI21_X1  g0805(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n700), .B1(new_n1007), .B2(new_n292), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n218), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1009), .B(new_n757), .C1(new_n274), .C2(new_n218), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n743), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n364), .A2(new_n768), .B1(new_n842), .B2(new_n774), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n587), .B2(new_n769), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n781), .A2(new_n423), .B1(new_n777), .B2(new_n361), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n288), .B1(new_n773), .B2(new_n449), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n1014), .A2(new_n970), .A3(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1013), .B(new_n1016), .C1(new_n202), .C2(new_n979), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n979), .A2(new_n790), .ZN(new_n1018));
  XOR2_X1   g0818(.A(KEYINPUT114), .B(G322), .Z(new_n1019));
  AOI21_X1  g0819(.A(new_n1018), .B1(new_n763), .B2(new_n1019), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n834), .B2(new_n830), .C1(new_n971), .C2(new_n768), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT48), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(G283), .ZN(new_n1024));
  INV_X1    g0824(.A(G294), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n781), .A2(new_n1024), .B1(new_n777), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1023), .A2(KEYINPUT49), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n288), .B1(new_n795), .B2(G326), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(new_n473), .C2(new_n783), .ZN(new_n1030));
  AOI21_X1  g0830(.A(KEYINPUT49), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1017), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1002), .B(new_n1011), .C1(new_n1032), .C2(new_n756), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n945), .B2(new_n742), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1001), .A2(new_n1034), .ZN(G393));
  AND2_X1   g0835(.A1(new_n935), .A2(new_n937), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n999), .B1(new_n1036), .B2(new_n940), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n939), .A2(new_n940), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n938), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1037), .B(new_n698), .C1(new_n1040), .C2(new_n999), .ZN(new_n1041));
  OR3_X1    g0841(.A1(new_n1036), .A2(new_n940), .A3(new_n741), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT116), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n757), .B1(new_n253), .B2(new_n218), .C1(new_n247), .C2(new_n750), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n965), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G150), .A2(new_n763), .B1(new_n767), .B2(G159), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT51), .Z(new_n1048));
  OAI22_X1  g0848(.A1(new_n781), .A2(new_n361), .B1(new_n777), .B2(new_n202), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n288), .B1(new_n773), .B2(new_n985), .C1(new_n506), .C2(new_n783), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n765), .C2(new_n587), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1048), .B(new_n1051), .C1(new_n364), .C2(new_n830), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G311), .A2(new_n767), .B1(new_n763), .B2(G317), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT117), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1054), .A2(KEYINPUT52), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(KEYINPUT52), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n288), .B1(new_n795), .B2(new_n1019), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n274), .B2(new_n783), .C1(new_n1024), .C2(new_n777), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G294), .B2(new_n765), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1055), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n830), .A2(new_n790), .B1(new_n473), .B2(new_n781), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT118), .Z(new_n1062));
  OAI21_X1  g0862(.A(new_n1052), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1046), .B1(new_n1063), .B2(new_n756), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n924), .B2(new_n800), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1041), .A2(new_n1042), .A3(new_n1065), .ZN(G390));
  INV_X1    g0866(.A(KEYINPUT122), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n471), .A2(new_n878), .A3(G330), .A4(new_n631), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n642), .B(new_n1068), .C1(new_n734), .C2(new_n906), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n725), .A2(G330), .A3(new_n812), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n873), .A2(new_n875), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n876), .A2(new_n878), .A3(G330), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n894), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n686), .B(new_n812), .C1(new_n737), .C2(new_n654), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1076), .A2(new_n893), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n891), .A2(new_n725), .A3(G330), .A4(new_n812), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n814), .A2(new_n815), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n878), .A2(G330), .A3(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1077), .B(new_n1078), .C1(new_n1080), .C2(new_n891), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1069), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n894), .A2(new_n891), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n903), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n900), .B2(new_n901), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n871), .B(new_n903), .C1(new_n1071), .C2(new_n1077), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n1086), .A3(new_n1078), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n904), .B1(new_n894), .B2(new_n891), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n870), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n903), .B1(new_n897), .B2(new_n898), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1076), .A2(new_n893), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1093), .A2(new_n891), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1074), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1082), .A2(new_n1087), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT119), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n1098), .A3(new_n698), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1087), .A2(new_n1096), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1082), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1098), .B1(new_n1097), .B2(new_n698), .ZN(new_n1104));
  OAI21_X1  g0904(.A(KEYINPUT120), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1097), .A2(new_n698), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(KEYINPUT119), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT120), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1107), .A2(new_n1108), .A3(new_n1102), .A4(new_n1099), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1087), .A2(new_n1096), .A3(new_n742), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n743), .B1(new_n587), .B2(new_n826), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n781), .A2(new_n361), .B1(new_n783), .B2(new_n202), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n292), .B1(new_n773), .B2(new_n1025), .C1(new_n506), .C2(new_n777), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(new_n767), .C2(G116), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G97), .A2(new_n765), .B1(new_n763), .B2(G283), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(new_n830), .C2(new_n274), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n765), .A2(new_n1119), .B1(G159), .B2(new_n782), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n830), .B2(new_n841), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT121), .Z(new_n1122));
  OAI21_X1  g0922(.A(KEYINPUT53), .B1(new_n777), .B2(new_n449), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n292), .B1(new_n795), .B2(G125), .ZN(new_n1124));
  OR3_X1    g0924(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n449), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n784), .A2(G50), .ZN(new_n1126));
  AND4_X1   g0926(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(G128), .ZN(new_n1128));
  INV_X1    g0928(.A(G132), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1127), .B1(new_n1128), .B2(new_n842), .C1(new_n1129), .C2(new_n768), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1117), .B1(new_n1122), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1112), .B1(new_n1131), .B2(new_n756), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n902), .B2(new_n754), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1111), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1067), .B1(new_n1110), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(KEYINPUT122), .B(new_n1134), .C1(new_n1105), .C2(new_n1109), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(G378));
  NOR2_X1   g0940(.A1(new_n459), .A2(new_n677), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n641), .B2(new_n461), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n641), .A2(new_n461), .A3(new_n1142), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1146), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n884), .B2(new_n854), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1150), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1152), .A2(new_n882), .A3(G330), .A4(new_n883), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n905), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1151), .A2(new_n905), .A3(new_n1153), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n742), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1152), .A2(new_n754), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n743), .B1(G50), .B2(new_n826), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n322), .B(new_n292), .C1(new_n773), .C2(new_n1024), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G68), .B2(new_n782), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n778), .A2(G77), .B1(new_n784), .B2(G58), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n768), .C2(new_n274), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n253), .A2(new_n770), .B1(new_n979), .B2(new_n423), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(G116), .C2(new_n763), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT58), .Z(new_n1168));
  AOI21_X1  g0968(.A(G50), .B1(new_n476), .B2(new_n322), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n288), .B2(G41), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n781), .A2(new_n449), .B1(new_n777), .B2(new_n1118), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G125), .A2(new_n763), .B1(new_n767), .B2(G128), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n841), .B2(new_n979), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(G132), .C2(new_n769), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n784), .A2(G159), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G33), .B(G41), .C1(new_n795), .C2(G124), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1168), .B(new_n1170), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1181), .A2(KEYINPUT123), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n756), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1181), .B2(KEYINPUT123), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1161), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1160), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1159), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n698), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1069), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1156), .A2(new_n1157), .B1(new_n1189), .B2(new_n1097), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1188), .B1(new_n1190), .B2(KEYINPUT57), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1097), .A2(new_n1189), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1158), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1187), .B1(new_n1191), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(G375));
  NAND2_X1  g0997(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1198));
  OR3_X1    g0998(.A1(new_n1198), .A2(KEYINPUT124), .A3(new_n1189), .ZN(new_n1199));
  OAI21_X1  g0999(.A(KEYINPUT124), .B1(new_n1198), .B2(new_n1189), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1082), .A2(new_n947), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1071), .A2(new_n753), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n743), .B1(G68), .B2(new_n826), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n781), .A2(new_n364), .B1(new_n777), .B2(new_n774), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n288), .B1(new_n773), .B2(new_n1128), .C1(new_n201), .C2(new_n783), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(new_n767), .C2(G137), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G132), .A2(new_n763), .B1(new_n765), .B2(G150), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n830), .C2(new_n1118), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n830), .A2(new_n473), .B1(new_n274), .B2(new_n979), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT125), .Z(new_n1211));
  NOR2_X1   g1011(.A1(new_n842), .A2(new_n1025), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n768), .A2(new_n1024), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n292), .B1(new_n773), .B2(new_n790), .C1(new_n361), .C2(new_n783), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n781), .A2(new_n423), .B1(new_n777), .B2(new_n253), .ZN(new_n1215));
  OR4_X1    g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1209), .B1(new_n1211), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1204), .B1(new_n1217), .B2(new_n756), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1198), .A2(new_n742), .B1(new_n1203), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1202), .A2(new_n1219), .ZN(G381));
  NAND3_X1  g1020(.A1(new_n1001), .A2(new_n802), .A3(new_n1034), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(new_n1134), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1222), .A2(new_n1196), .A3(new_n995), .A4(new_n1224), .ZN(G407));
  NAND2_X1  g1025(.A1(new_n678), .A2(G213), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT126), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1196), .A2(new_n1224), .A3(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(G407), .A2(G213), .A3(new_n1228), .ZN(G409));
  AOI21_X1  g1029(.A(new_n802), .B1(new_n1001), .B2(new_n1034), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G390), .A2(new_n1221), .A3(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1042), .A2(new_n1065), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1221), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1041), .B(new_n1233), .C1(new_n1234), .C2(new_n1230), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(G387), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n995), .A2(new_n1232), .A3(new_n1235), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT62), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1196), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1193), .A2(new_n947), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1224), .B1(new_n1242), .B2(new_n1187), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1245), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1198), .A2(new_n1189), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1188), .B1(new_n1247), .B2(KEYINPUT60), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  OR2_X1    g1049(.A1(G384), .A2(KEYINPUT127), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1249), .A2(new_n1219), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G384), .A2(KEYINPUT127), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1249), .A2(new_n1219), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  AND4_X1   g1054(.A1(new_n1240), .A2(new_n1244), .A3(new_n1226), .A4(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1254), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1256), .B2(KEYINPUT62), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1227), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n678), .A2(G213), .A3(G2897), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1254), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1227), .A2(G2897), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1261), .A2(new_n1240), .A3(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1257), .B1(new_n1258), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1239), .B1(new_n1255), .B2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1244), .A2(new_n1226), .A3(new_n1254), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1237), .A2(new_n1270), .A3(new_n1238), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1256), .A2(new_n1268), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1271), .B1(new_n1258), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1244), .A2(new_n1226), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1269), .A2(new_n1273), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1266), .A2(new_n1277), .ZN(G405));
  INV_X1    g1078(.A(new_n1241), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1196), .A2(new_n1134), .A3(new_n1223), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1254), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1280), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1241), .A3(new_n1256), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1239), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1281), .A2(new_n1283), .A3(new_n1238), .A4(new_n1237), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(G402));
endmodule


