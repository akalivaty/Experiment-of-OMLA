//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n193), .B(KEYINPUT69), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT5), .ZN(new_n197));
  OR2_X1    g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G113), .B1(new_n190), .B2(KEYINPUT5), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n195), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT77), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT77), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G104), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(G107), .B1(new_n203), .B2(new_n205), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT78), .B1(new_n211), .B2(new_n207), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT78), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT77), .B(G104), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n213), .B(KEYINPUT3), .C1(new_n214), .C2(G107), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n210), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n208), .A2(G104), .ZN(new_n220));
  OAI21_X1  g034(.A(G101), .B1(new_n211), .B2(new_n220), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n219), .B1(new_n218), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n201), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n210), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n204), .A2(G104), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n202), .A2(KEYINPUT77), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n208), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n213), .B1(new_n228), .B2(KEYINPUT3), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n211), .A2(KEYINPUT78), .A3(new_n207), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n225), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT79), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n216), .A2(KEYINPUT79), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(G101), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT80), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(new_n216), .B2(new_n217), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n236), .B1(new_n235), .B2(new_n238), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n195), .B1(new_n196), .B2(new_n194), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT81), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n212), .A2(new_n215), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT79), .B1(new_n245), .B2(new_n225), .ZN(new_n246));
  AOI211_X1 g060(.A(new_n232), .B(new_n210), .C1(new_n212), .C2(new_n215), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n244), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND4_X1   g064(.A1(new_n244), .A2(new_n233), .A3(new_n234), .A4(new_n249), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n243), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n224), .B1(new_n241), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT86), .ZN(new_n254));
  XNOR2_X1  g068(.A(G110), .B(G122), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(KEYINPUT6), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n224), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n246), .A2(new_n247), .A3(new_n217), .ZN(new_n259));
  INV_X1    g073(.A(new_n238), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT80), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n233), .A2(new_n234), .A3(new_n249), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT81), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n248), .A2(new_n244), .A3(new_n249), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n242), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n258), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n256), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT86), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n257), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n268), .B2(new_n255), .ZN(new_n273));
  INV_X1    g087(.A(new_n255), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n253), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n277));
  INV_X1    g091(.A(G128), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G146), .ZN(new_n281));
  INV_X1    g095(.A(G146), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT65), .B1(new_n282), .B2(G143), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(new_n280), .A3(G146), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n281), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT68), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n279), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  XOR2_X1   g104(.A(G143), .B(G146), .Z(new_n291));
  INV_X1    g105(.A(new_n281), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n277), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G128), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n288), .A2(new_n290), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G125), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(KEYINPUT0), .A2(G128), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(KEYINPUT0), .A2(G128), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n286), .A2(new_n299), .B1(new_n291), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G125), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G224), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G953), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n305), .B(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n271), .A2(new_n276), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT87), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n271), .A2(new_n276), .A3(new_n311), .A4(new_n308), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT89), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT7), .B1(new_n306), .B2(G953), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n305), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n315), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n297), .A2(KEYINPUT89), .A3(new_n304), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n255), .B(KEYINPUT8), .Z(new_n320));
  AND2_X1   g134(.A1(new_n218), .A2(new_n221), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT88), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n193), .B2(new_n197), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(new_n200), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n193), .A2(new_n322), .A3(new_n197), .ZN(new_n325));
  OAI22_X1  g139(.A1(new_n324), .A2(new_n325), .B1(new_n194), .B2(new_n193), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n320), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n218), .A2(new_n221), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n201), .A2(new_n328), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n327), .A2(new_n329), .B1(new_n305), .B2(new_n315), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n319), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n268), .B2(new_n255), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT90), .B1(new_n332), .B2(G902), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT90), .ZN(new_n334));
  INV_X1    g148(.A(G902), .ZN(new_n335));
  AOI211_X1 g149(.A(new_n274), .B(new_n258), .C1(new_n263), .C2(new_n267), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n334), .B(new_n335), .C1(new_n336), .C2(new_n331), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n188), .B1(new_n313), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n188), .ZN(new_n341));
  AOI211_X1 g155(.A(new_n341), .B(new_n338), .C1(new_n310), .C2(new_n312), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n187), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT91), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(KEYINPUT91), .B(new_n187), .C1(new_n340), .C2(new_n342), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G140), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT76), .ZN(new_n348));
  AND2_X1   g162(.A1(KEYINPUT71), .A2(G953), .ZN(new_n349));
  NOR2_X1   g163(.A1(KEYINPUT71), .A2(G953), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n351), .A2(G227), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n348), .B(new_n352), .Z(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n303), .B1(new_n265), .B2(new_n266), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n294), .A2(new_n291), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n279), .A2(new_n289), .A3(new_n286), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n289), .B1(new_n279), .B2(new_n286), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n222), .B2(new_n223), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT10), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n278), .B1(new_n292), .B2(KEYINPUT1), .ZN(new_n363));
  OAI22_X1  g177(.A1(new_n357), .A2(new_n358), .B1(new_n286), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n321), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n263), .A2(new_n355), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT11), .ZN(new_n367));
  INV_X1    g181(.A(G134), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(G137), .ZN(new_n369));
  INV_X1    g183(.A(G137), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(KEYINPUT11), .A3(G134), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(G137), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G131), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(KEYINPUT66), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n373), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n366), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n321), .A2(new_n364), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n328), .A2(new_n295), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(KEYINPUT83), .A3(new_n380), .ZN(new_n381));
  OR2_X1    g195(.A1(new_n380), .A2(KEYINPUT83), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(new_n376), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT12), .B1(new_n376), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n385), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n381), .A2(new_n382), .A3(new_n376), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n354), .B1(new_n378), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n391), .B1(new_n366), .B2(new_n377), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n263), .A2(new_n355), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n361), .A2(new_n365), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT85), .A3(new_n376), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n395), .A2(new_n376), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(new_n353), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n390), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G469), .B1(new_n400), .B2(G902), .ZN(new_n401));
  INV_X1    g215(.A(G469), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n354), .B1(new_n397), .B2(new_n378), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n378), .A2(new_n354), .A3(new_n389), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n402), .B(new_n335), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT9), .B(G234), .ZN(new_n407));
  OAI21_X1  g221(.A(G221), .B1(new_n407), .B2(G902), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n191), .A2(G122), .ZN(new_n410));
  INV_X1    g224(.A(G122), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(G116), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(new_n208), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n278), .A2(G143), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n280), .A2(G128), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n368), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n415), .A2(KEYINPUT13), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n415), .A2(KEYINPUT13), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n419), .A2(new_n420), .A3(new_n416), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n414), .B(new_n418), .C1(new_n368), .C2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n417), .B(new_n368), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n413), .A2(new_n208), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT14), .B1(new_n411), .B2(G116), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(KEYINPUT94), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT14), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n410), .B1(new_n428), .B2(new_n412), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n208), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n422), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G217), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n407), .A2(new_n432), .A3(G953), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n431), .B(new_n433), .Z(new_n434));
  AND2_X1   g248(.A1(new_n434), .A2(new_n335), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT95), .ZN(new_n436));
  INV_X1    g250(.A(G478), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(KEYINPUT15), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n436), .B(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G113), .B(G122), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(new_n202), .ZN(new_n442));
  INV_X1    g256(.A(G140), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G125), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n296), .A2(G140), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(G146), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT73), .ZN(new_n448));
  INV_X1    g262(.A(new_n446), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n282), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G237), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n351), .A2(G214), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n280), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n351), .A2(G143), .A3(G214), .A4(new_n451), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(KEYINPUT18), .A3(G131), .ZN(new_n456));
  NAND2_X1  g270(.A1(KEYINPUT18), .A2(G131), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n453), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(G131), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n453), .A2(new_n374), .A3(new_n454), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(KEYINPUT17), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT16), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n443), .A3(G125), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT72), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n465), .B1(new_n446), .B2(new_n464), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(new_n468), .B2(KEYINPUT72), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n469), .A2(G146), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(G146), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n460), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n442), .B(new_n459), .C1(new_n463), .C2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n446), .B(KEYINPUT19), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n475), .A2(G146), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n471), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT92), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(KEYINPUT92), .A3(new_n471), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n462), .A3(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n481), .A2(new_n459), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n474), .B1(new_n482), .B2(new_n442), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT93), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT20), .ZN(new_n485));
  NOR2_X1   g299(.A1(G475), .A2(G902), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n483), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n474), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n442), .B1(new_n481), .B2(new_n459), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n485), .B(new_n486), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT93), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT20), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n487), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n459), .B1(new_n463), .B2(new_n473), .ZN(new_n495));
  INV_X1    g309(.A(new_n442), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(G902), .B1(new_n497), .B2(new_n474), .ZN(new_n498));
  INV_X1    g312(.A(G475), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(G234), .A2(G237), .ZN(new_n502));
  INV_X1    g316(.A(G953), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(G952), .A3(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT96), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n351), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n507), .A2(G902), .A3(new_n502), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT21), .B(G898), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n440), .A2(new_n501), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n409), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n345), .A2(new_n346), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT97), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G472), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT31), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n351), .A2(G210), .A3(new_n451), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n519), .B(KEYINPUT27), .Z(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT26), .B(G101), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n520), .B(new_n521), .Z(new_n522));
  NAND2_X1  g336(.A1(new_n373), .A2(new_n374), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n370), .A2(G134), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n372), .A3(G131), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI22_X1  g341(.A1(new_n295), .A2(new_n527), .B1(new_n377), .B2(new_n303), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT64), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT30), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n359), .A2(new_n526), .B1(new_n376), .B2(new_n302), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(KEYINPUT64), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n242), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n242), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT70), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI211_X1 g351(.A(KEYINPUT70), .B(new_n242), .C1(new_n530), .C2(new_n533), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n518), .B(new_n522), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n522), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT28), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n528), .A2(new_n243), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n535), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT28), .B1(new_n532), .B2(new_n242), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT70), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n534), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n534), .B2(new_n536), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n518), .B1(new_n549), .B2(new_n522), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n517), .B(new_n335), .C1(new_n546), .C2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT32), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n537), .A2(new_n538), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT31), .B1(new_n554), .B2(new_n540), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n545), .A3(new_n539), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n556), .A2(KEYINPUT32), .A3(new_n517), .A4(new_n335), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n540), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n543), .A2(new_n540), .A3(new_n544), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(KEYINPUT29), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(G902), .B1(new_n559), .B2(KEYINPUT29), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(G472), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n553), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n470), .A2(new_n471), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT23), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n189), .B2(G128), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n278), .A2(KEYINPUT23), .A3(G119), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n568), .B(new_n569), .C1(G119), .C2(new_n278), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G110), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT24), .B(G110), .Z(new_n572));
  XNOR2_X1  g386(.A(G119), .B(G128), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n566), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n351), .A2(G221), .A3(G234), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT22), .B(G137), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  OAI22_X1  g394(.A1(new_n570), .A2(G110), .B1(new_n573), .B2(new_n572), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n471), .A2(new_n448), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n580), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n575), .B1(new_n470), .B2(new_n471), .ZN(new_n585));
  INV_X1    g399(.A(new_n582), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n583), .A2(new_n587), .A3(new_n335), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT25), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n583), .A2(new_n587), .A3(KEYINPUT25), .A4(new_n335), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n432), .B1(G234), .B2(new_n335), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT74), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n592), .A2(KEYINPUT74), .A3(new_n593), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n583), .A2(new_n587), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n599), .B(KEYINPUT75), .Z(new_n600));
  NOR3_X1   g414(.A1(new_n600), .A2(G902), .A3(new_n593), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n565), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n345), .A2(KEYINPUT97), .A3(new_n346), .A4(new_n513), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n516), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT98), .B(G101), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G3));
  NOR2_X1   g422(.A1(new_n343), .A2(new_n510), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n556), .A2(new_n335), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(new_n551), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n602), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n409), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n494), .A2(new_n500), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n434), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(G478), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n437), .A2(new_n335), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n435), .B2(new_n437), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n609), .A2(new_n614), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT99), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT34), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n628));
  OAI22_X1  g442(.A1(new_n490), .A2(new_n628), .B1(new_n498), .B2(new_n499), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n490), .A2(new_n628), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n629), .B1(new_n630), .B2(new_n493), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n631), .A2(new_n439), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n609), .A2(new_n614), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NAND2_X1  g449(.A1(new_n577), .A2(new_n582), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n584), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n638), .B(new_n335), .C1(new_n432), .C2(G234), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n596), .A2(new_n597), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n612), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT101), .Z(new_n642));
  NAND3_X1  g456(.A1(new_n516), .A2(new_n605), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  INV_X1    g459(.A(new_n187), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n257), .A2(new_n270), .B1(new_n273), .B2(new_n275), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n311), .B1(new_n647), .B2(new_n308), .ZN(new_n648));
  INV_X1    g462(.A(new_n312), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n339), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n341), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n313), .A2(new_n188), .A3(new_n339), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n646), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n653), .A2(new_n565), .ZN(new_n654));
  INV_X1    g468(.A(new_n408), .ZN(new_n655));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n506), .B1(new_n656), .B2(new_n508), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n631), .A2(new_n640), .A3(new_n439), .A4(new_n658), .ZN(new_n659));
  AOI211_X1 g473(.A(new_n655), .B(new_n659), .C1(new_n401), .C2(new_n405), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G128), .ZN(G30));
  NAND2_X1  g476(.A1(new_n651), .A2(new_n652), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT38), .ZN(new_n664));
  NOR4_X1   g478(.A1(new_n440), .A2(new_n501), .A3(new_n646), .A4(new_n640), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n655), .B1(new_n401), .B2(new_n405), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n657), .B(new_n668), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT40), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n554), .A2(new_n522), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n542), .A2(new_n535), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n335), .B1(new_n676), .B2(new_n522), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n553), .A2(new_n557), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT102), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n553), .A2(new_n557), .A3(new_n681), .A4(new_n678), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n666), .A2(new_n672), .A3(new_n673), .A4(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n664), .A2(new_n683), .A3(new_n665), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT104), .B1(new_n685), .B2(new_n671), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n280), .ZN(G45));
  NAND4_X1  g502(.A1(new_n615), .A2(new_n640), .A3(new_n621), .A4(new_n658), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n655), .B(new_n689), .C1(new_n401), .C2(new_n405), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n654), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  INV_X1    g506(.A(new_n404), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n398), .B1(new_n392), .B2(new_n396), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n693), .B1(new_n694), .B2(new_n354), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n335), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n408), .A3(new_n405), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n603), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n609), .A2(new_n623), .A3(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT41), .B(G113), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT105), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n700), .B(new_n702), .ZN(G15));
  NAND3_X1  g517(.A1(new_n609), .A2(new_n632), .A3(new_n699), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  OAI21_X1  g519(.A(KEYINPUT106), .B1(new_n343), .B2(new_n698), .ZN(new_n706));
  INV_X1    g520(.A(new_n405), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n402), .B1(new_n695), .B2(new_n335), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n707), .A2(new_n708), .A3(new_n655), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n653), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n565), .A2(new_n640), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n512), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  INV_X1    g530(.A(new_n613), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n440), .A2(new_n501), .A3(new_n510), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(new_n653), .A3(new_n709), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  NOR2_X1   g534(.A1(new_n622), .A2(new_n657), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n612), .A2(new_n640), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n706), .B2(new_n711), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n296), .ZN(G27));
  AND2_X1   g538(.A1(new_n539), .A2(new_n545), .ZN(new_n725));
  AOI21_X1  g539(.A(G902), .B1(new_n725), .B2(new_n555), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n727), .A3(KEYINPUT32), .A4(new_n517), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT108), .B1(new_n551), .B2(new_n552), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT107), .B1(new_n551), .B2(new_n552), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n731), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n729), .A3(new_n728), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n734), .A3(new_n564), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n602), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n340), .A2(new_n342), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n187), .A3(new_n667), .A4(new_n721), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT42), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n663), .A2(new_n409), .A3(new_n646), .ZN(new_n740));
  INV_X1    g554(.A(new_n721), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(KEYINPUT42), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n604), .A3(new_n742), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NAND2_X1  g559(.A1(new_n632), .A2(new_n658), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n746), .B(KEYINPUT109), .Z(new_n747));
  NAND3_X1  g561(.A1(new_n740), .A2(new_n604), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT110), .B(G134), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G36));
  OR2_X1    g564(.A1(new_n400), .A2(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n400), .A2(KEYINPUT45), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(G469), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(G469), .A2(G902), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n707), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n756), .B2(new_n755), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n408), .A3(new_n669), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT111), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(new_n761), .A3(new_n408), .A4(new_n669), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n663), .A2(new_n646), .ZN(new_n763));
  INV_X1    g577(.A(new_n612), .ZN(new_n764));
  INV_X1    g578(.A(new_n621), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n766));
  OAI22_X1  g580(.A1(new_n765), .A2(new_n615), .B1(KEYINPUT112), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n501), .A2(new_n621), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n764), .A2(new_n640), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n763), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n772), .B2(new_n771), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n760), .A2(new_n762), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  NOR3_X1   g590(.A1(new_n741), .A2(new_n565), .A3(new_n602), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n763), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT113), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n758), .A2(KEYINPUT47), .A3(new_n408), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT47), .B1(new_n758), .B2(new_n408), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT114), .B(G140), .Z(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G42));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n786));
  INV_X1    g600(.A(new_n722), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n712), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n653), .B(new_n565), .C1(new_n660), .C2(new_n690), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n640), .A2(new_n657), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n655), .B(new_n790), .C1(new_n405), .C2(new_n401), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n440), .A2(new_n501), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n653), .A2(new_n683), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n786), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n789), .A2(new_n793), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n723), .A2(new_n796), .A3(KEYINPUT116), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n785), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n622), .B1(new_n440), .B2(new_n615), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n511), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n345), .A2(new_n614), .A3(new_n346), .A4(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n606), .A2(new_n643), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n440), .A2(new_n631), .A3(new_n658), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n722), .B1(new_n713), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n740), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n739), .A2(new_n743), .A3(new_n748), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n715), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n700), .A2(new_n704), .A3(new_n719), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n788), .A2(new_n794), .A3(new_n786), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT116), .B1(new_n723), .B2(new_n796), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT52), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n798), .A2(new_n802), .A3(new_n809), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n700), .A2(new_n704), .A3(new_n719), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n748), .A2(new_n805), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n744), .A2(new_n817), .A3(new_n715), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n606), .A2(new_n643), .A3(new_n801), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n785), .B1(new_n788), .B2(new_n794), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n821), .A2(KEYINPUT53), .A3(new_n798), .A4(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n815), .A2(new_n816), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT117), .B1(new_n813), .B2(new_n814), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT52), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(new_n810), .B2(new_n811), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT53), .A4(new_n821), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n798), .A2(new_n823), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n802), .A2(new_n809), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n814), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n826), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n825), .B1(KEYINPUT54), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n663), .A2(new_n698), .A3(new_n646), .ZN(new_n838));
  INV_X1    g652(.A(new_n683), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n602), .A3(new_n506), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n501), .A3(new_n765), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n770), .A2(new_n506), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n641), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n664), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n717), .A2(new_n843), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n646), .A2(new_n847), .A3(new_n709), .A4(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(KEYINPUT50), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(KEYINPUT50), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n842), .B(new_n846), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n848), .A2(new_n763), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n780), .A2(new_n781), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n707), .A2(new_n708), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n655), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n853), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n837), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n844), .ZN(new_n859));
  INV_X1    g673(.A(new_n736), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(KEYINPUT119), .A3(KEYINPUT48), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n841), .A2(new_n623), .ZN(new_n862));
  XOR2_X1   g676(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n844), .B2(new_n736), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n712), .A2(new_n848), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n858), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n852), .A2(new_n857), .A3(new_n837), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n836), .A2(new_n869), .A3(KEYINPUT118), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(G952), .A3(new_n503), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n836), .A2(new_n869), .ZN(new_n872));
  OAI21_X1  g686(.A(G953), .B1(new_n872), .B2(KEYINPUT118), .ZN(new_n873));
  INV_X1    g687(.A(new_n768), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n602), .A3(new_n187), .A4(new_n408), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT115), .Z(new_n876));
  INV_X1    g690(.A(KEYINPUT49), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n855), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n855), .A2(new_n877), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n839), .A3(new_n847), .A4(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n871), .A2(new_n873), .A3(new_n881), .ZN(G75));
  NOR2_X1   g696(.A1(new_n351), .A2(G952), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n335), .B1(new_n815), .B2(new_n824), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n885), .B2(G210), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n647), .B(new_n308), .Z(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n884), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n886), .B2(new_n888), .ZN(G51));
  INV_X1    g704(.A(new_n825), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n815), .A2(new_n824), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n754), .B(KEYINPUT57), .Z(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n695), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n885), .A2(G469), .A3(new_n752), .A4(new_n751), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n883), .B1(new_n897), .B2(new_n898), .ZN(G54));
  NAND3_X1  g713(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n900));
  INV_X1    g714(.A(new_n483), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n903), .A3(new_n883), .ZN(G60));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n619), .B(KEYINPUT59), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n835), .A2(KEYINPUT54), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(new_n891), .ZN(new_n908));
  INV_X1    g722(.A(new_n617), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g724(.A(KEYINPUT120), .B(new_n617), .C1(new_n836), .C2(new_n906), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n617), .A2(new_n906), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n883), .B1(new_n894), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(G63));
  XNOR2_X1  g728(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n432), .A2(new_n335), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n892), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT122), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n892), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n600), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n892), .B2(new_n917), .ZN(new_n923));
  INV_X1    g737(.A(new_n917), .ZN(new_n924));
  AOI211_X1 g738(.A(KEYINPUT122), .B(new_n924), .C1(new_n815), .C2(new_n824), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n638), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n926), .A3(new_n884), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n922), .A2(new_n926), .A3(KEYINPUT61), .A4(new_n884), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(G66));
  OAI21_X1  g745(.A(G953), .B1(new_n509), .B2(new_n306), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n802), .A2(new_n715), .A3(new_n817), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n934), .B2(new_n507), .ZN(new_n935));
  INV_X1    g749(.A(new_n647), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(G898), .B2(new_n351), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT123), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n935), .B(new_n938), .ZN(G69));
  NAND2_X1  g753(.A1(new_n530), .A2(new_n533), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n475), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(G900), .B2(new_n507), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n788), .A2(new_n789), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n782), .A2(new_n748), .A3(new_n943), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n343), .A2(new_n501), .A3(new_n440), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n760), .A2(new_n860), .A3(new_n762), .A4(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n944), .A2(new_n744), .A3(new_n775), .A4(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n942), .B1(new_n947), .B2(new_n507), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n684), .A2(new_n943), .A3(new_n686), .A4(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n740), .A2(new_n604), .A3(new_n669), .A4(new_n799), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n775), .A2(new_n782), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n684), .A2(new_n943), .A3(new_n686), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(KEYINPUT62), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n507), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n941), .B(KEYINPUT124), .Z(new_n958));
  OAI21_X1  g772(.A(new_n948), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT126), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n961), .B(new_n948), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n351), .B1(G227), .B2(G900), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n960), .A2(new_n964), .A3(new_n962), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(G72));
  AND3_X1   g782(.A1(new_n952), .A2(new_n675), .A3(new_n956), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n947), .A2(new_n522), .A3(new_n554), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n934), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  NOR2_X1   g787(.A1(new_n554), .A2(new_n540), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n974), .A2(KEYINPUT127), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(new_n558), .Z(new_n976));
  NAND3_X1  g790(.A1(new_n835), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n974), .A2(new_n973), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n883), .B1(new_n978), .B2(new_n558), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n971), .A2(new_n977), .A3(new_n979), .ZN(G57));
endmodule


