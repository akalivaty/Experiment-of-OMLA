//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n612, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(G125), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n463), .B(G125), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G101), .A3(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  OAI211_X1 g049(.A(G137), .B(new_n472), .C1(new_n466), .C2(new_n467), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT69), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n464), .A2(new_n477), .A3(G137), .A4(new_n472), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n474), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT70), .ZN(new_n485));
  OR2_X1    g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n472), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n489));
  AOI22_X1  g064(.A1(G124), .A2(new_n488), .B1(new_n489), .B2(G136), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n485), .A2(new_n490), .ZN(G162));
  OR2_X1    g066(.A1(new_n472), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n472), .C1(new_n466), .C2(new_n467), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n464), .A2(new_n500), .A3(G138), .A4(new_n472), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(G164));
  OR2_X1    g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  INV_X1    g088(.A(new_n504), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n512), .A2(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n508), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  XOR2_X1   g097(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n526), .B1(new_n509), .B2(new_n510), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n518), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n525), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n530), .B1(new_n528), .B2(new_n529), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n507), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT73), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT74), .B(G90), .Z(new_n540));
  AOI22_X1  g115(.A1(new_n532), .A2(new_n540), .B1(G52), .B2(new_n527), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n507), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n512), .A2(new_n546), .B1(new_n518), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  OAI211_X1 g130(.A(G53), .B(G543), .C1(new_n516), .C2(new_n517), .ZN(new_n556));
  XNOR2_X1  g131(.A(KEYINPUT76), .B(KEYINPUT9), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT77), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(KEYINPUT76), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n527), .A2(new_n559), .A3(G53), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n558), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n556), .A2(KEYINPUT75), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n511), .A2(new_n568), .A3(G53), .A4(G543), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n569), .A3(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n566), .A2(new_n570), .A3(KEYINPUT78), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n514), .A2(new_n515), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(new_n532), .B2(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n575), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G168), .ZN(G286));
  NAND2_X1  g157(.A1(new_n532), .A2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n527), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  OAI211_X1 g161(.A(G48), .B(G543), .C1(new_n516), .C2(new_n517), .ZN(new_n587));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n518), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(G61), .B1(new_n514), .B2(new_n515), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n507), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n532), .A2(G85), .B1(G47), .B2(new_n527), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n507), .B2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(new_n532), .A2(G92), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n577), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G54), .B2(new_n527), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G284));
  OAI21_X1  g183(.A(new_n607), .B1(G171), .B2(new_n606), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT79), .ZN(new_n611));
  INV_X1    g186(.A(new_n580), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n573), .B2(new_n574), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n611), .B1(G868), .B2(new_n613), .ZN(G297));
  OAI21_X1  g189(.A(new_n611), .B1(G868), .B2(new_n613), .ZN(G280));
  INV_X1    g190(.A(new_n605), .ZN(new_n616));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G860), .ZN(G148));
  OR2_X1    g193(.A1(new_n545), .A2(new_n548), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n606), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n605), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n489), .A2(G2104), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n624), .B(KEYINPUT81), .ZN(new_n629));
  INV_X1    g204(.A(new_n627), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n489), .A2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n488), .A2(G123), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n472), .A2(G111), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n637), .B(new_n638), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT82), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n635), .A2(new_n636), .A3(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  OAI21_X1  g231(.A(G14), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n655), .B2(new_n656), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n655), .A2(new_n658), .A3(new_n656), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(G401));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT84), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT18), .Z(new_n668));
  OR2_X1    g243(.A1(new_n664), .A2(new_n666), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n666), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n665), .B(KEYINPUT17), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n665), .B(KEYINPUT85), .Z(new_n673));
  OAI211_X1 g248(.A(new_n668), .B(new_n672), .C1(new_n669), .C2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n678), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1981), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT86), .B(KEYINPUT87), .Z(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  INV_X1    g268(.A(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n692), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  NAND3_X1  g272(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT26), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT98), .ZN(new_n701));
  AOI211_X1 g276(.A(new_n699), .B(new_n701), .C1(G141), .C2(new_n489), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n488), .A2(G129), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT97), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n707), .B2(G32), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT27), .B(G1996), .ZN(new_n710));
  INV_X1    g285(.A(G2078), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(G27), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT101), .Z(new_n713));
  AOI22_X1  g288(.A1(new_n488), .A2(G126), .B1(new_n492), .B2(new_n494), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n500), .B1(new_n489), .B2(G138), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n713), .B1(new_n717), .B2(G29), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n709), .A2(new_n710), .B1(new_n711), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n709), .B2(new_n710), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n707), .A2(G35), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G162), .B2(new_n707), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT29), .B(G2090), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G5), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G171), .B2(new_n725), .ZN(new_n727));
  OAI221_X1 g302(.A(new_n724), .B1(new_n711), .B2(new_n718), .C1(new_n727), .C2(G1961), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n707), .B1(KEYINPUT24), .B2(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(KEYINPUT24), .B2(G34), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n480), .B2(G29), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT30), .B(G28), .ZN(new_n734));
  OR2_X1    g309(.A1(KEYINPUT31), .A2(G11), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n734), .A2(new_n707), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n642), .B2(new_n707), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT100), .Z(new_n739));
  OR4_X1    g314(.A1(new_n720), .A2(new_n728), .A3(new_n733), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n489), .A2(G140), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n488), .A2(G128), .ZN(new_n742));
  OR2_X1    g317(.A1(G104), .A2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n743), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT94), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n707), .A2(G26), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT28), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G2067), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n725), .A2(G19), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n549), .B2(new_n725), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1341), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n616), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G4), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1348), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n752), .B(new_n759), .C1(new_n758), .C2(new_n757), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT95), .ZN(new_n761));
  INV_X1    g336(.A(G21), .ZN(new_n762));
  AOI21_X1  g337(.A(KEYINPUT99), .B1(new_n725), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G286), .A2(new_n725), .ZN(new_n764));
  MUX2_X1   g339(.A(new_n763), .B(KEYINPUT99), .S(new_n764), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1966), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n464), .A2(G127), .ZN(new_n767));
  AND2_X1   g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(G2105), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT96), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(KEYINPUT96), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT25), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n489), .A2(G139), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n770), .A2(new_n771), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  MUX2_X1   g350(.A(G33), .B(new_n775), .S(G29), .Z(new_n776));
  AND2_X1   g351(.A1(new_n776), .A2(G2072), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G1961), .B2(new_n727), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G2072), .B2(new_n776), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n740), .A2(new_n761), .A3(new_n766), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n725), .A2(G22), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G166), .B2(new_n725), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G1971), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n725), .A2(G23), .ZN(new_n784));
  INV_X1    g359(.A(G288), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n725), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT33), .B(G1976), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT93), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n786), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G6), .A2(G16), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n593), .B2(G16), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT32), .B(G1981), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n783), .A2(new_n789), .A3(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n707), .A2(G25), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n488), .A2(G119), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT88), .Z(new_n798));
  NOR2_X1   g373(.A1(G95), .A2(G2105), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT89), .Z(new_n800));
  INV_X1    g375(.A(G2104), .ZN(new_n801));
  INV_X1    g376(.A(G107), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G2105), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n800), .A2(new_n803), .B1(G131), .B2(new_n489), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT90), .Z(new_n806));
  AOI21_X1  g381(.A(new_n796), .B1(new_n806), .B2(G29), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G1991), .Z(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n807), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n725), .A2(G24), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT91), .Z(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G290), .B2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT92), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(new_n694), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n794), .A2(KEYINPUT34), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n795), .A2(new_n810), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT36), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n725), .A2(G20), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT23), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n613), .B2(new_n725), .ZN(new_n821));
  INV_X1    g396(.A(G1956), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n780), .A2(new_n818), .A3(new_n823), .ZN(G150));
  INV_X1    g399(.A(G150), .ZN(G311));
  NAND2_X1  g400(.A1(new_n616), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  INV_X1    g403(.A(G67), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n577), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT102), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n832), .B(new_n828), .C1(new_n577), .C2(new_n829), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(G651), .A3(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT103), .B(G93), .Z(new_n835));
  AOI22_X1  g410(.A1(new_n532), .A2(new_n835), .B1(G55), .B2(new_n527), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n549), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n549), .B1(new_n834), .B2(new_n836), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n827), .B(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT104), .B(G860), .Z(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n844), .B1(new_n834), .B2(new_n836), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(G145));
  XOR2_X1   g423(.A(new_n480), .B(G162), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT105), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n642), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n849), .A2(KEYINPUT105), .ZN(new_n852));
  INV_X1    g427(.A(new_n642), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(KEYINPUT105), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  INV_X1    g432(.A(G118), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(G2105), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(G130), .B2(new_n488), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n489), .A2(G142), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n628), .B2(new_n631), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n805), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n628), .A2(new_n631), .A3(new_n862), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n628), .A2(new_n631), .A3(new_n862), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n805), .B1(new_n868), .B2(new_n863), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n745), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n775), .B(new_n705), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n499), .A2(new_n501), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n874), .A2(new_n875), .A3(new_n714), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n874), .B2(new_n714), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n867), .A2(new_n869), .A3(new_n745), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n873), .A2(new_n878), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n872), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n872), .A2(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n856), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n872), .A2(new_n880), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n879), .A2(new_n881), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n889), .A2(new_n855), .A3(new_n851), .A4(new_n882), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n885), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(G395));
  XOR2_X1   g468(.A(new_n840), .B(new_n621), .Z(new_n894));
  NAND2_X1  g469(.A1(G299), .A2(new_n616), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n613), .A2(new_n605), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(KEYINPUT108), .A3(new_n896), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n613), .A2(new_n605), .A3(KEYINPUT108), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OR3_X1    g474(.A1(new_n894), .A2(new_n899), .A3(KEYINPUT109), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n897), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n902), .A3(new_n896), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n894), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT109), .B1(new_n894), .B2(new_n899), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(G303), .B(new_n785), .ZN(new_n907));
  XNOR2_X1  g482(.A(G290), .B(new_n593), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT42), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n900), .A2(new_n910), .A3(new_n904), .A4(new_n905), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n606), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n834), .A2(new_n836), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n606), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n914), .A2(new_n917), .ZN(G295));
  OR3_X1    g493(.A1(new_n914), .A2(KEYINPUT110), .A3(new_n917), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT110), .B1(new_n914), .B2(new_n917), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(G331));
  INV_X1    g496(.A(new_n909), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n902), .B1(new_n895), .B2(new_n896), .ZN(new_n923));
  OAI21_X1  g498(.A(G168), .B1(new_n838), .B2(new_n839), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n915), .A2(new_n619), .ZN(new_n925));
  NAND3_X1  g500(.A1(G286), .A2(new_n925), .A3(new_n837), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(G301), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n926), .A3(G171), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n923), .B(new_n930), .C1(new_n902), .C2(new_n899), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n924), .A2(new_n926), .A3(G171), .ZN(new_n932));
  AOI21_X1  g507(.A(G171), .B1(new_n924), .B2(new_n926), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n898), .B(new_n897), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT112), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n930), .A2(new_n936), .A3(new_n898), .A4(new_n897), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n922), .B1(new_n931), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n932), .A2(new_n933), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n901), .A3(new_n903), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(new_n909), .A3(new_n934), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n942), .A2(new_n886), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n942), .A2(new_n886), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n909), .B1(new_n941), .B2(new_n934), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(KEYINPUT111), .A3(new_n948), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n948), .A2(KEYINPUT111), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n939), .A2(new_n943), .A3(KEYINPUT43), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(new_n956), .ZN(G397));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT45), .B1(new_n717), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT68), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n961), .A2(new_n468), .B1(G113), .B2(G2104), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n479), .B(G40), .C1(new_n962), .C2(new_n472), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G1384), .B1(new_n874), .B2(new_n714), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT45), .ZN(new_n966));
  AOI21_X1  g541(.A(G1966), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n476), .A2(new_n478), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(G40), .A3(new_n473), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n961), .A2(new_n468), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n472), .B1(new_n970), .B2(new_n462), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n965), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n975));
  AND4_X1   g550(.A1(new_n732), .A2(new_n972), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(KEYINPUT122), .B(G8), .C1(new_n967), .C2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  NOR2_X1   g553(.A1(G168), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(KEYINPUT51), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(G164), .B2(G1384), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n972), .A2(new_n966), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1966), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n972), .A2(new_n974), .A3(new_n975), .A4(new_n732), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n978), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(KEYINPUT122), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT123), .B1(new_n981), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT122), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n992), .A2(new_n732), .B1(new_n984), .B2(new_n985), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n991), .B1(new_n993), .B2(new_n978), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT123), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n994), .A2(new_n995), .A3(new_n977), .A4(new_n980), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT51), .B1(new_n988), .B2(new_n979), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n990), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n979), .B1(new_n967), .B2(new_n976), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT62), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n1002), .A3(new_n999), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n717), .A2(KEYINPUT106), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n874), .A2(new_n875), .A3(new_n714), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(KEYINPUT45), .A3(new_n958), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n964), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1004), .B1(new_n1008), .B2(G2078), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1009), .A2(KEYINPUT124), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n992), .A2(G1961), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1011), .B1(new_n1009), .B2(KEYINPUT124), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1004), .A2(G2078), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n964), .A2(new_n966), .A3(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1010), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT115), .B(G1971), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n964), .B2(new_n1007), .ZN(new_n1017));
  INV_X1    g592(.A(G2090), .ZN(new_n1018));
  AND4_X1   g593(.A1(new_n1018), .A2(new_n972), .A3(new_n974), .A4(new_n975), .ZN(new_n1019));
  OAI21_X1  g594(.A(G8), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G303), .A2(G8), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1020), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n583), .A2(G1976), .A3(new_n584), .A4(new_n585), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n717), .A2(new_n958), .ZN(new_n1029));
  OAI211_X1 g604(.A(G8), .B(new_n1028), .C1(new_n963), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1030), .A2(new_n1031), .A3(KEYINPUT52), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1030), .B2(KEYINPUT52), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n978), .B1(new_n972), .B2(new_n965), .ZN(new_n1035));
  OAI21_X1  g610(.A(G1981), .B1(new_n589), .B2(new_n592), .ZN(new_n1036));
  INV_X1    g611(.A(G61), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n503), .B2(new_n504), .ZN(new_n1038));
  INV_X1    g613(.A(new_n591), .ZN(new_n1039));
  OAI21_X1  g614(.A(G651), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1981), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n505), .A2(new_n511), .A3(G86), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n587), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1036), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT49), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1036), .A2(new_n1043), .A3(KEYINPUT49), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1035), .B(new_n1046), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1976), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1035), .A2(new_n1028), .A3(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(G8), .B(new_n1025), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1027), .A2(new_n1034), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1015), .A2(G301), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1001), .A2(new_n1003), .A3(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1051), .B(new_n1054), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(new_n1056), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1051), .A2(new_n1052), .A3(new_n785), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1043), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1061), .B1(new_n1035), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n963), .B1(KEYINPUT50), .B2(new_n1029), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(new_n1018), .A3(new_n974), .ZN(new_n1066));
  INV_X1    g641(.A(G40), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1067), .B(new_n474), .C1(new_n476), .C2(new_n478), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n471), .B(new_n1068), .C1(new_n965), .C2(KEYINPUT45), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n876), .A2(new_n877), .A3(G1384), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(KEYINPUT45), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1066), .B1(new_n1071), .B2(new_n1016), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1025), .B1(new_n1072), .B2(G8), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1056), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1073), .A2(new_n1074), .A3(new_n1060), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n988), .A2(G168), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT63), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT63), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1057), .A2(new_n1079), .A3(new_n1076), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1064), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n972), .A2(new_n975), .ZN(new_n1084));
  INV_X1    g659(.A(new_n974), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n822), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n964), .A2(new_n1007), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n566), .A2(KEYINPUT78), .A3(new_n570), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT78), .B1(new_n566), .B2(new_n570), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT57), .B(new_n580), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n571), .A2(new_n580), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n575), .A2(new_n1093), .A3(KEYINPUT57), .A4(new_n580), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1097), .A2(new_n1098), .A3(KEYINPUT120), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT120), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1089), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1348), .B1(new_n1065), .B2(new_n974), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n972), .A2(new_n965), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(G2067), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n616), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n1089), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1107), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1101), .A2(new_n1112), .ZN(new_n1113));
  NOR4_X1   g688(.A1(new_n1102), .A2(new_n1104), .A3(KEYINPUT60), .A4(new_n605), .ZN(new_n1114));
  OAI221_X1 g689(.A(new_n605), .B1(G2067), .B2(new_n1103), .C1(new_n992), .C2(G1348), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1105), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1114), .B1(new_n1116), .B2(KEYINPUT60), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1103), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT58), .B(G1341), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1008), .A2(G1996), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n549), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT59), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1123), .A3(new_n549), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1113), .A2(new_n1117), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n1107), .B2(new_n1089), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1107), .A2(new_n1089), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1107), .A2(new_n1089), .A3(new_n1127), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT61), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1108), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n472), .B1(new_n962), .B2(KEYINPUT125), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n969), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1070), .B2(KEYINPUT45), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1139), .A2(new_n1007), .A3(new_n1013), .A4(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1142));
  XNOR2_X1  g717(.A(G301), .B(KEYINPUT54), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1010), .A2(new_n1012), .A3(new_n1014), .A4(new_n1143), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1057), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1133), .A2(new_n1000), .A3(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT118), .B(new_n1064), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1059), .A2(new_n1083), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(G290), .A2(G1986), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT113), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(G1986), .B2(G290), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1070), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT114), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1155), .B2(G1996), .ZN(new_n1158));
  INV_X1    g733(.A(G1996), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1154), .A2(KEYINPUT114), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n706), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n745), .B(new_n751), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n706), .B2(new_n1159), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1154), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n805), .B(new_n809), .ZN(new_n1167));
  AOI211_X1 g742(.A(new_n1156), .B(new_n1166), .C1(new_n1154), .C2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1150), .A2(new_n1168), .ZN(new_n1169));
  OR3_X1    g744(.A1(new_n1166), .A2(new_n806), .A3(new_n809), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n871), .A2(new_n751), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1155), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT48), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1167), .A2(new_n1154), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1162), .A2(new_n1174), .A3(new_n1165), .A4(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1155), .B1(new_n706), .B2(new_n1163), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT46), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1161), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1158), .A2(KEYINPUT46), .A3(new_n1160), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT47), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1176), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1172), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1169), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n1189));
  NOR2_X1   g763(.A1(G227), .A2(new_n460), .ZN(new_n1190));
  INV_X1    g764(.A(new_n1190), .ZN(new_n1191));
  OAI21_X1  g765(.A(new_n1189), .B1(G401), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g766(.A(new_n661), .ZN(new_n1193));
  NOR2_X1   g767(.A1(new_n1193), .A2(new_n659), .ZN(new_n1194));
  OAI211_X1 g768(.A(KEYINPUT127), .B(new_n1190), .C1(new_n1194), .C2(new_n657), .ZN(new_n1195));
  AND4_X1   g769(.A1(new_n696), .A2(new_n1192), .A3(new_n891), .A4(new_n1195), .ZN(new_n1196));
  AND3_X1   g770(.A1(new_n1196), .A2(new_n949), .A3(new_n950), .ZN(G308));
  NAND3_X1  g771(.A1(new_n1196), .A2(new_n949), .A3(new_n950), .ZN(G225));
endmodule


