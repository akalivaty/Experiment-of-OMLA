//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT74), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT76), .ZN(new_n195));
  OR3_X1    g009(.A1(new_n191), .A2(KEYINPUT76), .A3(G125), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT16), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT16), .B1(new_n191), .B2(G125), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G125), .B(G140), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT64), .B(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT24), .B(G110), .Z(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G119), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G128), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT75), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n207), .A2(G119), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n206), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n217), .B(new_n212), .C1(new_n210), .C2(KEYINPUT23), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(G110), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n205), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT77), .B1(new_n202), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n216), .A2(new_n219), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n222), .A2(new_n223), .A3(new_n201), .A4(new_n205), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n197), .A2(new_n225), .A3(new_n199), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n201), .A2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n211), .A2(new_n215), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n228), .A2(new_n206), .B1(G110), .B2(new_n218), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n221), .A2(new_n224), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT22), .B(G137), .ZN(new_n232));
  INV_X1    g046(.A(G221), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n233), .A2(new_n187), .A3(G953), .ZN(new_n234));
  XOR2_X1   g048(.A(new_n232), .B(new_n234), .Z(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G902), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n221), .A2(new_n224), .A3(new_n230), .A4(new_n235), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n237), .A2(KEYINPUT25), .A3(new_n238), .A4(new_n239), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n190), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n237), .A2(new_n239), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n189), .A2(G902), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(KEYINPUT78), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT78), .ZN(new_n250));
  INV_X1    g064(.A(new_n248), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n244), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n256), .A3(G143), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n225), .A2(G143), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n207), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n254), .A2(new_n256), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(new_n263), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n261), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  INV_X1    g084(.A(G137), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(G134), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(G134), .ZN(new_n273));
  INV_X1    g087(.A(G134), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT65), .A3(G137), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G131), .ZN(new_n277));
  INV_X1    g091(.A(G131), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n271), .A2(G134), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(G134), .B2(new_n271), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n274), .A2(KEYINPUT11), .A3(G137), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n278), .B(new_n280), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(KEYINPUT69), .B(new_n261), .C1(new_n262), .C2(new_n266), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n269), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OR2_X1    g101(.A1(KEYINPUT67), .A2(G116), .ZN(new_n288));
  NAND2_X1  g102(.A1(KEYINPUT67), .A2(G116), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(G119), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G116), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(G119), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT2), .B(G113), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n293), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n295), .B(new_n290), .C1(new_n291), .C2(G119), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(KEYINPUT0), .A2(G128), .ZN(new_n299));
  NOR2_X1   g113(.A1(KEYINPUT0), .A2(G128), .ZN(new_n300));
  OR2_X1    g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n255), .A2(G146), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n263), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n264), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n257), .A2(new_n259), .A3(new_n299), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT68), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT11), .B1(new_n274), .B2(G137), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n281), .A2(new_n271), .A3(G134), .ZN(new_n310));
  AOI211_X1 g124(.A(G131), .B(new_n279), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n310), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n278), .B1(new_n312), .B2(new_n280), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n299), .A2(new_n300), .ZN(new_n315));
  AOI21_X1  g129(.A(G143), .B1(new_n254), .B2(new_n256), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(new_n264), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n257), .A2(new_n259), .A3(new_n299), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n308), .A2(new_n314), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n287), .A2(new_n298), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n325));
  NOR2_X1   g139(.A1(G237), .A2(G953), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G210), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n325), .B(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT26), .B(G101), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n267), .A2(new_n285), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n317), .B(new_n319), .C1(new_n311), .C2(new_n313), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n298), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n318), .B1(new_n317), .B2(new_n319), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n297), .B1(new_n336), .B2(new_n314), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n333), .B1(new_n337), .B2(new_n287), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n324), .B(new_n330), .C1(new_n338), .C2(new_n323), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n287), .A2(KEYINPUT30), .A3(new_n321), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT66), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n331), .A2(new_n332), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT30), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI211_X1 g160(.A(KEYINPUT66), .B(KEYINPUT30), .C1(new_n331), .C2(new_n332), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n297), .B(new_n342), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n330), .B1(new_n348), .B2(new_n322), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n238), .B1(new_n341), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n298), .B1(new_n287), .B2(new_n321), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT71), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n322), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI211_X1 g167(.A(KEYINPUT71), .B(new_n298), .C1(new_n287), .C2(new_n321), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT28), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT72), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n322), .A2(new_n356), .A3(new_n323), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n322), .B2(new_n323), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n330), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(new_n340), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n355), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G472), .B1(new_n350), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT73), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n362), .B(new_n238), .C1(new_n349), .C2(new_n341), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT73), .A3(G472), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n348), .A2(new_n322), .A3(new_n330), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT31), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n348), .A2(KEYINPUT31), .A3(new_n322), .A4(new_n330), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n324), .B1(new_n338), .B2(new_n323), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n360), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT32), .ZN(new_n378));
  NOR2_X1   g192(.A1(G472), .A2(G902), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n372), .A2(new_n373), .B1(new_n375), .B2(new_n360), .ZN(new_n381));
  INV_X1    g195(.A(new_n379), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT32), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n253), .B1(new_n369), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G237), .ZN(new_n386));
  INV_X1    g200(.A(G953), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(G214), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n263), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n326), .A2(G143), .A3(G214), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT17), .A3(G131), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n326), .A2(G143), .A3(G214), .ZN(new_n393));
  AOI21_X1  g207(.A(G143), .B1(new_n326), .B2(G214), .ZN(new_n394));
  OAI21_X1  g208(.A(G131), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT17), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n389), .A2(new_n278), .A3(new_n390), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n201), .A2(new_n226), .A3(new_n392), .A4(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G113), .B(G122), .ZN(new_n400));
  INV_X1    g214(.A(G104), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n191), .A2(KEYINPUT76), .A3(G125), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n203), .B2(KEYINPUT76), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G146), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n205), .ZN(new_n406));
  NAND2_X1  g220(.A1(KEYINPUT18), .A2(G131), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n389), .A2(new_n390), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n391), .A2(KEYINPUT18), .A3(G131), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n399), .A2(new_n402), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT89), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n399), .A2(KEYINPUT89), .A3(new_n402), .A4(new_n410), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n399), .A2(new_n410), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n415), .B1(new_n402), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n238), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n418), .A2(G475), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT90), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n413), .A2(new_n414), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n395), .A2(new_n397), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n198), .B1(new_n404), .B2(KEYINPUT16), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n422), .B1(new_n423), .B2(new_n225), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n425), .A2(KEYINPUT19), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(KEYINPUT19), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n203), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT86), .B1(new_n404), .B2(KEYINPUT19), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT86), .A4(KEYINPUT19), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n204), .B(new_n428), .C1(new_n429), .C2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n424), .B1(new_n432), .B2(KEYINPUT88), .ZN(new_n433));
  INV_X1    g247(.A(new_n428), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT19), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT86), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI211_X1 g251(.A(new_n265), .B(new_n434), .C1(new_n437), .C2(new_n430), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT88), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n402), .B1(new_n441), .B2(new_n410), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n420), .B1(new_n421), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(G475), .A2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n410), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n445), .B1(new_n433), .B2(new_n440), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n415), .B(KEYINPUT90), .C1(new_n402), .C2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n443), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n424), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n438), .B2(new_n439), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n432), .A2(KEYINPUT88), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n410), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n402), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n455), .A2(new_n456), .B1(new_n413), .B2(new_n414), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n444), .A2(new_n458), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n457), .A2(KEYINPUT91), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT91), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n411), .A2(new_n412), .ZN(new_n462));
  INV_X1    g276(.A(new_n414), .ZN(new_n463));
  OAI22_X1  g277(.A1(new_n462), .A2(new_n463), .B1(new_n446), .B2(new_n402), .ZN(new_n464));
  INV_X1    g278(.A(new_n459), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n419), .B1(new_n451), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT9), .B(G234), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(G217), .A3(new_n387), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n288), .A2(G122), .A3(new_n289), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n291), .A2(G122), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G107), .ZN(new_n476));
  INV_X1    g290(.A(G107), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n477), .A3(new_n474), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n263), .A2(G128), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n207), .A2(G143), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n274), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT13), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT13), .B1(new_n263), .B2(G128), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n485), .A2(KEYINPUT92), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(KEYINPUT92), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n479), .B(new_n482), .C1(new_n274), .C2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n480), .A2(new_n481), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G134), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n482), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n475), .A2(KEYINPUT14), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT14), .ZN(new_n494));
  OAI21_X1  g308(.A(G107), .B1(new_n473), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n478), .B(new_n492), .C1(new_n493), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(KEYINPUT93), .A3(new_n496), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n472), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT93), .B1(new_n489), .B2(new_n496), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(new_n471), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n238), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G478), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(KEYINPUT15), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI221_X1 g321(.A(new_n238), .B1(KEYINPUT15), .B2(new_n505), .C1(new_n501), .C2(new_n503), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n507), .A2(KEYINPUT94), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT94), .B1(new_n507), .B2(new_n508), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n468), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G101), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n477), .A2(G104), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n401), .A2(G107), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT3), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n477), .A3(G104), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n518), .A2(new_n515), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT79), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT3), .B1(new_n401), .B2(G107), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n513), .A4(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n521), .A2(new_n518), .A3(new_n513), .A4(new_n515), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT79), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n516), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n269), .A2(KEYINPUT10), .A3(new_n286), .A4(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT4), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n521), .A2(new_n518), .A3(new_n515), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(G101), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n523), .A2(KEYINPUT79), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n523), .A2(KEYINPUT79), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n527), .A3(G101), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT80), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n528), .A2(KEYINPUT80), .A3(new_n527), .A4(G101), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n532), .A2(new_n537), .A3(new_n308), .A4(new_n320), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n522), .A2(new_n524), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n258), .B1(new_n204), .B2(G143), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n207), .B1(new_n305), .B2(KEYINPUT1), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n261), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n516), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT10), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n526), .A2(new_n538), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n314), .ZN(new_n548));
  INV_X1    g362(.A(new_n314), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n526), .A2(new_n538), .A3(new_n546), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(KEYINPUT81), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(G110), .B(G140), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n387), .A2(G227), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n552), .B(new_n553), .Z(new_n554));
  INV_X1    g368(.A(KEYINPUT81), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n547), .A2(new_n555), .A3(new_n314), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n551), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n544), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n525), .A2(new_n267), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n314), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT12), .ZN(new_n561));
  INV_X1    g375(.A(new_n554), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n563), .B(new_n314), .C1(new_n558), .C2(new_n559), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n561), .A2(new_n562), .A3(new_n550), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G469), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n238), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n551), .A2(new_n556), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n562), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n561), .A2(new_n550), .A3(new_n564), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n554), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(G469), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(G469), .A2(G902), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n568), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n233), .B1(new_n470), .B2(new_n238), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(G210), .B1(G237), .B2(G902), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n539), .A2(new_n543), .ZN(new_n581));
  INV_X1    g395(.A(G113), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n291), .A2(G119), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT5), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n292), .B2(new_n584), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n296), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n525), .A2(new_n296), .A3(new_n586), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(G110), .B(G122), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n591), .B(KEYINPUT8), .Z(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT84), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT84), .ZN(new_n595));
  AOI211_X1 g409(.A(new_n595), .B(new_n592), .C1(new_n588), .C2(new_n589), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n532), .A2(new_n537), .A3(new_n297), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n589), .A3(new_n591), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n267), .A2(new_n193), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n317), .A2(G125), .A3(new_n319), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n387), .A2(G224), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(KEYINPUT7), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(KEYINPUT7), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n599), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n238), .B1(new_n597), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n598), .A2(new_n589), .ZN(new_n609));
  INV_X1    g423(.A(new_n591), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(KEYINPUT6), .A3(new_n599), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n603), .B(KEYINPUT83), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n602), .B(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT6), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n615), .A3(new_n610), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n580), .B1(new_n608), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n581), .A2(new_n587), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n539), .A2(new_n543), .B1(new_n586), .B2(new_n296), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n593), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n595), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n590), .A2(KEYINPUT84), .A3(new_n593), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n607), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n579), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n618), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n387), .A2(G952), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n187), .B2(new_n386), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AOI211_X1 g446(.A(new_n238), .B(new_n387), .C1(G234), .C2(G237), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT21), .B(G898), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(G214), .B1(G237), .B2(G902), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT82), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n629), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n512), .A2(new_n578), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n385), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT95), .B(G101), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G3));
  INV_X1    g458(.A(new_n468), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n497), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n472), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n497), .A2(new_n646), .A3(new_n471), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(KEYINPUT33), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n505), .A2(G902), .ZN(new_n651));
  INV_X1    g465(.A(new_n500), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n471), .B1(new_n652), .B2(new_n502), .ZN(new_n653));
  INV_X1    g467(.A(new_n503), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT33), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT97), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT97), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n658), .B(KEYINPUT33), .C1(new_n653), .C2(new_n654), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n650), .B(new_n651), .C1(new_n657), .C2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT99), .B(G478), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n504), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n645), .A2(KEYINPUT100), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n665));
  INV_X1    g479(.A(new_n650), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n656), .B1(new_n501), .B2(new_n503), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n658), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n655), .A2(KEYINPUT97), .A3(new_n656), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n670), .A2(new_n651), .B1(new_n504), .B2(new_n661), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n665), .B1(new_n468), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n626), .A2(new_n627), .A3(new_n579), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n579), .B1(new_n626), .B2(new_n627), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n639), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT96), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT96), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n629), .A2(new_n678), .A3(new_n639), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n635), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n575), .A2(new_n252), .A3(new_n249), .A4(new_n577), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n381), .B2(G902), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n377), .A2(new_n379), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n673), .A2(new_n680), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT34), .B(G104), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G6));
  INV_X1    g502(.A(new_n511), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n443), .A2(new_n447), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n444), .A3(new_n449), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n419), .B1(new_n691), .B2(new_n451), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n685), .A2(new_n680), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT35), .B(G107), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G9));
  NOR2_X1   g510(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n231), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n247), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n245), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n684), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n641), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT37), .B(G110), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G12));
  AOI21_X1  g521(.A(new_n578), .B1(new_n369), .B2(new_n384), .ZN(new_n708));
  INV_X1    g522(.A(G900), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n632), .B1(new_n633), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n689), .A2(new_n692), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n701), .B1(new_n677), .B2(new_n679), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n708), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G128), .ZN(G30));
  XOR2_X1   g529(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n710), .B(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n575), .A2(new_n577), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n718), .B(KEYINPUT105), .Z(new_n719));
  INV_X1    g533(.A(KEYINPUT40), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n353), .A2(new_n354), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n238), .B1(new_n723), .B2(new_n330), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n348), .A2(new_n322), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n360), .ZN(new_n726));
  OAI21_X1  g540(.A(G472), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n727), .B(KEYINPUT103), .Z(new_n728));
  INV_X1    g542(.A(new_n384), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n629), .B(KEYINPUT38), .Z(new_n731));
  NOR3_X1   g545(.A1(new_n731), .A2(new_n638), .A3(new_n700), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n468), .A2(new_n511), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n721), .A2(new_n722), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n263), .ZN(G45));
  NOR3_X1   g550(.A1(new_n468), .A2(new_n671), .A3(new_n710), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n708), .A2(new_n713), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G146), .ZN(G48));
  AOI21_X1  g553(.A(new_n567), .B1(new_n566), .B2(new_n238), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n577), .A3(new_n568), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n385), .A2(new_n673), .A3(new_n680), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND4_X1  g560(.A1(new_n385), .A2(new_n680), .A3(new_n693), .A4(new_n743), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G116), .ZN(G18));
  NOR3_X1   g562(.A1(new_n512), .A2(new_n635), .A3(new_n701), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n742), .B1(new_n677), .B2(new_n679), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT73), .B1(new_n367), .B2(G472), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n367), .A2(KEYINPUT73), .A3(G472), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n384), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n749), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G119), .ZN(G21));
  NOR3_X1   g569(.A1(new_n468), .A2(new_n511), .A3(new_n635), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n372), .A2(new_n373), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n330), .B1(new_n355), .B2(new_n359), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n379), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n244), .A2(new_n251), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n682), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n677), .A2(new_n679), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n756), .A2(new_n761), .A3(new_n762), .A4(new_n743), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT106), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n750), .A2(KEYINPUT106), .A3(new_n761), .A4(new_n756), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G122), .ZN(G24));
  OAI21_X1  g582(.A(KEYINPUT91), .B1(new_n457), .B2(new_n459), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n464), .A2(new_n461), .A3(new_n465), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n448), .B2(new_n450), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n663), .B(new_n711), .C1(new_n772), .C2(new_n419), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n682), .A2(new_n759), .A3(new_n700), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n750), .ZN(new_n776));
  XOR2_X1   g590(.A(KEYINPUT107), .B(G125), .Z(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(G27));
  AND4_X1   g592(.A1(new_n639), .A2(new_n618), .A3(new_n628), .A4(new_n577), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n572), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n571), .A2(KEYINPUT109), .A3(new_n554), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n570), .A2(new_n781), .A3(G469), .A4(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n574), .B(KEYINPUT108), .Z(new_n784));
  NAND3_X1  g598(.A1(new_n568), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n779), .A2(new_n785), .A3(KEYINPUT42), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n753), .A2(new_n786), .A3(new_n760), .A4(new_n737), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n760), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n369), .B2(new_n384), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n779), .A2(new_n785), .A3(KEYINPUT42), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n773), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n793), .A3(KEYINPUT110), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT42), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n779), .A2(new_n785), .ZN(new_n796));
  INV_X1    g610(.A(new_n253), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n753), .A2(new_n796), .A3(new_n797), .A4(new_n737), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n789), .A2(new_n794), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(new_n278), .ZN(G33));
  NAND3_X1  g614(.A1(new_n385), .A2(new_n712), .A3(new_n796), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G134), .ZN(G36));
  NAND2_X1  g616(.A1(new_n570), .A2(new_n572), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n570), .A2(new_n781), .A3(KEYINPUT45), .A4(new_n782), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(G469), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n784), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n568), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n808), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(KEYINPUT46), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n810), .B1(new_n812), .B2(KEYINPUT111), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n811), .B2(KEYINPUT46), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n576), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n816), .A2(new_n717), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n468), .A2(new_n663), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT43), .Z(new_n819));
  AOI21_X1  g633(.A(new_n701), .B1(new_n682), .B2(new_n683), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n819), .A2(KEYINPUT44), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT44), .B1(new_n819), .B2(new_n820), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n629), .A2(new_n638), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G137), .ZN(G39));
  XNOR2_X1  g641(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n816), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT47), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n816), .B1(KEYINPUT112), .B2(new_n830), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n753), .A2(new_n797), .A3(new_n773), .A4(new_n824), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  XOR2_X1   g647(.A(KEYINPUT113), .B(G140), .Z(new_n834));
  XNOR2_X1  g648(.A(new_n833), .B(new_n834), .ZN(G42));
  NOR2_X1   g649(.A1(G952), .A2(G953), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT121), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n819), .A2(new_n632), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n824), .A2(new_n742), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n791), .A3(new_n839), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT48), .Z(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n750), .A3(new_n761), .ZN(new_n842));
  INV_X1    g656(.A(new_n673), .ZN(new_n843));
  INV_X1    g657(.A(new_n730), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n797), .A3(new_n632), .A4(new_n839), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n842), .B(new_n630), .C1(new_n843), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n838), .A2(new_n761), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n731), .A2(new_n638), .A3(new_n743), .ZN(new_n849));
  OR4_X1    g663(.A1(KEYINPUT119), .A2(new_n848), .A3(KEYINPUT50), .A4(new_n849), .ZN(new_n850));
  XOR2_X1   g664(.A(KEYINPUT119), .B(KEYINPUT50), .Z(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(new_n848), .B2(new_n849), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n838), .A2(new_n839), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(new_n774), .ZN(new_n854));
  OR3_X1    g668(.A1(new_n845), .A2(new_n645), .A3(new_n663), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n850), .A2(new_n852), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n829), .A2(new_n831), .ZN(new_n857));
  INV_X1    g671(.A(new_n568), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n740), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n576), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n848), .A2(new_n824), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n847), .B1(new_n863), .B2(KEYINPUT51), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n854), .A2(new_n855), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(KEYINPUT51), .A3(new_n850), .A4(new_n852), .ZN(new_n867));
  INV_X1    g681(.A(new_n861), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n868), .A2(KEYINPUT120), .ZN(new_n869));
  INV_X1    g683(.A(new_n862), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n868), .B2(KEYINPUT120), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n867), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n762), .A2(new_n733), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n785), .A2(new_n577), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n701), .A2(KEYINPUT117), .A3(new_n711), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n700), .B2(new_n710), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n875), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n730), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n776), .A3(new_n714), .A4(new_n738), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT52), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n714), .A2(new_n776), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n738), .A4(new_n880), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n507), .A2(new_n508), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n710), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n692), .A2(new_n700), .A3(new_n823), .A4(new_n888), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n708), .A2(new_n889), .B1(new_n775), .B2(new_n796), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n641), .B1(new_n385), .B2(new_n702), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n681), .A2(new_n684), .A3(new_n640), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n451), .A2(new_n467), .ZN(new_n893));
  INV_X1    g707(.A(new_n419), .ZN(new_n894));
  AND4_X1   g708(.A1(KEYINPUT115), .A2(new_n893), .A3(new_n894), .A4(new_n887), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT115), .B1(new_n468), .B2(new_n887), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT114), .B1(new_n468), .B2(new_n671), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT114), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n663), .B(new_n899), .C1(new_n772), .C2(new_n419), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n892), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n890), .A2(new_n891), .A3(new_n801), .A4(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n799), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n765), .A2(new_n766), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n744), .A2(new_n747), .A3(new_n754), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n883), .A2(new_n884), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT53), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n886), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n886), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n767), .A2(new_n744), .A3(new_n747), .A4(new_n754), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT116), .ZN(new_n914));
  NOR4_X1   g728(.A1(new_n913), .A2(new_n799), .A3(new_n903), .A4(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT116), .B1(new_n904), .B2(new_n907), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n911), .B1(new_n919), .B2(KEYINPUT118), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT118), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n917), .A2(new_n922), .A3(new_n918), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n917), .B1(new_n918), .B2(new_n909), .ZN(new_n925));
  INV_X1    g739(.A(new_n919), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT54), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n837), .B1(new_n873), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n859), .B(KEYINPUT49), .Z(new_n930));
  NAND4_X1  g744(.A1(new_n731), .A2(new_n760), .A3(new_n639), .A4(new_n577), .ZN(new_n931));
  OR4_X1    g745(.A1(new_n730), .A2(new_n930), .A3(new_n931), .A4(new_n818), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n929), .A2(new_n932), .ZN(G75));
  NAND2_X1  g747(.A1(new_n798), .A2(new_n795), .ZN(new_n934));
  INV_X1    g748(.A(new_n794), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT110), .B1(new_n791), .B2(new_n793), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n891), .A2(new_n902), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n890), .A2(new_n801), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n914), .B1(new_n940), .B2(new_n913), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n904), .A2(KEYINPUT116), .A3(new_n907), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n886), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT118), .B1(new_n943), .B2(KEYINPUT53), .ZN(new_n944));
  INV_X1    g758(.A(new_n911), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n923), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(G210), .A3(G902), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT56), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n612), .A2(new_n616), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n614), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n947), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n951), .B1(new_n947), .B2(new_n948), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n387), .A2(G952), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G51));
  XOR2_X1   g769(.A(new_n784), .B(KEYINPUT57), .Z(new_n956));
  AOI21_X1  g770(.A(new_n921), .B1(new_n920), .B2(new_n923), .ZN(new_n957));
  AND4_X1   g771(.A1(new_n921), .A2(new_n944), .A3(new_n923), .A4(new_n945), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n566), .ZN(new_n960));
  INV_X1    g774(.A(new_n807), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n946), .A2(G902), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n954), .B1(new_n960), .B2(new_n962), .ZN(G54));
  NAND4_X1  g777(.A1(new_n946), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n964));
  INV_X1    g778(.A(new_n690), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n965), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n954), .ZN(G60));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT59), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n670), .B1(new_n928), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n670), .A2(new_n971), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n946), .A2(KEYINPUT54), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n973), .B1(new_n924), .B2(new_n974), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n972), .A2(new_n954), .A3(new_n975), .ZN(G63));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT60), .Z(new_n978));
  NAND2_X1  g792(.A1(new_n946), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n246), .B(KEYINPUT122), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n954), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n946), .A2(new_n698), .A3(new_n978), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT61), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n981), .A2(KEYINPUT61), .A3(new_n982), .A4(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(G66));
  NAND2_X1  g802(.A1(new_n907), .A2(new_n938), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n387), .ZN(new_n990));
  INV_X1    g804(.A(G224), .ZN(new_n991));
  OAI21_X1  g805(.A(G953), .B1(new_n634), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n949), .B1(G898), .B2(new_n387), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT123), .Z(new_n995));
  XNOR2_X1  g809(.A(new_n993), .B(new_n995), .ZN(G69));
  NAND2_X1  g810(.A1(new_n883), .A2(new_n738), .ZN(new_n997));
  OR3_X1    g811(.A1(new_n735), .A2(KEYINPUT62), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n719), .A2(new_n385), .A3(new_n823), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n897), .A2(new_n901), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n1001), .B1(new_n817), .B2(new_n825), .ZN(new_n1002));
  OAI21_X1  g816(.A(KEYINPUT62), .B1(new_n735), .B2(new_n997), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n998), .A2(new_n1002), .A3(new_n833), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n387), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n342), .B1(new_n346), .B2(new_n347), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT124), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n437), .A2(new_n430), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n428), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1007), .B(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n387), .B1(G227), .B2(G900), .ZN(new_n1011));
  AOI22_X1  g825(.A1(new_n1005), .A2(new_n1010), .B1(KEYINPUT125), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1010), .B1(G900), .B2(G953), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n874), .A2(new_n791), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n817), .B1(new_n825), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n801), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n997), .A2(new_n799), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n833), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1013), .B1(new_n1018), .B2(G953), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1012), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1011), .A2(KEYINPUT125), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1020), .B(new_n1021), .Z(G72));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  INV_X1    g838(.A(KEYINPUT126), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n370), .A2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(new_n349), .Z(new_n1027));
  OAI211_X1 g841(.A(new_n1024), .B(new_n1027), .C1(new_n925), .C2(new_n926), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1024), .B1(new_n1018), .B2(new_n989), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1029), .A2(new_n360), .A3(new_n725), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1024), .B1(new_n1004), .B2(new_n989), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n954), .B1(new_n1031), .B2(new_n726), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1028), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT127), .ZN(new_n1034));
  XNOR2_X1  g848(.A(new_n1033), .B(new_n1034), .ZN(G57));
endmodule


