//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n211), .B(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n207), .ZN(new_n226));
  INV_X1    g0026(.A(new_n201), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n213), .B(new_n224), .C1(new_n226), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(new_n216), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(new_n225), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G223), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT66), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(KEYINPUT66), .A3(G1698), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n250), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n255), .ZN(new_n262));
  INV_X1    g0062(.A(G222), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n262), .A2(new_n263), .B1(new_n264), .B2(new_n259), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n249), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n225), .B1(KEYINPUT65), .B2(new_n247), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT65), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G33), .A3(G41), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n267), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n268), .B2(new_n270), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n271), .B1(new_n274), .B2(G226), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n266), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G200), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n278), .A2(KEYINPUT68), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(G190), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n225), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n207), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n285), .A2(new_n287), .B1(G150), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n203), .A2(G20), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n283), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n282), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n206), .A2(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(G50), .A3(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(G50), .B2(new_n292), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g0098(.A(new_n298), .B(KEYINPUT9), .Z(new_n299));
  NAND3_X1  g0099(.A1(new_n279), .A2(new_n280), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n278), .A2(KEYINPUT68), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n299), .A2(new_n280), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n304), .A2(new_n279), .A3(new_n305), .A4(new_n301), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n276), .A2(new_n308), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n309), .B1(G169), .B2(new_n276), .C1(new_n291), .C2(new_n297), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT67), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n294), .A2(G77), .A3(new_n295), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(G77), .B2(new_n292), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n285), .A2(new_n288), .B1(G20), .B2(G77), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT15), .B(G87), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n286), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n314), .B1(new_n317), .B2(new_n282), .ZN(new_n318));
  INV_X1    g0118(.A(G238), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n256), .B2(new_n260), .ZN(new_n320));
  INV_X1    g0120(.A(G107), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n262), .A2(new_n216), .B1(new_n321), .B2(new_n259), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n249), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n271), .B1(new_n274), .B2(G244), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n312), .B(new_n318), .C1(new_n326), .C2(new_n277), .ZN(new_n327));
  INV_X1    g0127(.A(new_n318), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n277), .B1(new_n323), .B2(new_n324), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT67), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n327), .B(new_n330), .C1(new_n331), .C2(new_n325), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n326), .A2(new_n308), .ZN(new_n333));
  INV_X1    g0133(.A(G169), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n325), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n328), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G68), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n293), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT12), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n338), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n264), .B2(new_n286), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT11), .A3(new_n282), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n294), .A2(G68), .A3(new_n295), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT11), .B1(new_n342), .B2(new_n282), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n274), .A2(KEYINPUT69), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n247), .A2(KEYINPUT65), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(new_n270), .A3(new_n246), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n272), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT69), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n350), .A2(new_n355), .A3(G238), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n216), .A2(G1698), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(G226), .B2(G1698), .ZN(new_n359));
  INV_X1    g0159(.A(G33), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n359), .A2(new_n254), .B1(new_n360), .B2(new_n217), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n271), .B1(new_n361), .B2(new_n249), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n356), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n357), .B1(new_n356), .B2(new_n362), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n349), .B(G169), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n365), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n363), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n366), .B1(new_n308), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n349), .B1(new_n368), .B2(G169), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n348), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(G200), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n347), .C1(new_n331), .C2(new_n368), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n257), .A2(new_n207), .A3(new_n258), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n338), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n288), .A2(G159), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT70), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n288), .A2(KEYINPUT70), .A3(G159), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g0185(.A(G58), .B(G68), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n375), .B1(new_n380), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT7), .B1(new_n254), .B2(new_n207), .ZN(new_n390));
  NOR4_X1   g0190(.A1(new_n252), .A2(new_n253), .A3(new_n377), .A4(G20), .ZN(new_n391));
  OAI21_X1  g0191(.A(G68), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n383), .A2(new_n384), .B1(new_n386), .B2(G20), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(KEYINPUT16), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n389), .A2(new_n394), .A3(new_n282), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n284), .B1(new_n206), .B2(G20), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(new_n294), .B1(new_n293), .B2(new_n284), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n352), .A2(G232), .A3(new_n272), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n352), .A2(G274), .A3(new_n273), .ZN(new_n400));
  INV_X1    g0200(.A(G87), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n360), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(G223), .A2(G1698), .ZN(new_n403));
  INV_X1    g0203(.A(G226), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n403), .B1(new_n404), .B2(G1698), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n402), .B1(new_n405), .B2(new_n259), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n399), .B(new_n400), .C1(new_n406), .C2(new_n248), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G169), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n308), .B2(new_n407), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n398), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT18), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n398), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT71), .ZN(new_n416));
  OR2_X1    g0216(.A1(G223), .A2(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n404), .A2(G1698), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n252), .C2(new_n253), .ZN(new_n419));
  INV_X1    g0219(.A(new_n402), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n271), .B1(new_n421), .B2(new_n249), .ZN(new_n422));
  AOI21_X1  g0222(.A(G200), .B1(new_n422), .B2(new_n399), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n248), .B1(new_n419), .B2(new_n420), .ZN(new_n424));
  NOR2_X1   g0224(.A1(G41), .A2(G45), .ZN(new_n425));
  OAI21_X1  g0225(.A(G232), .B1(new_n425), .B2(G1), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n270), .B2(new_n268), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n424), .A2(new_n427), .A3(new_n271), .A4(G190), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n416), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n407), .A2(new_n277), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n421), .A2(new_n249), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n431), .A2(new_n331), .A3(new_n400), .A4(new_n399), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(KEYINPUT71), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n429), .A2(new_n395), .A3(new_n397), .A4(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT72), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n397), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n392), .A2(new_n393), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n283), .B1(new_n441), .B2(new_n375), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n440), .B1(new_n442), .B2(new_n394), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n443), .A2(KEYINPUT72), .A3(new_n429), .A4(new_n433), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n415), .B(new_n437), .C1(new_n445), .C2(new_n435), .ZN(new_n446));
  NOR4_X1   g0246(.A1(new_n311), .A2(new_n337), .A3(new_n374), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n206), .A2(G33), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n292), .A2(new_n448), .A3(new_n225), .A4(new_n281), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT74), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G107), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n293), .B(new_n321), .C1(KEYINPUT80), .C2(KEYINPUT25), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT80), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT25), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n453), .B(new_n454), .C1(new_n292), .C2(G107), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n452), .B(new_n455), .C1(new_n453), .C2(new_n454), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n321), .A2(G20), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT23), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n459), .B(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n207), .B(G87), .C1(new_n252), .C2(new_n253), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n462), .A2(KEYINPUT22), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n462), .A2(KEYINPUT22), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n458), .B(new_n461), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT24), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n283), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n461), .A2(new_n458), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n468), .B(KEYINPUT24), .C1(new_n463), .C2(new_n464), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n457), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(G250), .A2(G1698), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n218), .B2(G1698), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n473), .A2(new_n259), .B1(G33), .B2(G294), .ZN(new_n474));
  OR2_X1    g0274(.A1(new_n474), .A2(new_n248), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n352), .A2(new_n481), .A3(G264), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n206), .A2(G45), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT5), .ZN(new_n484));
  INV_X1    g0284(.A(G41), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n483), .B1(new_n486), .B2(new_n478), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(new_n352), .A3(G274), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n475), .A2(KEYINPUT81), .A3(new_n482), .A4(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n482), .B(new_n488), .C1(new_n474), .C2(new_n248), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n489), .A2(G169), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n490), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G179), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n471), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(G190), .B1(new_n489), .B2(new_n492), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n494), .A2(G200), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n470), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT82), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT82), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n497), .A2(new_n503), .A3(new_n500), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n352), .A2(new_n481), .A3(G270), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n488), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(G257), .B(new_n255), .C1(new_n252), .C2(new_n253), .ZN(new_n508));
  OAI211_X1 g0308(.A(G264), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n509));
  INV_X1    g0309(.A(G303), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n259), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n249), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G116), .ZN(new_n514));
  OR2_X1    g0314(.A1(new_n449), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n293), .A2(new_n514), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n281), .A2(new_n225), .B1(G20), .B2(new_n514), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G283), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n518), .B(new_n207), .C1(G33), .C2(new_n217), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n517), .A2(KEYINPUT20), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT20), .B1(new_n517), .B2(new_n519), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n515), .B(new_n516), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n513), .A2(G169), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT21), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n512), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n488), .A2(new_n506), .ZN(new_n527));
  OAI21_X1  g0327(.A(G200), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n522), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n507), .A2(G190), .A3(new_n512), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n513), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(G179), .A3(new_n522), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n513), .A2(KEYINPUT21), .A3(G169), .A4(new_n522), .ZN(new_n534));
  AND4_X1   g0334(.A1(new_n525), .A2(new_n531), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(G244), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n536));
  OAI211_X1 g0336(.A(G238), .B(new_n255), .C1(new_n252), .C2(new_n253), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n536), .B(new_n537), .C1(new_n360), .C2(new_n514), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n249), .ZN(new_n539));
  AOI21_X1  g0339(.A(G250), .B1(new_n206), .B2(G45), .ZN(new_n540));
  INV_X1    g0340(.A(G274), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(new_n477), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n352), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n308), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT78), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n539), .A2(new_n543), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n334), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT78), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n539), .A2(new_n548), .A3(new_n308), .A4(new_n543), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n259), .A2(new_n207), .A3(G68), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n286), .B2(new_n217), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n401), .A2(new_n217), .A3(new_n321), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT79), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT79), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(new_n401), .A3(new_n217), .A4(new_n321), .ZN(new_n557));
  NAND3_X1  g0357(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n555), .A2(new_n557), .B1(new_n207), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n282), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT74), .ZN(new_n561));
  OR2_X1    g0361(.A1(new_n449), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n449), .A2(new_n561), .ZN(new_n563));
  INV_X1    g0363(.A(new_n316), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n316), .A2(new_n293), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n560), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n545), .A2(new_n547), .A3(new_n549), .A4(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n560), .A2(new_n566), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n546), .A2(G200), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n539), .A2(G190), .A3(new_n543), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n450), .A2(G87), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n569), .A2(new_n570), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n488), .ZN(new_n576));
  OAI211_X1 g0376(.A(G244), .B(new_n255), .C1(new_n252), .C2(new_n253), .ZN(new_n577));
  XNOR2_X1  g0377(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n255), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n259), .A2(G250), .A3(G1698), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n518), .A4(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n576), .B1(new_n582), .B2(new_n249), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n352), .A2(new_n481), .A3(G257), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n584), .B(KEYINPUT77), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n585), .A3(new_n308), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n583), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n334), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n217), .B1(new_n562), .B2(new_n563), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n292), .A2(new_n217), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT75), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT75), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n593), .B(new_n590), .C1(new_n450), .C2(new_n217), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(G107), .B1(new_n390), .B2(new_n391), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n288), .A2(G77), .ZN(new_n597));
  XNOR2_X1  g0397(.A(G97), .B(G107), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT73), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(KEYINPUT6), .ZN(new_n600));
  MUX2_X1   g0400(.A(new_n599), .B(G97), .S(KEYINPUT6), .Z(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n596), .B(new_n597), .C1(new_n207), .C2(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n603), .A2(new_n282), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n586), .B(new_n588), .C1(new_n595), .C2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n592), .A2(new_n594), .B1(new_n282), .B2(new_n603), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n587), .A2(G190), .ZN(new_n607));
  AOI21_X1  g0407(.A(G200), .B1(new_n583), .B2(new_n585), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n535), .A2(new_n575), .A3(new_n605), .A4(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n447), .A2(new_n505), .A3(new_n610), .ZN(G372));
  XNOR2_X1  g0411(.A(KEYINPUT86), .B(KEYINPUT26), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n605), .A2(new_n574), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT26), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT83), .B1(new_n542), .B2(new_n352), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n542), .A2(KEYINPUT83), .A3(new_n352), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n616), .A2(new_n617), .B1(new_n249), .B2(new_n538), .ZN(new_n618));
  OAI211_X1 g0418(.A(KEYINPUT84), .B(new_n544), .C1(new_n618), .C2(G169), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n617), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n539), .B1(new_n621), .B2(new_n615), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n334), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT84), .B1(new_n623), .B2(new_n544), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n567), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n588), .A2(new_n586), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(new_n606), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT85), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n622), .B2(G200), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n618), .A2(KEYINPUT85), .A3(new_n277), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n625), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n613), .B1(new_n614), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n605), .A2(new_n632), .A3(new_n609), .A4(new_n500), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n525), .A2(new_n533), .A3(new_n534), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n496), .B2(new_n471), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n625), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n447), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n435), .B1(new_n439), .B2(new_n444), .ZN(new_n641));
  INV_X1    g0441(.A(new_n336), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n373), .A2(new_n642), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n436), .B(new_n641), .C1(new_n643), .C2(new_n371), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n307), .B1(new_n644), .B2(new_n414), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(new_n310), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n646), .ZN(G369));
  NAND3_X1  g0447(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n649), .A2(new_n650), .A3(G213), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G343), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n505), .B1(new_n470), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n652), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n471), .A2(new_n496), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n522), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n535), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n636), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(KEYINPUT87), .B(G330), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n656), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n471), .A2(new_n496), .A3(new_n652), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n502), .A2(new_n504), .A3(new_n636), .A4(new_n652), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(G399));
  NAND3_X1  g0468(.A1(new_n555), .A2(new_n514), .A3(new_n557), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n210), .A2(new_n485), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n671), .A3(G1), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n228), .B2(new_n671), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT29), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n639), .A2(new_n675), .A3(new_n652), .ZN(new_n676));
  INV_X1    g0476(.A(new_n638), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n625), .A2(new_n627), .A3(KEYINPUT26), .A4(new_n632), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n612), .B1(new_n605), .B2(new_n574), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n654), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n676), .B1(new_n675), .B2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n610), .A2(new_n502), .A3(new_n504), .A4(new_n652), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n539), .A2(new_n543), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n474), .A2(new_n248), .ZN(new_n685));
  INV_X1    g0485(.A(new_n482), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n684), .A2(new_n583), .A3(new_n687), .A4(new_n585), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT88), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n513), .B2(new_n308), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n507), .A2(KEYINPUT88), .A3(new_n512), .A4(G179), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n689), .A2(KEYINPUT30), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n692), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n688), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n532), .A2(new_n618), .A3(G179), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n494), .B1(new_n583), .B2(new_n585), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT89), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n693), .B(new_n696), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n654), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n683), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n662), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n682), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n674), .B1(new_n710), .B2(G1), .ZN(G364));
  AOI21_X1  g0511(.A(new_n225), .B1(G20), .B2(new_n334), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n207), .A2(new_n331), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n308), .A2(G200), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n207), .A2(G190), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(G58), .A2(new_n717), .B1(new_n720), .B2(G77), .ZN(new_n721));
  NAND3_X1  g0521(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n331), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n721), .B1(new_n202), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT92), .Z(new_n726));
  NOR2_X1   g0526(.A1(new_n277), .A2(G179), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n714), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n259), .B1(new_n728), .B2(new_n401), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n718), .A2(new_n727), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n729), .B1(G107), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G179), .A2(G200), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n207), .B1(new_n733), .B2(G190), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n217), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n722), .A2(G190), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n736), .B2(G68), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n718), .A2(new_n733), .ZN(new_n738));
  INV_X1    g0538(.A(G159), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT32), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n726), .A2(new_n732), .A3(new_n737), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT93), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n254), .B1(new_n728), .B2(new_n510), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(G326), .B2(new_n723), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G322), .A2(new_n717), .B1(new_n731), .B2(G283), .ZN(new_n746));
  INV_X1    g0546(.A(new_n738), .ZN(new_n747));
  AOI22_X1  g0547(.A1(G311), .A2(new_n720), .B1(new_n747), .B2(G329), .ZN(new_n748));
  INV_X1    g0548(.A(new_n734), .ZN(new_n749));
  XNOR2_X1  g0549(.A(KEYINPUT33), .B(G317), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n749), .A2(G294), .B1(new_n736), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n745), .A2(new_n746), .A3(new_n748), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n743), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT94), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n713), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n754), .B2(new_n753), .ZN(new_n756));
  INV_X1    g0556(.A(new_n671), .ZN(new_n757));
  INV_X1    g0557(.A(G13), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n206), .B1(new_n759), .B2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n210), .A2(new_n259), .ZN(new_n763));
  INV_X1    g0563(.A(G355), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n763), .A2(new_n764), .B1(G116), .B2(new_n210), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n241), .A2(new_n476), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n210), .A2(new_n254), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n476), .B2(new_n229), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n765), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n712), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT90), .Z(new_n774));
  OAI21_X1  g0574(.A(new_n762), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT91), .ZN(new_n776));
  INV_X1    g0576(.A(new_n772), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n756), .B(new_n776), .C1(new_n660), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n664), .A2(new_n762), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n662), .B2(new_n660), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(G396));
  NOR2_X1   g0582(.A1(new_n336), .A2(new_n654), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n328), .A2(new_n654), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n332), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n783), .B1(new_n785), .B2(new_n336), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n786), .B(new_n652), .C1(new_n634), .C2(new_n638), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(KEYINPUT96), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n786), .B1(new_n639), .B2(new_n652), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n789), .B(new_n790), .Z(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n709), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n762), .B1(new_n791), .B2(new_n709), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(new_n793), .B2(KEYINPUT97), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(KEYINPUT97), .B2(new_n793), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n712), .A2(new_n770), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n761), .B(new_n757), .C1(new_n264), .C2(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G143), .A2(new_n717), .B1(new_n720), .B2(G159), .ZN(new_n798));
  INV_X1    g0598(.A(G137), .ZN(new_n799));
  INV_X1    g0599(.A(G150), .ZN(new_n800));
  INV_X1    g0600(.A(new_n736), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n798), .B1(new_n724), .B2(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT34), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n259), .B1(new_n730), .B2(new_n338), .ZN(new_n806));
  INV_X1    g0606(.A(G132), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n728), .A2(new_n202), .B1(new_n738), .B2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n806), .B(new_n808), .C1(G58), .C2(new_n749), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n804), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n254), .B1(new_n728), .B2(new_n321), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n735), .B(new_n811), .C1(G303), .C2(new_n723), .ZN(new_n812));
  INV_X1    g0612(.A(G294), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n716), .A2(new_n813), .B1(new_n719), .B2(new_n514), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n730), .A2(new_n401), .B1(new_n738), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G283), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n801), .A2(KEYINPUT95), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n801), .A2(KEYINPUT95), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n812), .B(new_n817), .C1(new_n818), .C2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n810), .A2(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n797), .B1(new_n713), .B2(new_n823), .C1(new_n786), .C2(new_n771), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n795), .A2(new_n824), .ZN(G384));
  INV_X1    g0625(.A(KEYINPUT35), .ZN(new_n826));
  OAI211_X1 g0626(.A(G116), .B(new_n226), .C1(new_n602), .C2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n826), .B2(new_n602), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT36), .Z(new_n829));
  OAI21_X1  g0629(.A(G77), .B1(new_n215), .B2(new_n338), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n228), .A2(new_n830), .B1(G50), .B2(new_n338), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n831), .A2(G1), .A3(new_n758), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT98), .Z(new_n834));
  INV_X1    g0634(.A(KEYINPUT100), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n395), .A2(new_n835), .A3(new_n397), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n395), .B2(new_n397), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n651), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n446), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n409), .B1(new_n836), .B2(new_n837), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n841), .A2(new_n838), .A3(new_n439), .A4(new_n444), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n398), .A2(new_n651), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n410), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n445), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT38), .B1(new_n840), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n439), .A2(new_n444), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n436), .B1(new_n851), .B2(KEYINPUT17), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n838), .B1(new_n852), .B2(new_n415), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n842), .A2(KEYINPUT37), .B1(new_n445), .B2(new_n847), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT102), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n840), .A2(KEYINPUT38), .A3(new_n849), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n855), .B1(new_n853), .B2(new_n854), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT102), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n347), .A2(new_n652), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT99), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n371), .B2(new_n373), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n371), .A2(new_n373), .A3(new_n864), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n702), .A2(KEYINPUT105), .A3(new_n654), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT105), .B1(new_n702), .B2(new_n654), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT31), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n683), .A2(new_n706), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n868), .B(new_n786), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT40), .B1(new_n862), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT104), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n641), .A2(new_n414), .A3(new_n436), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n877), .B2(new_n844), .ZN(new_n878));
  INV_X1    g0678(.A(new_n844), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n446), .A2(KEYINPUT104), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n434), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n846), .B1(new_n845), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n848), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n878), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n858), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n873), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n875), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n870), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n702), .A2(KEYINPUT105), .A3(new_n654), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(new_n704), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(new_n706), .A3(new_n683), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n447), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n662), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n890), .B2(new_n895), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n371), .A2(new_n654), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT39), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n856), .B1(new_n884), .B2(new_n885), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n899), .B(new_n900), .C1(new_n901), .C2(KEYINPUT39), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n371), .A2(new_n373), .A3(new_n864), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n903), .A2(new_n865), .ZN(new_n904));
  INV_X1    g0704(.A(new_n783), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n787), .B2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n860), .B1(new_n858), .B2(new_n859), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n651), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n414), .A2(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n902), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n682), .A2(new_n447), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n646), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n912), .B(new_n914), .Z(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n897), .A2(new_n916), .B1(new_n206), .B2(new_n759), .ZN(new_n917));
  INV_X1    g0717(.A(new_n897), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n915), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n834), .B1(new_n917), .B2(new_n919), .ZN(G367));
  OAI211_X1 g0720(.A(new_n605), .B(new_n609), .C1(new_n606), .C2(new_n652), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n627), .A2(new_n654), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n667), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT42), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n605), .B1(new_n921), .B2(new_n497), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n652), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n569), .A2(new_n572), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n654), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n625), .A2(new_n632), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n625), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT43), .B1(new_n933), .B2(KEYINPUT106), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(KEYINPUT106), .B2(new_n933), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n929), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n929), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n665), .A2(new_n924), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n938), .B(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n671), .B(KEYINPUT41), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n667), .A2(new_n666), .A3(new_n923), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT107), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(KEYINPUT107), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT45), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n923), .B1(new_n667), .B2(new_n666), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT108), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT44), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n948), .A2(new_n951), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(KEYINPUT108), .C2(KEYINPUT44), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n943), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n665), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n653), .B(new_n655), .C1(new_n659), .C2(new_n654), .ZN(new_n959));
  AOI211_X1 g0759(.A(KEYINPUT109), .B(new_n663), .C1(new_n959), .C2(new_n667), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n663), .A2(KEYINPUT109), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n663), .A2(KEYINPUT109), .ZN(new_n963));
  AND4_X1   g0763(.A1(new_n667), .A2(new_n959), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n710), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n956), .A2(new_n957), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n958), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n941), .B1(new_n969), .B2(new_n710), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n940), .B1(new_n970), .B2(new_n761), .ZN(new_n971));
  INV_X1    g0771(.A(new_n774), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n210), .B2(new_n316), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n237), .A2(new_n767), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n762), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n731), .A2(G77), .ZN(new_n976));
  INV_X1    g0776(.A(G143), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n976), .B(new_n259), .C1(new_n977), .C2(new_n724), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G68), .B2(new_n749), .ZN(new_n979));
  INV_X1    g0779(.A(new_n821), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(G159), .ZN(new_n981));
  INV_X1    g0781(.A(new_n728), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G58), .A2(new_n982), .B1(new_n717), .B2(G150), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G50), .A2(new_n720), .B1(new_n747), .B2(G137), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n979), .A2(new_n981), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n724), .A2(new_n815), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n259), .B(new_n986), .C1(G317), .C2(new_n747), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n321), .B2(new_n734), .C1(new_n821), .C2(new_n813), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT110), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n728), .B2(new_n514), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT46), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(KEYINPUT46), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n717), .A2(G303), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G97), .A2(new_n731), .B1(new_n720), .B2(G283), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n985), .B1(new_n988), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT47), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n975), .B1(new_n997), .B2(new_n712), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n933), .B2(new_n777), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n971), .A2(new_n999), .ZN(G387));
  INV_X1    g0800(.A(new_n965), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n653), .A2(new_n655), .A3(new_n772), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n670), .A2(new_n763), .B1(G107), .B2(new_n210), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n767), .B1(new_n234), .B2(G45), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n670), .A2(KEYINPUT111), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n670), .A2(KEYINPUT111), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n284), .A2(G50), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT50), .ZN(new_n1008));
  AOI21_X1  g0808(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1003), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n762), .B1(new_n1011), .B2(new_n774), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n734), .A2(new_n316), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n254), .B(new_n1013), .C1(G97), .C2(new_n731), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n723), .A2(G159), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT112), .Z(new_n1016));
  OAI22_X1  g0816(.A1(new_n202), .A2(new_n716), .B1(new_n728), .B2(new_n264), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n719), .A2(new_n338), .B1(new_n738), .B2(new_n800), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n285), .A2(new_n736), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1014), .A2(new_n1016), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n259), .B1(new_n747), .B2(G326), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n728), .A2(new_n813), .B1(new_n734), .B2(new_n818), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G317), .A2(new_n717), .B1(new_n720), .B2(G303), .ZN(new_n1024));
  INV_X1    g0824(.A(G322), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n724), .C1(new_n821), .C2(new_n815), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT48), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT49), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1022), .B1(new_n514), .B2(new_n730), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1021), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1012), .B1(new_n1033), .B2(new_n712), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1001), .A2(new_n761), .B1(new_n1002), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n757), .B1(new_n965), .B2(new_n966), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1001), .A2(new_n710), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(G393));
  NAND3_X1  g0838(.A1(new_n958), .A2(new_n761), .A3(new_n968), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n972), .B1(new_n217), .B2(new_n210), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n244), .A2(new_n767), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n762), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n980), .A2(G50), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n724), .A2(new_n800), .B1(new_n716), .B2(new_n739), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT51), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n728), .A2(new_n338), .B1(new_n738), .B2(new_n977), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n285), .B2(new_n720), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n734), .A2(new_n264), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n254), .B(new_n1048), .C1(G87), .C2(new_n731), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n719), .A2(new_n813), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n254), .B1(new_n730), .B2(new_n321), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(G116), .C2(new_n749), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n728), .A2(new_n818), .B1(new_n738), .B2(new_n1025), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT113), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(new_n821), .C2(new_n510), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n717), .A2(G311), .B1(G317), .B2(new_n723), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1050), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1042), .B1(new_n1059), .B2(new_n712), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n923), .B2(new_n777), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n969), .A2(new_n757), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n967), .B1(new_n968), .B2(new_n958), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1039), .B(new_n1061), .C1(new_n1062), .C2(new_n1063), .ZN(G390));
  INV_X1    g0864(.A(KEYINPUT115), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n787), .A2(new_n905), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n868), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1065), .B1(new_n1067), .B2(new_n898), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n906), .A2(KEYINPUT115), .A3(new_n899), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n900), .B1(new_n901), .B2(KEYINPUT39), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n785), .A2(new_n336), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n783), .B1(new_n681), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n898), .B1(new_n1074), .B2(new_n904), .ZN(new_n1075));
  OAI21_X1  g0875(.A(KEYINPUT114), .B1(new_n1075), .B2(new_n901), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n680), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n652), .B(new_n1073), .C1(new_n1077), .C2(new_n638), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n905), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n899), .B1(new_n1079), .B2(new_n868), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT114), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n887), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n868), .A2(new_n707), .A3(new_n662), .A4(new_n786), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1072), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1071), .A2(new_n1070), .B1(new_n1076), .B2(new_n1082), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n894), .A2(G330), .A3(new_n786), .A4(new_n868), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n786), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n904), .B1(new_n708), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n894), .A2(G330), .A3(new_n786), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n904), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1084), .A2(new_n1074), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1066), .A2(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n447), .A2(G330), .A3(new_n894), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n913), .A2(new_n646), .A3(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1088), .A2(KEYINPUT116), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT116), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .C1(new_n1098), .C2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1102), .A3(new_n757), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1085), .B(new_n761), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n796), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n762), .B1(new_n285), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n980), .A2(G137), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n734), .A2(new_n739), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n259), .B1(new_n730), .B2(new_n202), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(G128), .C2(new_n723), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n728), .A2(new_n800), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT53), .ZN(new_n1112));
  INV_X1    g0912(.A(G125), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n716), .A2(new_n807), .B1(new_n738), .B2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT54), .B(G143), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1114), .B1(new_n720), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1107), .A2(new_n1110), .A3(new_n1112), .A4(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n821), .A2(new_n321), .B1(new_n217), .B2(new_n719), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT117), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n716), .A2(new_n514), .B1(new_n730), .B2(new_n338), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G294), .B2(new_n747), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n254), .B1(new_n728), .B2(new_n401), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1048), .B(new_n1123), .C1(G283), .C2(new_n723), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1120), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1119), .A2(KEYINPUT117), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1118), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1106), .B1(new_n1127), .B2(new_n712), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1071), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n771), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1104), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1103), .A2(new_n1131), .ZN(G378));
  INV_X1    g0932(.A(KEYINPUT121), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n298), .A2(new_n910), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n311), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n307), .B(new_n310), .C1(new_n298), .C2(new_n910), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n894), .A2(KEYINPUT40), .A3(new_n786), .A4(new_n868), .ZN(new_n1143));
  OAI21_X1  g0943(.A(G330), .B1(new_n1143), .B2(new_n901), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1142), .B1(new_n875), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n874), .B1(new_n907), .B2(new_n908), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n888), .ZN(new_n1147));
  INV_X1    g0947(.A(G330), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n889), .B2(new_n887), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1145), .A2(new_n912), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n912), .B1(new_n1145), .B2(new_n1151), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1133), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n912), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n875), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1150), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1145), .A2(new_n1151), .A3(new_n912), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(KEYINPUT121), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1154), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1085), .B(new_n1098), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1097), .B(KEYINPUT122), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT57), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT57), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n757), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  AOI211_X1 g0970(.A(G41), .B(new_n259), .C1(new_n747), .C2(G283), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n215), .B2(new_n730), .C1(new_n264), .C2(new_n728), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT119), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n716), .A2(new_n321), .B1(new_n719), .B2(new_n316), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G68), .B2(new_n749), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n736), .A2(G97), .B1(new_n723), .B2(G116), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT58), .ZN(new_n1178));
  OR2_X1    g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(G33), .A2(G41), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT118), .Z(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(new_n202), .C1(G41), .C2(new_n259), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1179), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n801), .A2(new_n807), .B1(new_n800), .B2(new_n734), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G128), .A2(new_n717), .B1(new_n982), .B2(new_n1116), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n799), .B2(new_n719), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G125), .C2(new_n723), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1182), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G159), .A2(new_n731), .B1(new_n747), .B2(G124), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n713), .B1(new_n1184), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n762), .B1(G50), .B2(new_n1105), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n1142), .C2(new_n770), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT120), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1161), .B2(new_n761), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1170), .A2(new_n1199), .ZN(G375));
  AND2_X1   g1000(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT123), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n941), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT123), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1202), .A2(new_n1203), .A3(new_n1099), .A4(new_n1206), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(KEYINPUT124), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(KEYINPUT124), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1095), .A2(new_n760), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n259), .B1(new_n730), .B2(new_n215), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G50), .B2(new_n749), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G150), .A2(new_n720), .B1(new_n747), .B2(G128), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n739), .C2(new_n728), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT125), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n717), .A2(G137), .B1(G132), .B2(new_n723), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n821), .B2(new_n1115), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n980), .A2(G116), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1013), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n723), .A2(G294), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1221), .A2(new_n976), .A3(new_n254), .A4(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n217), .A2(new_n728), .B1(new_n716), .B2(new_n818), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n719), .A2(new_n321), .B1(new_n738), .B2(new_n510), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1216), .A2(new_n1219), .B1(new_n1220), .B2(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n762), .B1(G68), .B2(new_n1105), .C1(new_n1227), .C2(new_n713), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n904), .B2(new_n770), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1210), .A2(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT126), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1208), .A2(new_n1209), .A3(new_n1231), .ZN(G381));
  AND2_X1   g1032(.A1(new_n1103), .A2(new_n1131), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1170), .A2(new_n1233), .A3(new_n1199), .ZN(new_n1234));
  OR2_X1    g1034(.A1(G393), .A2(G396), .ZN(new_n1235));
  OR4_X1    g1035(.A1(G384), .A2(G387), .A3(new_n1235), .A4(G390), .ZN(new_n1236));
  OR3_X1    g1036(.A1(new_n1234), .A2(new_n1236), .A3(G381), .ZN(G407));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(G343), .C2(new_n1234), .ZN(G409));
  AOI21_X1  g1038(.A(G390), .B1(new_n971), .B2(new_n999), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(G393), .B(new_n781), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n971), .A2(new_n999), .A3(G390), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1241), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1242), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1244), .B1(new_n1245), .B2(new_n1239), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G378), .B(new_n1199), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1152), .A2(new_n1153), .A3(new_n1133), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT121), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1203), .B(new_n1164), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1197), .B1(new_n1167), .B2(new_n761), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1233), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1248), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(G343), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(G213), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1257), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(G2897), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1202), .B(new_n1206), .C1(new_n1262), .C2(new_n1098), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n671), .B1(new_n1201), .B2(KEYINPUT60), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1265), .A2(G384), .A3(new_n1231), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G384), .B1(new_n1265), .B2(new_n1231), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1261), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1231), .ZN(new_n1269));
  INV_X1    g1069(.A(G384), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1265), .A2(new_n1231), .A3(G384), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(new_n1260), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1268), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT61), .B1(new_n1258), .B2(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1255), .A2(new_n1257), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT62), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1277), .A2(KEYINPUT62), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1247), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1266), .A2(new_n1267), .A3(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1255), .A2(new_n1257), .A3(new_n1283), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1259), .B1(new_n1248), .B2(new_n1254), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT63), .B1(new_n1287), .B2(new_n1276), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT127), .B1(new_n1289), .B2(new_n1275), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1277), .A2(new_n1282), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1247), .B1(new_n1287), .B2(new_n1283), .ZN(new_n1292));
  AND4_X1   g1092(.A1(KEYINPUT127), .A2(new_n1275), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1281), .B1(new_n1290), .B2(new_n1293), .ZN(G405));
  AOI21_X1  g1094(.A(G378), .B1(new_n1170), .B2(new_n1199), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1248), .ZN(new_n1296));
  OR3_X1    g1096(.A1(new_n1295), .A2(new_n1296), .A3(new_n1276), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1276), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(new_n1247), .ZN(G402));
endmodule


