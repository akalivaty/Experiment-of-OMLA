//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT64), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G134), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  OAI211_X1 g008(.A(KEYINPUT64), .B(new_n194), .C1(new_n188), .C2(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n190), .A2(new_n198), .A3(new_n193), .A4(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT0), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(G143), .B(G146), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n206), .B2(new_n207), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n200), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G128), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n219), .B1(G143), .B2(new_n201), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n205), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n202), .A2(new_n204), .A3(new_n219), .A4(G128), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n188), .A2(G137), .ZN(new_n224));
  OAI21_X1  g038(.A(G131), .B1(new_n192), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n199), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n214), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G113), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT2), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G116), .B(G119), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G116), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT2), .B(G113), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n235), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT67), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n234), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n227), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n187), .B1(new_n246), .B2(KEYINPUT28), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n223), .A2(new_n199), .A3(new_n225), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n200), .B2(new_n213), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n244), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(KEYINPUT69), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n214), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n200), .A2(KEYINPUT65), .A3(new_n213), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n226), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n246), .B1(new_n245), .B2(new_n256), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n247), .B(new_n252), .C1(new_n257), .C2(new_n251), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT68), .A2(G953), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT68), .A2(G953), .ZN(new_n260));
  OR2_X1    g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G237), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(G210), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(G101), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n214), .A2(KEYINPUT30), .A3(new_n226), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n269), .B1(new_n256), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n246), .B1(new_n271), .B2(new_n245), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT31), .B1(new_n272), .B2(new_n266), .ZN(new_n273));
  INV_X1    g087(.A(new_n269), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n200), .A2(KEYINPUT65), .A3(new_n213), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT65), .B1(new_n200), .B2(new_n213), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n275), .A2(new_n276), .A3(new_n248), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n245), .B(new_n274), .C1(new_n277), .C2(KEYINPUT30), .ZN(new_n278));
  AND4_X1   g092(.A1(KEYINPUT31), .A2(new_n278), .A3(new_n250), .A4(new_n266), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n268), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(G472), .A2(G902), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n280), .A2(KEYINPUT32), .A3(new_n281), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT32), .B1(new_n280), .B2(new_n281), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OR2_X1    g101(.A1(new_n258), .A2(KEYINPUT29), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n266), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n272), .A2(new_n267), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT29), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n227), .A2(new_n245), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n250), .A2(KEYINPUT71), .A3(new_n292), .ZN(new_n293));
  OR3_X1    g107(.A1(new_n249), .A2(KEYINPUT71), .A3(new_n244), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(new_n251), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n247), .A2(new_n252), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n288), .A2(new_n266), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G472), .B1(new_n291), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT32), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n287), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(G101), .ZN(new_n306));
  INV_X1    g120(.A(G107), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G104), .ZN(new_n308));
  INV_X1    g122(.A(G104), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT3), .B1(new_n309), .B2(G107), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT74), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n312), .B(KEYINPUT3), .C1(new_n309), .C2(G107), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n308), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n307), .A3(G104), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n315), .A2(new_n307), .A3(KEYINPUT75), .A4(G104), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n306), .B1(new_n314), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n244), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n308), .ZN(new_n324));
  INV_X1    g138(.A(new_n313), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n307), .A2(G104), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n312), .B1(new_n326), .B2(KEYINPUT3), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n324), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n318), .A2(new_n319), .ZN(new_n329));
  OAI21_X1  g143(.A(G101), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n311), .A2(new_n313), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n331), .A2(new_n320), .A3(new_n306), .A4(new_n324), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(KEYINPUT4), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n323), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n324), .A2(new_n326), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G101), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n242), .A2(new_n243), .ZN(new_n338));
  INV_X1    g152(.A(new_n237), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n228), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n233), .A2(KEYINPUT5), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n342), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n337), .A2(new_n338), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n334), .A2(new_n347), .ZN(new_n348));
  XOR2_X1   g162(.A(G110), .B(G122), .Z(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n351));
  INV_X1    g165(.A(new_n349), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n334), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n350), .A2(new_n351), .A3(new_n353), .A4(KEYINPUT6), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n334), .A2(new_n347), .A3(new_n352), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n352), .B1(new_n334), .B2(new_n347), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT6), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n348), .A2(new_n357), .A3(new_n349), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT80), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n354), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G125), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n223), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n213), .A2(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G953), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G224), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(G224), .A3(new_n367), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n361), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT7), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n369), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n366), .A2(new_n374), .A3(new_n368), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n343), .B(KEYINPUT81), .ZN(new_n379));
  INV_X1    g193(.A(new_n341), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n338), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n337), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n349), .B(KEYINPUT8), .Z(new_n383));
  NAND2_X1  g197(.A1(new_n346), .A2(new_n338), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n382), .B(new_n383), .C1(new_n337), .C2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n378), .A2(new_n353), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n373), .A2(new_n300), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G210), .B1(G237), .B2(G902), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(G902), .B1(new_n361), .B2(new_n372), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n388), .A3(new_n386), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(G214), .B(new_n262), .C1(new_n259), .C2(new_n260), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n394), .A2(new_n203), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n203), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n198), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT17), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n198), .A3(new_n396), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n362), .A2(G140), .ZN(new_n402));
  XNOR2_X1  g216(.A(G125), .B(G140), .ZN(new_n403));
  MUX2_X1   g217(.A(new_n402), .B(new_n403), .S(KEYINPUT16), .Z(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(new_n201), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n395), .A2(new_n396), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT17), .A3(G131), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n397), .A2(KEYINPUT84), .A3(KEYINPUT17), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n401), .A2(new_n406), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT18), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n413), .A2(new_n198), .A3(KEYINPUT82), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT83), .B1(new_n403), .B2(new_n201), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n403), .A2(new_n201), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n414), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n395), .A2(new_n396), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n415), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n412), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G113), .B(G122), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(new_n309), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT86), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n300), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n422), .A2(new_n426), .ZN(new_n429));
  OAI21_X1  g243(.A(G475), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n404), .A2(new_n201), .ZN(new_n432));
  INV_X1    g246(.A(new_n403), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT19), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n403), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n436), .A3(new_n201), .ZN(new_n437));
  INV_X1    g251(.A(new_n400), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n432), .B(new_n437), .C1(new_n438), .C2(new_n397), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n439), .A2(new_n421), .A3(new_n425), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n422), .B2(new_n424), .ZN(new_n441));
  NOR2_X1   g255(.A1(G475), .A2(G902), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT85), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n431), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n425), .B1(new_n412), .B2(new_n421), .ZN(new_n446));
  NOR4_X1   g260(.A1(new_n446), .A2(KEYINPUT20), .A3(new_n440), .A4(new_n443), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n430), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT66), .B(G128), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT87), .B1(new_n450), .B2(new_n203), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n218), .A2(new_n452), .A3(G143), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n203), .A2(G128), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT13), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n449), .B(G134), .C1(new_n455), .C2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n453), .B2(new_n451), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT88), .B1(new_n460), .B2(new_n188), .ZN(new_n461));
  XNOR2_X1  g275(.A(G116), .B(G122), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(G107), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n451), .A2(new_n453), .B1(G128), .B2(new_n203), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n464), .B2(new_n188), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n238), .A2(G122), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n307), .B1(new_n467), .B2(KEYINPUT14), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n468), .A2(new_n470), .B1(new_n307), .B2(new_n462), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n464), .A2(new_n188), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n454), .A2(new_n188), .A3(new_n456), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n466), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT89), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n466), .A2(new_n474), .A3(KEYINPUT89), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT9), .B(G234), .Z(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G217), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n480), .A2(new_n481), .A3(G953), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n475), .A2(new_n476), .A3(new_n482), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n300), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G478), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(KEYINPUT15), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n488), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n484), .A2(new_n300), .A3(new_n485), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n367), .A2(G952), .ZN(new_n493));
  INV_X1    g307(.A(G234), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n493), .B1(new_n494), .B2(new_n262), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT21), .B(G898), .Z(new_n497));
  AOI21_X1  g311(.A(new_n300), .B1(G234), .B2(G237), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n261), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n448), .A2(new_n492), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n210), .A2(new_n212), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n321), .B2(new_n322), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n333), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n200), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n332), .A2(KEYINPUT10), .A3(new_n223), .A4(new_n336), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT76), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n222), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n211), .A2(KEYINPUT76), .A3(new_n219), .A4(G128), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n205), .B1(new_n220), .B2(new_n207), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n332), .A2(new_n513), .A3(new_n336), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT77), .B(KEYINPUT10), .Z(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n506), .A2(new_n507), .A3(new_n508), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n261), .A2(G227), .ZN(new_n518));
  XNOR2_X1  g332(.A(G110), .B(G140), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT78), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n506), .A2(new_n508), .A3(new_n516), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n200), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n517), .A2(KEYINPUT78), .A3(new_n520), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n520), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n514), .B1(new_n337), .B2(new_n223), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT12), .B1(new_n529), .B2(new_n200), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n332), .A2(new_n513), .A3(new_n336), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n223), .B1(new_n332), .B2(new_n336), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT12), .B(new_n200), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n517), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n528), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n527), .A2(G469), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G469), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(new_n300), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n535), .A2(new_n521), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n520), .B1(new_n525), .B2(new_n517), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n539), .B(new_n300), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n538), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(G221), .B1(new_n480), .B2(G902), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AND4_X1   g362(.A1(new_n305), .A2(new_n393), .A3(new_n503), .A4(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n236), .A2(KEYINPUT23), .A3(G128), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n207), .A2(G119), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n551), .B1(new_n218), .B2(G119), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n552), .B2(KEYINPUT23), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(G110), .ZN(new_n554));
  XOR2_X1   g368(.A(KEYINPUT24), .B(G110), .Z(new_n555));
  NOR2_X1   g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  OAI221_X1 g370(.A(new_n432), .B1(G146), .B2(new_n433), .C1(new_n554), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n552), .A2(new_n555), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(G110), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n405), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n261), .A2(G221), .A3(G234), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(G137), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT72), .B(KEYINPUT22), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n563), .B(new_n564), .Z(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n563), .B(new_n564), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n560), .A3(new_n557), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n481), .B1(G234), .B2(new_n300), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(G902), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n568), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n567), .B1(new_n557), .B2(new_n560), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT25), .B(new_n300), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT73), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT25), .B1(new_n569), .B2(new_n300), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT25), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n573), .A2(new_n574), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n570), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n572), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n304), .A2(new_n549), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  NAND3_X1  g401(.A1(new_n390), .A2(KEYINPUT90), .A3(new_n392), .ZN(new_n588));
  INV_X1    g402(.A(new_n305), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n388), .B1(new_n391), .B2(new_n386), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT90), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n278), .A2(new_n250), .A3(new_n266), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT31), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n272), .A2(KEYINPUT31), .A3(new_n266), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n597), .A2(new_n598), .B1(new_n267), .B2(new_n258), .ZN(new_n599));
  OAI21_X1  g413(.A(G472), .B1(new_n599), .B2(G902), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n282), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n601), .A2(new_n584), .A3(new_n547), .ZN(new_n602));
  INV_X1    g416(.A(new_n502), .ZN(new_n603));
  INV_X1    g417(.A(new_n448), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n484), .A2(new_n605), .A3(new_n485), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT91), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n475), .A2(KEYINPUT92), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(new_n483), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT33), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n607), .A2(G478), .A3(new_n300), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT93), .B(G478), .Z(new_n612));
  NAND2_X1  g426(.A1(new_n486), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n604), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n594), .A2(new_n602), .A3(new_n603), .A4(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(new_n615), .B(KEYINPUT94), .Z(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT34), .B(G104), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  OR3_X1    g432(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT95), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT95), .B1(new_n445), .B2(new_n447), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n430), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n489), .A2(new_n491), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n502), .B(KEYINPUT96), .Z(new_n623));
  NOR3_X1   g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n594), .A2(new_n602), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  INV_X1    g441(.A(new_n601), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n567), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(new_n561), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n571), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n578), .B2(new_n583), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n549), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  INV_X1    g449(.A(G900), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n501), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n499), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n638), .A2(KEYINPUT97), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(KEYINPUT97), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n495), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n621), .A2(new_n622), .A3(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n582), .A2(new_n570), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n576), .A2(new_n577), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n644), .A2(new_n645), .B1(new_n571), .B2(new_n630), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n547), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n304), .A2(new_n594), .A3(new_n643), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  XNOR2_X1  g463(.A(new_n641), .B(KEYINPUT39), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n548), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n646), .B1(new_n651), .B2(KEYINPUT40), .ZN(new_n652));
  AOI211_X1 g466(.A(new_n589), .B(new_n652), .C1(KEYINPUT40), .C2(new_n651), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n295), .A2(new_n267), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n300), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n272), .A2(new_n267), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n287), .A2(new_n303), .A3(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n658), .A2(KEYINPUT98), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(KEYINPUT98), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n604), .A2(new_n622), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n393), .B(KEYINPUT38), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n653), .A2(new_n662), .A3(new_n663), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  NAND2_X1  g480(.A1(new_n611), .A2(new_n613), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n448), .A3(new_n641), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n669), .A2(new_n304), .A3(new_n594), .A4(new_n647), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G146), .ZN(G48));
  OR2_X1    g485(.A1(new_n542), .A2(new_n543), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n539), .A2(KEYINPUT99), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n672), .A2(new_n300), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n672), .B2(new_n300), .ZN(new_n675));
  INV_X1    g489(.A(new_n546), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AND4_X1   g491(.A1(new_n603), .A2(new_n588), .A3(new_n592), .A4(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n678), .A2(new_n304), .A3(new_n585), .A4(new_n614), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  AND3_X1   g495(.A1(new_n588), .A2(new_n592), .A3(new_n677), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n304), .A2(new_n682), .A3(new_n585), .A4(new_n624), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G116), .ZN(G18));
  AND2_X1   g498(.A1(new_n503), .A2(new_n632), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n304), .A2(new_n594), .A3(new_n677), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G119), .ZN(G21));
  AND3_X1   g501(.A1(new_n588), .A2(new_n592), .A3(new_n663), .ZN(new_n688));
  INV_X1    g502(.A(G472), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n280), .B2(new_n300), .ZN(new_n690));
  INV_X1    g504(.A(new_n281), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n597), .A2(new_n598), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n267), .B1(new_n296), .B2(new_n297), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR4_X1   g508(.A1(new_n584), .A2(new_n690), .A3(new_n623), .A4(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n688), .A2(new_n677), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT100), .B(G122), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G24));
  OR2_X1    g512(.A1(new_n690), .A2(new_n694), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n646), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n614), .A2(KEYINPUT101), .A3(new_n641), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT101), .B1(new_n614), .B2(new_n641), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n682), .B(new_n700), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  NAND3_X1  g519(.A1(new_n390), .A2(new_n305), .A3(new_n392), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT103), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n390), .A2(new_n708), .A3(new_n305), .A4(new_n392), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n545), .A2(KEYINPUT102), .A3(new_n546), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT102), .B1(new_n545), .B2(new_n546), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n707), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n707), .A2(new_n712), .A3(KEYINPUT104), .A4(new_n709), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT101), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n668), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n701), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n285), .A2(new_n286), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n584), .B1(new_n302), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n717), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT42), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n304), .A2(new_n585), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n715), .B2(new_n716), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n720), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n643), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G134), .ZN(G36));
  NAND2_X1  g546(.A1(new_n667), .A2(new_n604), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT43), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT43), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n667), .A2(new_n735), .A3(new_n604), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n734), .A2(new_n601), .A3(new_n632), .A4(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n707), .A2(new_n709), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n745));
  INV_X1    g559(.A(new_n537), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n527), .A2(KEYINPUT45), .A3(new_n537), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(G469), .A3(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n749), .A2(KEYINPUT105), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(KEYINPUT105), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n540), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n544), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n752), .B2(KEYINPUT46), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n676), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n650), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n743), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n191), .ZN(G39));
  XOR2_X1   g574(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n761));
  NAND2_X1  g575(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n544), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n546), .B(new_n761), .C1(new_n763), .C2(new_n753), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT106), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n764), .B(new_n669), .C1(new_n757), .C2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n304), .A2(new_n585), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(KEYINPUT107), .A3(new_n742), .A4(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n546), .B1(new_n763), .B2(new_n753), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n766), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n669), .A3(new_n742), .A4(new_n764), .ZN(new_n775));
  INV_X1    g589(.A(new_n770), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n771), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n679), .A2(new_n683), .A3(new_n686), .A4(new_n696), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n782));
  INV_X1    g596(.A(new_n623), .ZN(new_n783));
  INV_X1    g597(.A(new_n392), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n305), .B(new_n783), .C1(new_n784), .C2(new_n590), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n492), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n489), .A2(KEYINPUT110), .A3(new_n491), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n448), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n782), .B1(new_n785), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n589), .B1(new_n390), .B2(new_n392), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(KEYINPUT111), .A3(new_n783), .A4(new_n789), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n602), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n602), .A2(new_n792), .A3(new_n614), .A4(new_n783), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n794), .A2(new_n586), .A3(new_n633), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n781), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n724), .A3(new_n728), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n699), .A2(new_n646), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n719), .B2(new_n701), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n717), .A2(new_n800), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n646), .A2(new_n621), .A3(new_n547), .A4(new_n642), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n304), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n742), .A3(new_n788), .A4(new_n787), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n643), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n806), .B(new_n725), .C1(new_n715), .C2(new_n716), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT112), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n731), .A2(new_n801), .A3(new_n809), .A4(new_n804), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n798), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n646), .A2(new_n548), .A3(new_n641), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n688), .A3(new_n658), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n704), .A2(new_n648), .A3(new_n815), .A4(new_n670), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT53), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n808), .A2(new_n810), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n797), .A2(new_n724), .A3(new_n728), .ZN(new_n821));
  AND4_X1   g635(.A1(KEYINPUT53), .A2(new_n820), .A3(new_n818), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n780), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n820), .A2(new_n821), .ZN(new_n825));
  INV_X1    g639(.A(new_n818), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n811), .A2(KEYINPUT53), .A3(new_n818), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n823), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n734), .A2(new_n736), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n831), .A2(new_n496), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n832), .A2(new_n677), .A3(new_n742), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n833), .A2(new_n722), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT48), .ZN(new_n836));
  INV_X1    g650(.A(new_n614), .ZN(new_n837));
  INV_X1    g651(.A(new_n677), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n741), .A2(new_n584), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n661), .A2(new_n496), .A3(new_n839), .ZN(new_n840));
  XOR2_X1   g654(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n841));
  OAI221_X1 g655(.A(new_n493), .B1(new_n837), .B2(new_n840), .C1(new_n834), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n674), .A2(new_n675), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT109), .Z(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n546), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n774), .A2(new_n764), .B1(KEYINPUT114), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(KEYINPUT114), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n699), .A2(new_n584), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n831), .A2(new_n496), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n741), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT51), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n849), .A2(new_n305), .A3(new_n838), .ZN(new_n852));
  INV_X1    g666(.A(new_n664), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT50), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n852), .A2(new_n856), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n833), .A2(new_n700), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OR3_X1    g673(.A1(new_n840), .A2(new_n448), .A3(new_n667), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n851), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n855), .A2(new_n860), .A3(new_n857), .A4(new_n858), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n845), .B1(new_n774), .B2(new_n764), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n863), .A2(new_n741), .A3(new_n849), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT51), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n842), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n830), .A2(new_n836), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n849), .A2(new_n593), .A3(new_n838), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n867), .A2(new_n868), .B1(G952), .B2(G953), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n844), .B(KEYINPUT49), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n664), .A3(new_n733), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n584), .A2(new_n589), .A3(new_n676), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT108), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n871), .A2(new_n661), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n869), .A2(new_n874), .ZN(G75));
  AOI21_X1  g689(.A(new_n300), .B1(new_n827), .B2(new_n828), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(G210), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT56), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n361), .B(new_n371), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT55), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n877), .B2(new_n878), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n261), .A2(G952), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G51));
  XNOR2_X1  g698(.A(new_n540), .B(KEYINPUT57), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n823), .A2(new_n829), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n823), .A2(new_n829), .A3(KEYINPUT116), .A4(new_n885), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n672), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n750), .A2(new_n751), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n876), .A2(KEYINPUT117), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT117), .B1(new_n876), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n883), .B1(new_n890), .B2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n876), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  INV_X1    g711(.A(new_n441), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n883), .ZN(G60));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT59), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n823), .A2(new_n829), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n607), .A2(new_n610), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n883), .ZN(G63));
  NAND2_X1  g722(.A1(new_n827), .A2(new_n828), .ZN(new_n909));
  XNOR2_X1  g723(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n481), .A2(new_n300), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n581), .ZN(new_n914));
  INV_X1    g728(.A(new_n883), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n630), .B(KEYINPUT119), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n909), .A2(new_n912), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n914), .A2(KEYINPUT61), .A3(new_n915), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(G66));
  AOI21_X1  g736(.A(new_n367), .B1(new_n497), .B2(G224), .ZN(new_n923));
  INV_X1    g737(.A(new_n797), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n261), .ZN(new_n925));
  INV_X1    g739(.A(new_n361), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(G898), .B2(new_n261), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT120), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n925), .B(new_n928), .ZN(G69));
  INV_X1    g743(.A(new_n778), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n704), .A2(new_n648), .A3(new_n670), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n743), .B2(new_n758), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT123), .ZN(new_n933));
  INV_X1    g747(.A(new_n758), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n722), .A2(new_n688), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n807), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n937), .B(new_n931), .C1(new_n743), .C2(new_n758), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n933), .A2(new_n729), .A3(new_n936), .A4(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n261), .B1(new_n930), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n637), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n434), .A2(new_n436), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n271), .B(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n665), .A2(new_n931), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n759), .B1(new_n946), .B2(KEYINPUT62), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n651), .B1(new_n837), .B2(new_n790), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n949), .A2(new_n742), .A3(new_n304), .A4(new_n585), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT122), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n778), .A2(new_n947), .A3(new_n948), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n261), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n943), .B(KEYINPUT121), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n261), .B1(G227), .B2(G900), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT124), .Z(new_n957));
  AND3_X1   g771(.A1(new_n945), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n945), .B2(new_n955), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(G72));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n933), .A2(new_n729), .A3(new_n938), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n962), .A2(new_n778), .A3(new_n797), .A4(new_n936), .ZN(new_n963));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  AND2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n290), .B(KEYINPUT125), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n961), .B(new_n915), .C1(new_n966), .C2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n965), .B1(new_n952), .B2(new_n924), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n272), .A2(new_n266), .ZN(new_n971));
  INV_X1    g785(.A(new_n595), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n827), .B2(new_n828), .ZN(new_n975));
  INV_X1    g789(.A(new_n965), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n971), .B2(new_n973), .ZN(new_n977));
  AOI22_X1  g791(.A1(new_n970), .A2(new_n656), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n968), .B1(new_n963), .B2(new_n965), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT126), .B1(new_n979), .B2(new_n883), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n969), .A2(new_n978), .A3(new_n980), .ZN(G57));
endmodule


