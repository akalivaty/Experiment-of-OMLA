

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U560 ( .A1(n528), .A2(n529), .ZN(n553) );
  NOR2_X1 U561 ( .A1(n722), .A2(n721), .ZN(n725) );
  NOR2_X1 U562 ( .A1(n783), .A2(n766), .ZN(n767) );
  NOR2_X1 U563 ( .A1(G651), .A2(n633), .ZN(n648) );
  NOR2_X1 U564 ( .A1(n596), .A2(n595), .ZN(n991) );
  AND2_X1 U565 ( .A1(n535), .A2(n534), .ZN(G160) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X1 U567 ( .A(KEYINPUT17), .B(n526), .Z(n574) );
  NAND2_X1 U568 ( .A1(n574), .A2(G137), .ZN(n535) );
  INV_X1 U569 ( .A(G2104), .ZN(n528) );
  NOR2_X1 U570 ( .A1(n528), .A2(G2105), .ZN(n554) );
  NAND2_X1 U571 ( .A1(G101), .A2(n554), .ZN(n527) );
  XNOR2_X1 U572 ( .A(KEYINPUT23), .B(n527), .ZN(n533) );
  INV_X1 U573 ( .A(G2105), .ZN(n529) );
  NAND2_X1 U574 ( .A1(G113), .A2(n553), .ZN(n531) );
  NOR2_X2 U575 ( .A1(G2104), .A2(n529), .ZN(n878) );
  NAND2_X1 U576 ( .A1(G125), .A2(n878), .ZN(n530) );
  NAND2_X1 U577 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U578 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  NAND2_X1 U580 ( .A1(n648), .A2(G51), .ZN(n539) );
  XNOR2_X1 U581 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n537) );
  XNOR2_X1 U582 ( .A(KEYINPUT67), .B(G651), .ZN(n541) );
  NOR2_X1 U583 ( .A1(G543), .A2(n541), .ZN(n536) );
  XNOR2_X1 U584 ( .A(n537), .B(n536), .ZN(n655) );
  NAND2_X1 U585 ( .A1(G63), .A2(n655), .ZN(n538) );
  NAND2_X1 U586 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U587 ( .A(KEYINPUT6), .B(n540), .Z(n549) );
  NOR2_X2 U588 ( .A1(n633), .A2(n541), .ZN(n651) );
  NAND2_X1 U589 ( .A1(G76), .A2(n651), .ZN(n542) );
  XNOR2_X1 U590 ( .A(KEYINPUT75), .B(n542), .ZN(n545) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n647) );
  NAND2_X1 U592 ( .A1(n647), .A2(G89), .ZN(n543) );
  XOR2_X1 U593 ( .A(n543), .B(KEYINPUT4), .Z(n544) );
  NOR2_X1 U594 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U595 ( .A(KEYINPUT5), .B(n546), .Z(n547) );
  XNOR2_X1 U596 ( .A(KEYINPUT76), .B(n547), .ZN(n548) );
  NAND2_X1 U597 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U598 ( .A(KEYINPUT7), .B(n550), .ZN(G168) );
  XOR2_X1 U599 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U600 ( .A1(n574), .A2(G138), .ZN(n552) );
  INV_X1 U601 ( .A(KEYINPUT85), .ZN(n551) );
  XNOR2_X1 U602 ( .A(n552), .B(n551), .ZN(n560) );
  AND2_X1 U603 ( .A1(n553), .A2(G114), .ZN(n558) );
  BUF_X1 U604 ( .A(n554), .Z(n875) );
  NAND2_X1 U605 ( .A1(G102), .A2(n875), .ZN(n556) );
  NAND2_X1 U606 ( .A1(G126), .A2(n878), .ZN(n555) );
  NAND2_X1 U607 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U608 ( .A1(n558), .A2(n557), .ZN(n559) );
  AND2_X1 U609 ( .A1(n560), .A2(n559), .ZN(G164) );
  NAND2_X1 U610 ( .A1(n648), .A2(G52), .ZN(n562) );
  NAND2_X1 U611 ( .A1(G64), .A2(n655), .ZN(n561) );
  NAND2_X1 U612 ( .A1(n562), .A2(n561), .ZN(n568) );
  NAND2_X1 U613 ( .A1(n647), .A2(G90), .ZN(n564) );
  NAND2_X1 U614 ( .A1(G77), .A2(n651), .ZN(n563) );
  NAND2_X1 U615 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  XNOR2_X1 U617 ( .A(KEYINPUT70), .B(n566), .ZN(n567) );
  NOR2_X1 U618 ( .A1(n568), .A2(n567), .ZN(G171) );
  AND2_X1 U619 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U620 ( .A1(G111), .A2(n553), .ZN(n570) );
  NAND2_X1 U621 ( .A1(G99), .A2(n875), .ZN(n569) );
  NAND2_X1 U622 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U623 ( .A1(n878), .A2(G123), .ZN(n571) );
  XOR2_X1 U624 ( .A(KEYINPUT18), .B(n571), .Z(n572) );
  NOR2_X1 U625 ( .A1(n573), .A2(n572), .ZN(n576) );
  BUF_X1 U626 ( .A(n574), .Z(n874) );
  NAND2_X1 U627 ( .A1(n874), .A2(G135), .ZN(n575) );
  NAND2_X1 U628 ( .A1(n576), .A2(n575), .ZN(n925) );
  XNOR2_X1 U629 ( .A(G2096), .B(n925), .ZN(n577) );
  OR2_X1 U630 ( .A1(G2100), .A2(n577), .ZN(G156) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  NAND2_X1 U632 ( .A1(n647), .A2(G88), .ZN(n579) );
  NAND2_X1 U633 ( .A1(G75), .A2(n651), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U635 ( .A1(n648), .A2(G50), .ZN(n581) );
  NAND2_X1 U636 ( .A1(G62), .A2(n655), .ZN(n580) );
  NAND2_X1 U637 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U638 ( .A1(n583), .A2(n582), .ZN(G166) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U640 ( .A(n584), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U641 ( .A(G223), .ZN(n829) );
  NAND2_X1 U642 ( .A1(n829), .A2(G567), .ZN(n585) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U644 ( .A1(G56), .A2(n655), .ZN(n586) );
  XNOR2_X1 U645 ( .A(n586), .B(KEYINPUT14), .ZN(n588) );
  NAND2_X1 U646 ( .A1(G43), .A2(n648), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n588), .A2(n587), .ZN(n596) );
  NAND2_X1 U648 ( .A1(G68), .A2(n651), .ZN(n589) );
  XNOR2_X1 U649 ( .A(KEYINPUT71), .B(n589), .ZN(n592) );
  NAND2_X1 U650 ( .A1(n647), .A2(G81), .ZN(n590) );
  XOR2_X1 U651 ( .A(n590), .B(KEYINPUT12), .Z(n591) );
  NOR2_X1 U652 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U653 ( .A(KEYINPUT13), .B(n593), .Z(n594) );
  XOR2_X1 U654 ( .A(KEYINPUT72), .B(n594), .Z(n595) );
  NAND2_X1 U655 ( .A1(n991), .A2(G860), .ZN(G153) );
  NAND2_X1 U656 ( .A1(G92), .A2(n647), .ZN(n598) );
  NAND2_X1 U657 ( .A1(G54), .A2(n648), .ZN(n597) );
  NAND2_X1 U658 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U659 ( .A1(G79), .A2(n651), .ZN(n600) );
  NAND2_X1 U660 ( .A1(G66), .A2(n655), .ZN(n599) );
  NAND2_X1 U661 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U662 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U663 ( .A(KEYINPUT15), .B(n603), .Z(n971) );
  NOR2_X1 U664 ( .A1(n971), .A2(G868), .ZN(n604) );
  XOR2_X1 U665 ( .A(KEYINPUT74), .B(n604), .Z(n607) );
  INV_X1 U666 ( .A(G868), .ZN(n620) );
  NOR2_X1 U667 ( .A1(G171), .A2(n620), .ZN(n605) );
  XNOR2_X1 U668 ( .A(KEYINPUT73), .B(n605), .ZN(n606) );
  NAND2_X1 U669 ( .A1(n607), .A2(n606), .ZN(G284) );
  NAND2_X1 U670 ( .A1(n648), .A2(G53), .ZN(n609) );
  NAND2_X1 U671 ( .A1(G65), .A2(n655), .ZN(n608) );
  NAND2_X1 U672 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U673 ( .A1(n647), .A2(G91), .ZN(n611) );
  NAND2_X1 U674 ( .A1(G78), .A2(n651), .ZN(n610) );
  NAND2_X1 U675 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U676 ( .A1(n613), .A2(n612), .ZN(n978) );
  INV_X1 U677 ( .A(n978), .ZN(G299) );
  NOR2_X1 U678 ( .A1(G286), .A2(n620), .ZN(n615) );
  NOR2_X1 U679 ( .A1(G868), .A2(G299), .ZN(n614) );
  NOR2_X1 U680 ( .A1(n615), .A2(n614), .ZN(G297) );
  INV_X1 U681 ( .A(G860), .ZN(n624) );
  NAND2_X1 U682 ( .A1(n624), .A2(G559), .ZN(n616) );
  NAND2_X1 U683 ( .A1(n616), .A2(n971), .ZN(n617) );
  XNOR2_X1 U684 ( .A(n617), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G559), .A2(n620), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n971), .A2(n618), .ZN(n619) );
  XNOR2_X1 U687 ( .A(n619), .B(KEYINPUT77), .ZN(n622) );
  AND2_X1 U688 ( .A1(n991), .A2(n620), .ZN(n621) );
  NOR2_X1 U689 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U690 ( .A1(G559), .A2(n971), .ZN(n623) );
  XNOR2_X1 U691 ( .A(n623), .B(n991), .ZN(n665) );
  NAND2_X1 U692 ( .A1(n624), .A2(n665), .ZN(n632) );
  NAND2_X1 U693 ( .A1(G93), .A2(n647), .ZN(n625) );
  XNOR2_X1 U694 ( .A(n625), .B(KEYINPUT78), .ZN(n627) );
  NAND2_X1 U695 ( .A1(G67), .A2(n655), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U697 ( .A1(n648), .A2(G55), .ZN(n629) );
  NAND2_X1 U698 ( .A1(G80), .A2(n651), .ZN(n628) );
  NAND2_X1 U699 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U700 ( .A1(n631), .A2(n630), .ZN(n667) );
  XOR2_X1 U701 ( .A(n632), .B(n667), .Z(G145) );
  NAND2_X1 U702 ( .A1(G87), .A2(n633), .ZN(n635) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U705 ( .A1(n655), .A2(n636), .ZN(n639) );
  NAND2_X1 U706 ( .A1(G49), .A2(n648), .ZN(n637) );
  XOR2_X1 U707 ( .A(KEYINPUT79), .B(n637), .Z(n638) );
  NAND2_X1 U708 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U709 ( .A1(n647), .A2(G85), .ZN(n641) );
  NAND2_X1 U710 ( .A1(G72), .A2(n651), .ZN(n640) );
  NAND2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U712 ( .A(KEYINPUT68), .B(n642), .Z(n646) );
  NAND2_X1 U713 ( .A1(n655), .A2(G60), .ZN(n644) );
  NAND2_X1 U714 ( .A1(n648), .A2(G47), .ZN(n643) );
  AND2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n646), .A2(n645), .ZN(G290) );
  NAND2_X1 U717 ( .A1(G86), .A2(n647), .ZN(n650) );
  NAND2_X1 U718 ( .A1(G48), .A2(n648), .ZN(n649) );
  NAND2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U720 ( .A1(n651), .A2(G73), .ZN(n652) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(n652), .Z(n653) );
  NOR2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U723 ( .A1(G61), .A2(n655), .ZN(n656) );
  NAND2_X1 U724 ( .A1(n657), .A2(n656), .ZN(G305) );
  XNOR2_X1 U725 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n659) );
  XNOR2_X1 U726 ( .A(G288), .B(KEYINPUT19), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U728 ( .A(G166), .B(n660), .ZN(n662) );
  XNOR2_X1 U729 ( .A(G290), .B(n978), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n667), .B(n663), .ZN(n664) );
  XNOR2_X1 U732 ( .A(n664), .B(G305), .ZN(n900) );
  XNOR2_X1 U733 ( .A(n900), .B(n665), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n666), .A2(G868), .ZN(n669) );
  OR2_X1 U735 ( .A1(G868), .A2(n667), .ZN(n668) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U739 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U740 ( .A(n672), .B(KEYINPUT82), .ZN(n673) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U742 ( .A1(G2072), .A2(n674), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U744 ( .A1(G69), .A2(G120), .ZN(n675) );
  NOR2_X1 U745 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U746 ( .A1(G108), .A2(n676), .ZN(n833) );
  NAND2_X1 U747 ( .A1(n833), .A2(G567), .ZN(n683) );
  XOR2_X1 U748 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n678) );
  NAND2_X1 U749 ( .A1(G132), .A2(G82), .ZN(n677) );
  XNOR2_X1 U750 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X1 U751 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U752 ( .A1(G96), .A2(n680), .ZN(n681) );
  XNOR2_X1 U753 ( .A(KEYINPUT84), .B(n681), .ZN(n834) );
  NAND2_X1 U754 ( .A1(G2106), .A2(n834), .ZN(n682) );
  NAND2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n835) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U757 ( .A1(n835), .A2(n684), .ZN(n832) );
  NAND2_X1 U758 ( .A1(n832), .A2(G36), .ZN(G176) );
  INV_X1 U759 ( .A(G166), .ZN(G303) );
  NAND2_X1 U760 ( .A1(G140), .A2(n874), .ZN(n686) );
  NAND2_X1 U761 ( .A1(G104), .A2(n875), .ZN(n685) );
  NAND2_X1 U762 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U763 ( .A(KEYINPUT34), .B(n687), .ZN(n692) );
  NAND2_X1 U764 ( .A1(G116), .A2(n553), .ZN(n689) );
  NAND2_X1 U765 ( .A1(G128), .A2(n878), .ZN(n688) );
  NAND2_X1 U766 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U767 ( .A(n690), .B(KEYINPUT35), .Z(n691) );
  NOR2_X1 U768 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U769 ( .A(KEYINPUT36), .B(n693), .Z(n694) );
  XOR2_X1 U770 ( .A(KEYINPUT88), .B(n694), .Z(n895) );
  XOR2_X1 U771 ( .A(G2067), .B(KEYINPUT37), .Z(n695) );
  XNOR2_X1 U772 ( .A(KEYINPUT87), .B(n695), .ZN(n820) );
  NOR2_X1 U773 ( .A1(n895), .A2(n820), .ZN(n928) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n698) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n700) );
  NOR2_X1 U776 ( .A1(n698), .A2(n700), .ZN(n697) );
  XNOR2_X1 U777 ( .A(n697), .B(KEYINPUT86), .ZN(n822) );
  NAND2_X1 U778 ( .A1(n928), .A2(n822), .ZN(n818) );
  INV_X1 U779 ( .A(n818), .ZN(n787) );
  INV_X1 U780 ( .A(KEYINPUT94), .ZN(n699) );
  XNOR2_X1 U781 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U782 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X2 U783 ( .A(n702), .B(KEYINPUT64), .ZN(n719) );
  NAND2_X1 U784 ( .A1(n719), .A2(G8), .ZN(n783) );
  INV_X1 U785 ( .A(n719), .ZN(n731) );
  NAND2_X1 U786 ( .A1(n731), .A2(G2067), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n719), .A2(G1348), .ZN(n703) );
  NAND2_X1 U788 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U789 ( .A(n705), .B(KEYINPUT98), .Z(n706) );
  OR2_X1 U790 ( .A1(n971), .A2(n706), .ZN(n717) );
  NAND2_X1 U791 ( .A1(n706), .A2(n971), .ZN(n715) );
  INV_X1 U792 ( .A(G1996), .ZN(n707) );
  NOR2_X1 U793 ( .A1(n719), .A2(n707), .ZN(n709) );
  XOR2_X1 U794 ( .A(KEYINPUT66), .B(KEYINPUT26), .Z(n708) );
  XNOR2_X1 U795 ( .A(n709), .B(n708), .ZN(n711) );
  INV_X1 U796 ( .A(n731), .ZN(n746) );
  NAND2_X1 U797 ( .A1(n746), .A2(G1341), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U799 ( .A(n712), .B(KEYINPUT97), .ZN(n713) );
  NAND2_X1 U800 ( .A1(n713), .A2(n991), .ZN(n714) );
  NAND2_X1 U801 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U802 ( .A1(n717), .A2(n716), .ZN(n724) );
  NAND2_X1 U803 ( .A1(G2072), .A2(n731), .ZN(n718) );
  XNOR2_X1 U804 ( .A(n718), .B(KEYINPUT27), .ZN(n722) );
  NAND2_X1 U805 ( .A1(n719), .A2(G1956), .ZN(n720) );
  XOR2_X1 U806 ( .A(KEYINPUT96), .B(n720), .Z(n721) );
  NAND2_X1 U807 ( .A1(n725), .A2(n978), .ZN(n723) );
  NAND2_X1 U808 ( .A1(n724), .A2(n723), .ZN(n728) );
  NOR2_X1 U809 ( .A1(n725), .A2(n978), .ZN(n726) );
  XOR2_X1 U810 ( .A(n726), .B(KEYINPUT28), .Z(n727) );
  NAND2_X1 U811 ( .A1(n728), .A2(n727), .ZN(n730) );
  XNOR2_X1 U812 ( .A(KEYINPUT29), .B(KEYINPUT99), .ZN(n729) );
  XNOR2_X1 U813 ( .A(n730), .B(n729), .ZN(n735) );
  XNOR2_X1 U814 ( .A(KEYINPUT25), .B(G2078), .ZN(n950) );
  NAND2_X1 U815 ( .A1(n731), .A2(n950), .ZN(n733) );
  INV_X1 U816 ( .A(G1961), .ZN(n1011) );
  NAND2_X1 U817 ( .A1(n746), .A2(n1011), .ZN(n732) );
  NAND2_X1 U818 ( .A1(n733), .A2(n732), .ZN(n740) );
  NAND2_X1 U819 ( .A1(n740), .A2(G171), .ZN(n734) );
  NAND2_X1 U820 ( .A1(n735), .A2(n734), .ZN(n745) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n783), .ZN(n757) );
  NOR2_X1 U822 ( .A1(n719), .A2(G2084), .ZN(n754) );
  INV_X1 U823 ( .A(n754), .ZN(n736) );
  NAND2_X1 U824 ( .A1(G8), .A2(n736), .ZN(n737) );
  OR2_X1 U825 ( .A1(n757), .A2(n737), .ZN(n738) );
  XNOR2_X1 U826 ( .A(KEYINPUT30), .B(n738), .ZN(n739) );
  NOR2_X1 U827 ( .A1(G168), .A2(n739), .ZN(n742) );
  NOR2_X1 U828 ( .A1(G171), .A2(n740), .ZN(n741) );
  NOR2_X1 U829 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U830 ( .A(KEYINPUT31), .B(n743), .Z(n744) );
  NAND2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n755) );
  NAND2_X1 U832 ( .A1(n755), .A2(G286), .ZN(n751) );
  NOR2_X1 U833 ( .A1(n746), .A2(G2090), .ZN(n748) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n783), .ZN(n747) );
  NOR2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n749), .A2(G303), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n752), .A2(G8), .ZN(n753) );
  XNOR2_X1 U839 ( .A(n753), .B(KEYINPUT32), .ZN(n761) );
  NAND2_X1 U840 ( .A1(G8), .A2(n754), .ZN(n759) );
  INV_X1 U841 ( .A(n755), .ZN(n756) );
  NOR2_X1 U842 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U843 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U844 ( .A1(n761), .A2(n760), .ZN(n776) );
  NOR2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NOR2_X1 U846 ( .A1(G1971), .A2(G303), .ZN(n762) );
  NOR2_X1 U847 ( .A1(n974), .A2(n762), .ZN(n763) );
  NAND2_X1 U848 ( .A1(n776), .A2(n763), .ZN(n765) );
  NAND2_X1 U849 ( .A1(G288), .A2(G1976), .ZN(n764) );
  XNOR2_X1 U850 ( .A(n764), .B(KEYINPUT100), .ZN(n975) );
  NAND2_X1 U851 ( .A1(n765), .A2(n975), .ZN(n766) );
  XNOR2_X1 U852 ( .A(KEYINPUT65), .B(n767), .ZN(n768) );
  INV_X1 U853 ( .A(n768), .ZN(n769) );
  NOR2_X1 U854 ( .A1(KEYINPUT33), .A2(n769), .ZN(n772) );
  NAND2_X1 U855 ( .A1(n974), .A2(KEYINPUT33), .ZN(n770) );
  NOR2_X1 U856 ( .A1(n770), .A2(n783), .ZN(n771) );
  NOR2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U858 ( .A(G1981), .B(G305), .Z(n987) );
  NAND2_X1 U859 ( .A1(n773), .A2(n987), .ZN(n779) );
  NOR2_X1 U860 ( .A1(G2090), .A2(G303), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G8), .A2(n774), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n777), .A2(n783), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n785) );
  NOR2_X1 U865 ( .A1(G1981), .A2(G305), .ZN(n780) );
  XNOR2_X1 U866 ( .A(n780), .B(KEYINPUT95), .ZN(n781) );
  XNOR2_X1 U867 ( .A(KEYINPUT24), .B(n781), .ZN(n782) );
  NOR2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U869 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U870 ( .A1(n787), .A2(n786), .ZN(n810) );
  NAND2_X1 U871 ( .A1(G107), .A2(n553), .ZN(n789) );
  NAND2_X1 U872 ( .A1(G119), .A2(n878), .ZN(n788) );
  NAND2_X1 U873 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U874 ( .A(KEYINPUT89), .B(n790), .ZN(n794) );
  NAND2_X1 U875 ( .A1(G131), .A2(n874), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G95), .A2(n875), .ZN(n791) );
  AND2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n794), .A2(n793), .ZN(n891) );
  NAND2_X1 U879 ( .A1(G1991), .A2(n891), .ZN(n795) );
  XOR2_X1 U880 ( .A(KEYINPUT90), .B(n795), .Z(n807) );
  NAND2_X1 U881 ( .A1(G141), .A2(n874), .ZN(n805) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(KEYINPUT92), .Z(n797) );
  NAND2_X1 U883 ( .A1(G105), .A2(n875), .ZN(n796) );
  XNOR2_X1 U884 ( .A(n797), .B(n796), .ZN(n802) );
  NAND2_X1 U885 ( .A1(G117), .A2(n553), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G129), .A2(n878), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U888 ( .A(KEYINPUT91), .B(n800), .Z(n801) );
  NOR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U890 ( .A(KEYINPUT93), .B(n803), .Z(n804) );
  NAND2_X1 U891 ( .A1(n805), .A2(n804), .ZN(n892) );
  AND2_X1 U892 ( .A1(n892), .A2(G1996), .ZN(n806) );
  NOR2_X1 U893 ( .A1(n807), .A2(n806), .ZN(n811) );
  XOR2_X1 U894 ( .A(G1986), .B(G290), .Z(n972) );
  NAND2_X1 U895 ( .A1(n811), .A2(n972), .ZN(n808) );
  NAND2_X1 U896 ( .A1(n808), .A2(n822), .ZN(n809) );
  NAND2_X1 U897 ( .A1(n810), .A2(n809), .ZN(n825) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n892), .ZN(n931) );
  INV_X1 U899 ( .A(n811), .ZN(n937) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n891), .ZN(n924) );
  NOR2_X1 U902 ( .A1(n812), .A2(n924), .ZN(n813) );
  NOR2_X1 U903 ( .A1(n937), .A2(n813), .ZN(n814) );
  NOR2_X1 U904 ( .A1(n931), .A2(n814), .ZN(n817) );
  XOR2_X1 U905 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n815) );
  XNOR2_X1 U906 ( .A(KEYINPUT39), .B(n815), .ZN(n816) );
  XNOR2_X1 U907 ( .A(n817), .B(n816), .ZN(n819) );
  NAND2_X1 U908 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U909 ( .A1(n895), .A2(n820), .ZN(n941) );
  NAND2_X1 U910 ( .A1(n821), .A2(n941), .ZN(n823) );
  NAND2_X1 U911 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U912 ( .A1(n825), .A2(n824), .ZN(n828) );
  XOR2_X1 U913 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n826) );
  XNOR2_X1 U914 ( .A(KEYINPUT40), .B(n826), .ZN(n827) );
  XNOR2_X1 U915 ( .A(n828), .B(n827), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U918 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U920 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U922 ( .A(G132), .ZN(G219) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G82), .ZN(G220) );
  INV_X1 U926 ( .A(G69), .ZN(G235) );
  NOR2_X1 U927 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  INV_X1 U929 ( .A(n835), .ZN(G319) );
  XOR2_X1 U930 ( .A(KEYINPUT105), .B(G2090), .Z(n837) );
  XNOR2_X1 U931 ( .A(G2072), .B(G2084), .ZN(n836) );
  XNOR2_X1 U932 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U933 ( .A(n838), .B(G2096), .Z(n840) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2078), .ZN(n839) );
  XNOR2_X1 U935 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U936 ( .A(KEYINPUT43), .B(G2678), .Z(n842) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(G2100), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U939 ( .A(n844), .B(n843), .Z(G227) );
  XOR2_X1 U940 ( .A(G1981), .B(G1961), .Z(n846) );
  XNOR2_X1 U941 ( .A(G1966), .B(G1956), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U943 ( .A(n847), .B(G2474), .Z(n849) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G1976), .Z(n851) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1971), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G124), .A2(n878), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n854), .B(KEYINPUT106), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U953 ( .A1(G112), .A2(n553), .ZN(n856) );
  NAND2_X1 U954 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U955 ( .A1(G136), .A2(n874), .ZN(n859) );
  NAND2_X1 U956 ( .A1(G100), .A2(n875), .ZN(n858) );
  NAND2_X1 U957 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U958 ( .A1(n861), .A2(n860), .ZN(G162) );
  XNOR2_X1 U959 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n925), .B(KEYINPUT48), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n887) );
  NAND2_X1 U962 ( .A1(n875), .A2(G106), .ZN(n864) );
  XOR2_X1 U963 ( .A(KEYINPUT109), .B(n864), .Z(n866) );
  NAND2_X1 U964 ( .A1(n874), .A2(G142), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n867), .B(KEYINPUT45), .ZN(n873) );
  NAND2_X1 U967 ( .A1(n553), .A2(G118), .ZN(n868) );
  XOR2_X1 U968 ( .A(KEYINPUT107), .B(n868), .Z(n870) );
  NAND2_X1 U969 ( .A1(n878), .A2(G130), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U971 ( .A(KEYINPUT108), .B(n871), .Z(n872) );
  NAND2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n885) );
  NAND2_X1 U973 ( .A1(G139), .A2(n874), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G103), .A2(n875), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n883) );
  NAND2_X1 U976 ( .A1(G115), .A2(n553), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G127), .A2(n878), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U980 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U981 ( .A(KEYINPUT110), .B(n884), .Z(n919) );
  XNOR2_X1 U982 ( .A(n885), .B(n919), .ZN(n886) );
  XOR2_X1 U983 ( .A(n887), .B(n886), .Z(n889) );
  XNOR2_X1 U984 ( .A(G160), .B(G162), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n894) );
  XOR2_X1 U987 ( .A(G164), .B(n892), .Z(n893) );
  XNOR2_X1 U988 ( .A(n894), .B(n893), .ZN(n896) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U990 ( .A1(G37), .A2(n897), .ZN(G395) );
  XOR2_X1 U991 ( .A(G286), .B(G171), .Z(n899) );
  XNOR2_X1 U992 ( .A(n991), .B(n971), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U995 ( .A1(G37), .A2(n902), .ZN(n903) );
  XNOR2_X1 U996 ( .A(KEYINPUT112), .B(n903), .ZN(G397) );
  XOR2_X1 U997 ( .A(G2451), .B(G2430), .Z(n905) );
  XNOR2_X1 U998 ( .A(G2438), .B(G2443), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n911) );
  XOR2_X1 U1000 ( .A(G2435), .B(G2454), .Z(n907) );
  XNOR2_X1 U1001 ( .A(G1348), .B(G1341), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1003 ( .A(G2446), .B(G2427), .Z(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1005 ( .A(n911), .B(n910), .Z(n912) );
  NAND2_X1 U1006 ( .A1(G14), .A2(n912), .ZN(n918) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G171), .ZN(G301) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  INV_X1 U1016 ( .A(n918), .ZN(G401) );
  INV_X1 U1017 ( .A(KEYINPUT55), .ZN(n967) );
  XOR2_X1 U1018 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n944) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n921) );
  XNOR2_X1 U1020 ( .A(G2072), .B(n919), .ZN(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1022 ( .A(KEYINPUT50), .B(n922), .Z(n940) );
  XOR2_X1 U1023 ( .A(G160), .B(G2084), .Z(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1027 ( .A(KEYINPUT113), .B(n929), .Z(n935) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1030 ( .A(KEYINPUT51), .B(n932), .Z(n933) );
  XNOR2_X1 U1031 ( .A(KEYINPUT114), .B(n933), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(KEYINPUT115), .B(n938), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(n944), .B(n943), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n967), .A2(n945), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n946), .A2(G29), .ZN(n1031) );
  XNOR2_X1 U1040 ( .A(KEYINPUT117), .B(G2090), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(n947), .B(G35), .ZN(n965) );
  XNOR2_X1 U1042 ( .A(G2084), .B(G34), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(n948), .B(KEYINPUT54), .ZN(n963) );
  XOR2_X1 U1044 ( .A(G1991), .B(G25), .Z(n949) );
  NAND2_X1 U1045 ( .A1(n949), .A2(G28), .ZN(n960) );
  XNOR2_X1 U1046 ( .A(G27), .B(n950), .ZN(n958) );
  XNOR2_X1 U1047 ( .A(G1996), .B(G32), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(G2072), .B(G33), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(n951), .B(KEYINPUT118), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(G26), .B(G2067), .ZN(n952) );
  NOR2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(KEYINPUT119), .B(n954), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(n961), .B(KEYINPUT53), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(n967), .B(n966), .ZN(n969) );
  INV_X1 U1060 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n970), .ZN(n1029) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n997) );
  XNOR2_X1 U1064 ( .A(n971), .B(G1348), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n986) );
  INV_X1 U1066 ( .A(n974), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(n977), .B(KEYINPUT121), .ZN(n984) );
  XNOR2_X1 U1069 ( .A(G166), .B(G1971), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n978), .B(G1956), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(G1961), .B(G301), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n995) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(n989), .B(KEYINPUT120), .ZN(n990) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n990), .Z(n993) );
  XOR2_X1 U1080 ( .A(n991), .B(G1341), .Z(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n1027) );
  INV_X1 U1084 ( .A(G16), .ZN(n1025) );
  XOR2_X1 U1085 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n1007) );
  XNOR2_X1 U1086 ( .A(G1956), .B(G20), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G19), .B(G1341), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1005) );
  XOR2_X1 U1089 ( .A(KEYINPUT122), .B(G4), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(G1348), .B(KEYINPUT59), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(n1001), .B(n1000), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G1981), .B(G6), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(n1007), .B(n1006), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G21), .B(G1966), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT124), .B(n1010), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(n1011), .B(G5), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1022) );
  XOR2_X1 U1101 ( .A(G1971), .B(G22), .Z(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT125), .B(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(G23), .B(G1976), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1105 ( .A(KEYINPUT126), .B(n1017), .Z(n1019) );
  XNOR2_X1 U1106 ( .A(G1986), .B(G24), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1020), .Z(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1032), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

