

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760;

  XNOR2_X1 U366 ( .A(n374), .B(n449), .ZN(n473) );
  XNOR2_X1 U367 ( .A(n385), .B(G119), .ZN(n374) );
  INV_X1 U368 ( .A(n550), .ZN(n655) );
  NOR2_X2 U369 ( .A1(n411), .A2(n710), .ZN(n715) );
  NOR2_X2 U370 ( .A1(n600), .A2(n574), .ZN(n575) );
  XNOR2_X2 U371 ( .A(n581), .B(KEYINPUT33), .ZN(n688) );
  XNOR2_X2 U372 ( .A(n571), .B(KEYINPUT0), .ZN(n600) );
  XNOR2_X2 U373 ( .A(n435), .B(n434), .ZN(n455) );
  XNOR2_X2 U374 ( .A(KEYINPUT81), .B(G143), .ZN(n435) );
  XNOR2_X2 U375 ( .A(n455), .B(G134), .ZN(n477) );
  XOR2_X1 U376 ( .A(KEYINPUT41), .B(n469), .Z(n696) );
  NOR2_X1 U377 ( .A1(n657), .A2(n655), .ZN(n684) );
  NOR2_X2 U378 ( .A1(n759), .A2(n757), .ZN(n388) );
  INV_X1 U379 ( .A(n566), .ZN(n344) );
  XNOR2_X1 U380 ( .A(n465), .B(n464), .ZN(n535) );
  NOR2_X2 U381 ( .A1(G953), .A2(G237), .ZN(n470) );
  INV_X1 U382 ( .A(G128), .ZN(n434) );
  NOR2_X1 U383 ( .A1(n629), .A2(n727), .ZN(n630) );
  INV_X1 U384 ( .A(n717), .ZN(n723) );
  XNOR2_X1 U385 ( .A(n596), .B(n576), .ZN(n578) );
  BUF_X1 U386 ( .A(n535), .Z(n466) );
  XNOR2_X1 U387 ( .A(n548), .B(KEYINPUT6), .ZN(n594) );
  XNOR2_X1 U388 ( .A(n480), .B(n636), .ZN(n548) );
  XNOR2_X1 U389 ( .A(n422), .B(n498), .ZN(n724) );
  XNOR2_X1 U390 ( .A(n459), .B(G146), .ZN(n743) );
  XNOR2_X1 U391 ( .A(G113), .B(KEYINPUT71), .ZN(n449) );
  XNOR2_X1 U392 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n459) );
  XNOR2_X2 U393 ( .A(n345), .B(G469), .ZN(n554) );
  NOR2_X1 U394 ( .A1(n713), .A2(G902), .ZN(n345) );
  NAND2_X1 U395 ( .A1(n578), .A2(n577), .ZN(n634) );
  NOR2_X2 U396 ( .A1(n682), .A2(n683), .ZN(n469) );
  XNOR2_X2 U397 ( .A(n510), .B(n509), .ZN(n746) );
  XNOR2_X1 U398 ( .A(n384), .B(KEYINPUT68), .ZN(n476) );
  INV_X1 U399 ( .A(G131), .ZN(n384) );
  XNOR2_X1 U400 ( .A(n379), .B(n442), .ZN(n718) );
  XNOR2_X1 U401 ( .A(n448), .B(n349), .ZN(n379) );
  NAND2_X1 U402 ( .A1(n556), .A2(KEYINPUT47), .ZN(n540) );
  AND2_X1 U403 ( .A1(n391), .A2(n390), .ZN(n389) );
  NOR2_X1 U404 ( .A1(n425), .A2(n392), .ZN(n391) );
  NOR2_X1 U405 ( .A1(n651), .A2(n546), .ZN(n547) );
  AND2_X1 U406 ( .A1(n634), .A2(n635), .ZN(n593) );
  XNOR2_X1 U407 ( .A(n472), .B(G137), .ZN(n373) );
  XNOR2_X1 U408 ( .A(n444), .B(n443), .ZN(n744) );
  INV_X1 U409 ( .A(G140), .ZN(n443) );
  XNOR2_X1 U410 ( .A(KEYINPUT10), .B(G125), .ZN(n444) );
  XNOR2_X1 U411 ( .A(KEYINPUT67), .B(G101), .ZN(n460) );
  INV_X1 U412 ( .A(n519), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n744), .B(G146), .ZN(n497) );
  XNOR2_X1 U414 ( .A(G110), .B(KEYINPUT92), .ZN(n492) );
  NAND2_X1 U415 ( .A1(n403), .A2(n413), .ZN(n412) );
  NOR2_X1 U416 ( .A1(n414), .A2(n727), .ZN(n413) );
  NOR2_X1 U417 ( .A1(n419), .A2(G475), .ZN(n414) );
  NAND2_X1 U418 ( .A1(G234), .A2(G237), .ZN(n486) );
  AND2_X1 U419 ( .A1(n371), .A2(n368), .ZN(n367) );
  INV_X1 U420 ( .A(n583), .ZN(n369) );
  NAND2_X1 U421 ( .A1(n366), .A2(KEYINPUT34), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n421), .B(n505), .ZN(n663) );
  NOR2_X1 U423 ( .A1(n724), .A2(G902), .ZN(n421) );
  AND2_X1 U424 ( .A1(n406), .A2(KEYINPUT60), .ZN(n405) );
  XNOR2_X1 U425 ( .A(n540), .B(n539), .ZN(n545) );
  INV_X1 U426 ( .A(KEYINPUT86), .ZN(n612) );
  INV_X1 U427 ( .A(G237), .ZN(n463) );
  XNOR2_X1 U428 ( .A(G902), .B(KEYINPUT15), .ZN(n618) );
  XNOR2_X1 U429 ( .A(G113), .B(G143), .ZN(n445) );
  XNOR2_X1 U430 ( .A(G119), .B(G128), .ZN(n490) );
  NOR2_X1 U431 ( .A1(n719), .A2(n416), .ZN(n415) );
  INV_X1 U432 ( .A(G475), .ZN(n416) );
  XNOR2_X1 U433 ( .A(KEYINPUT18), .B(G125), .ZN(n453) );
  AND2_X1 U434 ( .A1(n398), .A2(n397), .ZN(n396) );
  NAND2_X1 U435 ( .A1(n394), .A2(n356), .ZN(n397) );
  INV_X1 U436 ( .A(KEYINPUT48), .ZN(n361) );
  NOR2_X1 U437 ( .A1(n605), .A2(n582), .ZN(n370) );
  INV_X1 U438 ( .A(G902), .ZN(n479) );
  XNOR2_X1 U439 ( .A(n473), .B(n372), .ZN(n474) );
  XNOR2_X1 U440 ( .A(n373), .B(n471), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n734) );
  XNOR2_X1 U442 ( .A(G107), .B(G104), .ZN(n377) );
  XNOR2_X1 U443 ( .A(KEYINPUT89), .B(G110), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n473), .B(n450), .ZN(n736) );
  XNOR2_X1 U445 ( .A(G107), .B(KEYINPUT99), .ZN(n426) );
  XOR2_X1 U446 ( .A(KEYINPUT7), .B(KEYINPUT100), .Z(n427) );
  AND2_X1 U447 ( .A1(n364), .A2(n594), .ZN(n580) );
  INV_X1 U448 ( .A(n598), .ZN(n364) );
  NOR2_X1 U449 ( .A1(n380), .A2(n550), .ZN(n561) );
  NAND2_X1 U450 ( .A1(n594), .A2(n381), .ZN(n380) );
  NOR2_X1 U451 ( .A1(n549), .A2(n382), .ZN(n381) );
  INV_X1 U452 ( .A(n679), .ZN(n382) );
  NOR2_X1 U453 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U454 ( .A1(n518), .A2(n354), .ZN(n524) );
  BUF_X1 U455 ( .A(n548), .Z(n667) );
  XNOR2_X1 U456 ( .A(n378), .B(n348), .ZN(n542) );
  OR2_X1 U457 ( .A1(n718), .A2(G902), .ZN(n378) );
  XNOR2_X1 U458 ( .A(n499), .B(n352), .ZN(n422) );
  XNOR2_X1 U459 ( .A(KEYINPUT91), .B(G140), .ZN(n512) );
  XNOR2_X1 U460 ( .A(n532), .B(n531), .ZN(n759) );
  AND2_X1 U461 ( .A1(n375), .A2(n655), .ZN(n532) );
  XNOR2_X1 U462 ( .A(n586), .B(n585), .ZN(n635) );
  AND2_X1 U463 ( .A1(n363), .A2(n418), .ZN(G63) );
  AND2_X1 U464 ( .A1(n410), .A2(n409), .ZN(n408) );
  AND2_X1 U465 ( .A1(n399), .A2(n357), .ZN(n346) );
  XOR2_X1 U466 ( .A(n554), .B(KEYINPUT108), .Z(n347) );
  XOR2_X1 U467 ( .A(KEYINPUT13), .B(G475), .Z(n348) );
  XOR2_X1 U468 ( .A(n441), .B(n440), .Z(n349) );
  AND2_X1 U469 ( .A1(n605), .A2(n582), .ZN(n350) );
  AND2_X1 U470 ( .A1(n347), .A2(n344), .ZN(n351) );
  AND2_X1 U471 ( .A1(n500), .A2(G221), .ZN(n352) );
  AND2_X1 U472 ( .A1(n591), .A2(n590), .ZN(n353) );
  INV_X1 U473 ( .A(n594), .ZN(n590) );
  AND2_X1 U474 ( .A1(n587), .A2(n360), .ZN(n354) );
  AND2_X1 U475 ( .A1(n565), .A2(n402), .ZN(n355) );
  INV_X1 U476 ( .A(KEYINPUT34), .ZN(n582) );
  AND2_X1 U477 ( .A1(n393), .A2(KEYINPUT65), .ZN(n356) );
  AND2_X1 U478 ( .A1(n402), .A2(n619), .ZN(n357) );
  AND2_X1 U479 ( .A1(KEYINPUT65), .A2(n401), .ZN(n358) );
  AND2_X1 U480 ( .A1(n719), .A2(n417), .ZN(n359) );
  AND2_X1 U481 ( .A1(n628), .A2(G953), .ZN(n727) );
  INV_X1 U482 ( .A(n727), .ZN(n418) );
  INV_X1 U483 ( .A(KEYINPUT60), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n362), .B(n361), .ZN(n383) );
  NAND2_X1 U485 ( .A1(n387), .A2(n389), .ZN(n362) );
  XNOR2_X1 U486 ( .A(n721), .B(n722), .ZN(n363) );
  NAND2_X1 U487 ( .A1(n367), .A2(n365), .ZN(n586) );
  INV_X1 U488 ( .A(n688), .ZN(n366) );
  NOR2_X1 U489 ( .A1(n370), .A2(n369), .ZN(n368) );
  NAND2_X1 U490 ( .A1(n688), .A2(n350), .ZN(n371) );
  NAND2_X1 U491 ( .A1(n375), .A2(n657), .ZN(n560) );
  XNOR2_X1 U492 ( .A(n528), .B(n527), .ZN(n375) );
  NAND2_X1 U493 ( .A1(n561), .A2(n466), .ZN(n552) );
  NAND2_X1 U494 ( .A1(n383), .A2(n565), .ZN(n701) );
  NAND2_X1 U495 ( .A1(n383), .A2(n355), .ZN(n394) );
  XNOR2_X2 U496 ( .A(G116), .B(KEYINPUT3), .ZN(n385) );
  NOR2_X1 U497 ( .A1(n702), .A2(n701), .ZN(n620) );
  NAND2_X1 U498 ( .A1(n702), .A2(n358), .ZN(n398) );
  NAND2_X1 U499 ( .A1(n702), .A2(n401), .ZN(n400) );
  XNOR2_X2 U500 ( .A(n617), .B(n616), .ZN(n702) );
  NAND2_X1 U501 ( .A1(n386), .A2(n668), .ZN(n596) );
  NAND2_X1 U502 ( .A1(n353), .A2(n386), .ZN(n592) );
  XNOR2_X1 U503 ( .A(n575), .B(KEYINPUT22), .ZN(n386) );
  NAND2_X1 U504 ( .A1(n344), .A2(n424), .ZN(n571) );
  XNOR2_X1 U505 ( .A(n547), .B(KEYINPUT82), .ZN(n390) );
  XNOR2_X1 U506 ( .A(n516), .B(n517), .ZN(n757) );
  XNOR2_X1 U507 ( .A(n388), .B(KEYINPUT46), .ZN(n387) );
  INV_X1 U508 ( .A(n662), .ZN(n392) );
  NAND2_X1 U509 ( .A1(n701), .A2(n401), .ZN(n399) );
  NAND2_X1 U510 ( .A1(n402), .A2(KEYINPUT2), .ZN(n393) );
  NAND2_X1 U511 ( .A1(n396), .A2(n395), .ZN(n622) );
  NAND2_X1 U512 ( .A1(n346), .A2(n400), .ZN(n395) );
  INV_X1 U513 ( .A(KEYINPUT2), .ZN(n401) );
  INV_X1 U514 ( .A(n618), .ZN(n402) );
  NAND2_X1 U515 ( .A1(n723), .A2(n415), .ZN(n403) );
  NAND2_X1 U516 ( .A1(n408), .A2(n404), .ZN(G60) );
  NAND2_X1 U517 ( .A1(n407), .A2(n405), .ZN(n404) );
  NAND2_X1 U518 ( .A1(n411), .A2(n719), .ZN(n406) );
  INV_X1 U519 ( .A(n412), .ZN(n407) );
  NAND2_X1 U520 ( .A1(n411), .A2(n359), .ZN(n409) );
  NAND2_X1 U521 ( .A1(n412), .A2(n417), .ZN(n410) );
  INV_X1 U522 ( .A(n723), .ZN(n411) );
  INV_X1 U523 ( .A(n719), .ZN(n419) );
  NAND2_X1 U524 ( .A1(n420), .A2(n351), .ZN(n556) );
  XNOR2_X1 U525 ( .A(n507), .B(KEYINPUT28), .ZN(n420) );
  AND2_X1 U526 ( .A1(n420), .A2(n347), .ZN(n538) );
  OR2_X1 U527 ( .A1(n614), .A2(KEYINPUT44), .ZN(n423) );
  AND2_X1 U528 ( .A1(n570), .A2(n569), .ZN(n424) );
  XOR2_X1 U529 ( .A(KEYINPUT74), .B(n558), .Z(n425) );
  INV_X1 U530 ( .A(KEYINPUT83), .ZN(n539) );
  INV_X1 U531 ( .A(KEYINPUT65), .ZN(n619) );
  NOR2_X1 U532 ( .A1(n667), .A2(n549), .ZN(n507) );
  XNOR2_X1 U533 ( .A(n520), .B(KEYINPUT107), .ZN(n521) );
  XNOR2_X1 U534 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U535 ( .A(n530), .B(KEYINPUT40), .ZN(n531) );
  XOR2_X1 U536 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n517) );
  XNOR2_X1 U537 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U538 ( .A(n428), .B(KEYINPUT9), .Z(n430) );
  XNOR2_X1 U539 ( .A(G116), .B(G122), .ZN(n429) );
  XNOR2_X1 U540 ( .A(n430), .B(n429), .ZN(n433) );
  INV_X4 U541 ( .A(G953), .ZN(n750) );
  NAND2_X1 U542 ( .A1(G234), .A2(n750), .ZN(n431) );
  XOR2_X1 U543 ( .A(KEYINPUT8), .B(n431), .Z(n500) );
  NAND2_X1 U544 ( .A1(G217), .A2(n500), .ZN(n432) );
  XNOR2_X1 U545 ( .A(n433), .B(n432), .ZN(n436) );
  XNOR2_X1 U546 ( .A(n436), .B(n477), .ZN(n722) );
  NAND2_X1 U547 ( .A1(n722), .A2(n479), .ZN(n437) );
  XNOR2_X1 U548 ( .A(n437), .B(G478), .ZN(n541) );
  XOR2_X1 U549 ( .A(n476), .B(KEYINPUT97), .Z(n439) );
  NAND2_X1 U550 ( .A1(G214), .A2(n470), .ZN(n438) );
  XNOR2_X1 U551 ( .A(n439), .B(n438), .ZN(n442) );
  XOR2_X1 U552 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n441) );
  XNOR2_X1 U553 ( .A(KEYINPUT98), .B(KEYINPUT96), .ZN(n440) );
  XOR2_X1 U554 ( .A(G104), .B(G122), .Z(n446) );
  XNOR2_X1 U555 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U556 ( .A(n497), .B(n447), .ZN(n448) );
  OR2_X1 U557 ( .A1(n541), .A2(n542), .ZN(n682) );
  XNOR2_X1 U558 ( .A(KEYINPUT16), .B(G122), .ZN(n450) );
  XOR2_X1 U559 ( .A(KEYINPUT17), .B(KEYINPUT79), .Z(n452) );
  NAND2_X1 U560 ( .A1(G224), .A2(n750), .ZN(n451) );
  XNOR2_X1 U561 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U562 ( .A(n454), .B(n453), .ZN(n457) );
  INV_X1 U563 ( .A(n455), .ZN(n456) );
  XNOR2_X1 U564 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U565 ( .A(n736), .B(n458), .ZN(n462) );
  XNOR2_X1 U566 ( .A(n743), .B(n460), .ZN(n475) );
  XNOR2_X1 U567 ( .A(n734), .B(KEYINPUT73), .ZN(n461) );
  XNOR2_X1 U568 ( .A(n475), .B(n461), .ZN(n514) );
  XNOR2_X1 U569 ( .A(n462), .B(n514), .ZN(n623) );
  NAND2_X1 U570 ( .A1(n623), .A2(n618), .ZN(n465) );
  NAND2_X1 U571 ( .A1(n479), .A2(n463), .ZN(n468) );
  AND2_X1 U572 ( .A1(n468), .A2(G210), .ZN(n464) );
  XNOR2_X1 U573 ( .A(KEYINPUT38), .B(KEYINPUT76), .ZN(n467) );
  XNOR2_X1 U574 ( .A(n466), .B(n467), .ZN(n526) );
  INV_X1 U575 ( .A(n526), .ZN(n680) );
  NAND2_X1 U576 ( .A1(n468), .A2(G214), .ZN(n679) );
  NAND2_X1 U577 ( .A1(n680), .A2(n679), .ZN(n683) );
  NAND2_X1 U578 ( .A1(n470), .A2(G210), .ZN(n472) );
  XOR2_X1 U579 ( .A(KEYINPUT5), .B(KEYINPUT95), .Z(n471) );
  XNOR2_X1 U580 ( .A(n475), .B(n474), .ZN(n478) );
  XNOR2_X2 U581 ( .A(n477), .B(n476), .ZN(n510) );
  XNOR2_X1 U582 ( .A(n478), .B(n510), .ZN(n637) );
  NAND2_X1 U583 ( .A1(n637), .A2(n479), .ZN(n480) );
  INV_X1 U584 ( .A(G472), .ZN(n636) );
  NOR2_X1 U585 ( .A1(G900), .A2(n750), .ZN(n481) );
  NAND2_X1 U586 ( .A1(n481), .A2(G902), .ZN(n482) );
  NAND2_X1 U587 ( .A1(n750), .A2(G952), .ZN(n567) );
  NAND2_X1 U588 ( .A1(n482), .A2(n567), .ZN(n489) );
  NAND2_X1 U589 ( .A1(G234), .A2(n618), .ZN(n483) );
  XNOR2_X1 U590 ( .A(KEYINPUT20), .B(n483), .ZN(n501) );
  AND2_X1 U591 ( .A1(n501), .A2(G221), .ZN(n485) );
  INV_X1 U592 ( .A(KEYINPUT21), .ZN(n484) );
  XNOR2_X1 U593 ( .A(n485), .B(n484), .ZN(n664) );
  XNOR2_X1 U594 ( .A(KEYINPUT75), .B(KEYINPUT14), .ZN(n487) );
  XNOR2_X1 U595 ( .A(n487), .B(n486), .ZN(n694) );
  NOR2_X1 U596 ( .A1(n664), .A2(n694), .ZN(n488) );
  NAND2_X1 U597 ( .A1(n489), .A2(n488), .ZN(n519) );
  XOR2_X1 U598 ( .A(n519), .B(KEYINPUT70), .Z(n506) );
  XOR2_X1 U599 ( .A(KEYINPUT93), .B(KEYINPUT24), .Z(n491) );
  XNOR2_X1 U600 ( .A(n491), .B(n490), .ZN(n495) );
  XOR2_X1 U601 ( .A(KEYINPUT23), .B(KEYINPUT72), .Z(n493) );
  XNOR2_X1 U602 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U603 ( .A(n495), .B(n494), .Z(n499) );
  INV_X1 U604 ( .A(KEYINPUT69), .ZN(n496) );
  XNOR2_X1 U605 ( .A(n496), .B(G137), .ZN(n508) );
  XNOR2_X1 U606 ( .A(n497), .B(n508), .ZN(n498) );
  XOR2_X1 U607 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n503) );
  NAND2_X1 U608 ( .A1(n501), .A2(G217), .ZN(n502) );
  XNOR2_X1 U609 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U610 ( .A(n504), .B(KEYINPUT94), .ZN(n505) );
  NAND2_X1 U611 ( .A1(n506), .A2(n663), .ZN(n549) );
  XNOR2_X1 U612 ( .A(n508), .B(KEYINPUT90), .ZN(n509) );
  NAND2_X1 U613 ( .A1(n750), .A2(G227), .ZN(n511) );
  XNOR2_X1 U614 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U615 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U616 ( .A(n515), .B(n746), .ZN(n713) );
  INV_X1 U617 ( .A(G469), .ZN(n710) );
  NAND2_X1 U618 ( .A1(n696), .A2(n538), .ZN(n516) );
  INV_X1 U619 ( .A(n663), .ZN(n587) );
  INV_X1 U620 ( .A(n554), .ZN(n518) );
  INV_X1 U621 ( .A(n548), .ZN(n602) );
  NAND2_X1 U622 ( .A1(n602), .A2(n679), .ZN(n522) );
  XOR2_X1 U623 ( .A(KEYINPUT30), .B(KEYINPUT106), .Z(n520) );
  XNOR2_X1 U624 ( .A(n525), .B(KEYINPUT77), .ZN(n533) );
  NOR2_X1 U625 ( .A1(n533), .A2(n526), .ZN(n528) );
  INV_X1 U626 ( .A(KEYINPUT39), .ZN(n527) );
  INV_X1 U627 ( .A(n542), .ZN(n529) );
  OR2_X1 U628 ( .A1(n541), .A2(n529), .ZN(n550) );
  INV_X1 U629 ( .A(KEYINPUT109), .ZN(n530) );
  AND2_X1 U630 ( .A1(n541), .A2(n542), .ZN(n583) );
  NAND2_X1 U631 ( .A1(n583), .A2(n466), .ZN(n534) );
  NOR2_X1 U632 ( .A1(n533), .A2(n534), .ZN(n651) );
  NAND2_X1 U633 ( .A1(n535), .A2(n679), .ZN(n537) );
  INV_X1 U634 ( .A(KEYINPUT19), .ZN(n536) );
  XNOR2_X1 U635 ( .A(n537), .B(n536), .ZN(n566) );
  INV_X1 U636 ( .A(n541), .ZN(n543) );
  NOR2_X1 U637 ( .A1(n543), .A2(n542), .ZN(n657) );
  NAND2_X1 U638 ( .A1(n684), .A2(KEYINPUT47), .ZN(n544) );
  NAND2_X1 U639 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U640 ( .A(KEYINPUT111), .B(KEYINPUT36), .Z(n551) );
  XNOR2_X1 U641 ( .A(n552), .B(n551), .ZN(n555) );
  XNOR2_X1 U642 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n553) );
  XNOR2_X2 U643 ( .A(n554), .B(n553), .ZN(n668) );
  XNOR2_X1 U644 ( .A(n668), .B(KEYINPUT88), .ZN(n588) );
  OR2_X1 U645 ( .A1(n555), .A2(n588), .ZN(n662) );
  XOR2_X1 U646 ( .A(n684), .B(KEYINPUT84), .Z(n606) );
  NOR2_X1 U647 ( .A1(n556), .A2(KEYINPUT47), .ZN(n557) );
  NAND2_X1 U648 ( .A1(n606), .A2(n557), .ZN(n558) );
  INV_X1 U649 ( .A(KEYINPUT112), .ZN(n559) );
  XNOR2_X1 U650 ( .A(n560), .B(n559), .ZN(n756) );
  XOR2_X1 U651 ( .A(KEYINPUT105), .B(n561), .Z(n562) );
  AND2_X1 U652 ( .A1(n562), .A2(n668), .ZN(n563) );
  XNOR2_X1 U653 ( .A(n563), .B(KEYINPUT43), .ZN(n564) );
  NOR2_X1 U654 ( .A1(n564), .A2(n466), .ZN(n631) );
  NOR2_X1 U655 ( .A1(n756), .A2(n631), .ZN(n565) );
  NOR2_X1 U656 ( .A1(G898), .A2(n750), .ZN(n738) );
  NAND2_X1 U657 ( .A1(n738), .A2(G902), .ZN(n568) );
  NAND2_X1 U658 ( .A1(n568), .A2(n567), .ZN(n570) );
  INV_X1 U659 ( .A(n694), .ZN(n569) );
  INV_X1 U660 ( .A(n682), .ZN(n573) );
  INV_X1 U661 ( .A(n664), .ZN(n572) );
  NAND2_X1 U662 ( .A1(n573), .A2(n572), .ZN(n574) );
  INV_X1 U663 ( .A(n668), .ZN(n579) );
  INV_X1 U664 ( .A(KEYINPUT104), .ZN(n576) );
  AND2_X1 U665 ( .A1(n663), .A2(n667), .ZN(n577) );
  OR2_X1 U666 ( .A1(n663), .A2(n664), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n580), .A2(n579), .ZN(n581) );
  INV_X1 U668 ( .A(n600), .ZN(n605) );
  INV_X1 U669 ( .A(KEYINPUT80), .ZN(n584) );
  XNOR2_X1 U670 ( .A(n584), .B(KEYINPUT35), .ZN(n585) );
  OR2_X1 U671 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U672 ( .A(n589), .B(KEYINPUT103), .ZN(n591) );
  XNOR2_X1 U673 ( .A(n592), .B(KEYINPUT32), .ZN(n632) );
  NAND2_X1 U674 ( .A1(n593), .A2(n632), .ZN(n614) );
  NAND2_X1 U675 ( .A1(n614), .A2(KEYINPUT44), .ZN(n611) );
  OR2_X1 U676 ( .A1(n663), .A2(n594), .ZN(n595) );
  NOR2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U678 ( .A(n597), .B(KEYINPUT102), .ZN(n760) );
  NOR2_X1 U679 ( .A1(n598), .A2(n667), .ZN(n599) );
  NAND2_X1 U680 ( .A1(n599), .A2(n579), .ZN(n673) );
  OR2_X1 U681 ( .A1(n673), .A2(n600), .ZN(n601) );
  XNOR2_X1 U682 ( .A(n601), .B(KEYINPUT31), .ZN(n658) );
  NOR2_X1 U683 ( .A1(n598), .A2(n602), .ZN(n603) );
  AND2_X1 U684 ( .A1(n603), .A2(n518), .ZN(n604) );
  AND2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n644) );
  OR2_X1 U686 ( .A1(n658), .A2(n644), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U688 ( .A(n608), .B(KEYINPUT101), .ZN(n609) );
  NOR2_X1 U689 ( .A1(n760), .A2(n609), .ZN(n610) );
  NAND2_X1 U690 ( .A1(n611), .A2(n610), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n613), .B(n612), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n615), .A2(n423), .ZN(n617) );
  INV_X1 U693 ( .A(KEYINPUT45), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n620), .A2(KEYINPUT2), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n717) );
  INV_X1 U696 ( .A(n717), .ZN(n720) );
  NAND2_X1 U697 ( .A1(n720), .A2(G210), .ZN(n627) );
  XOR2_X1 U698 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n625) );
  BUF_X1 U699 ( .A(n623), .Z(n624) );
  XOR2_X1 U700 ( .A(n625), .B(n624), .Z(n626) );
  XNOR2_X1 U701 ( .A(n627), .B(n626), .ZN(n629) );
  INV_X1 U702 ( .A(G952), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n630), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U704 ( .A(G140), .B(n631), .Z(G42) );
  XOR2_X1 U705 ( .A(G119), .B(KEYINPUT126), .Z(n633) );
  XOR2_X1 U706 ( .A(n633), .B(n632), .Z(G21) );
  XNOR2_X1 U707 ( .A(n634), .B(G110), .ZN(G12) );
  XNOR2_X1 U708 ( .A(n635), .B(G122), .ZN(G24) );
  NOR2_X1 U709 ( .A1(n717), .A2(n636), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n637), .B(KEYINPUT62), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X1 U712 ( .A1(n640), .A2(n727), .ZN(n642) );
  XNOR2_X1 U713 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(G57) );
  NAND2_X1 U715 ( .A1(n644), .A2(n655), .ZN(n643) );
  XNOR2_X1 U716 ( .A(n643), .B(G104), .ZN(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n646) );
  NAND2_X1 U718 ( .A1(n644), .A2(n657), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U720 ( .A(G107), .B(n647), .ZN(G9) );
  XOR2_X1 U721 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n649) );
  INV_X1 U722 ( .A(n556), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n652), .A2(n657), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U725 ( .A(G128), .B(n650), .Z(G30) );
  XOR2_X1 U726 ( .A(G143), .B(n651), .Z(G45) );
  NAND2_X1 U727 ( .A1(n652), .A2(n655), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n653), .B(KEYINPUT114), .ZN(n654) );
  XNOR2_X1 U729 ( .A(G146), .B(n654), .ZN(G48) );
  NAND2_X1 U730 ( .A1(n658), .A2(n655), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n656), .B(G113), .ZN(G15) );
  XOR2_X1 U732 ( .A(G116), .B(KEYINPUT115), .Z(n660) );
  NAND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U734 ( .A(n660), .B(n659), .ZN(G18) );
  XOR2_X1 U735 ( .A(G125), .B(KEYINPUT37), .Z(n661) );
  XNOR2_X1 U736 ( .A(n662), .B(n661), .ZN(G27) );
  XOR2_X1 U737 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n709) );
  INV_X1 U738 ( .A(n696), .ZN(n678) );
  NAND2_X1 U739 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U740 ( .A(KEYINPUT49), .B(n665), .Z(n666) );
  NAND2_X1 U741 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n668), .A2(n598), .ZN(n669) );
  XOR2_X1 U743 ( .A(n669), .B(KEYINPUT50), .Z(n670) );
  NOR2_X1 U744 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U745 ( .A(KEYINPUT117), .B(n672), .ZN(n674) );
  NAND2_X1 U746 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U747 ( .A(n675), .B(KEYINPUT51), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n676), .B(KEYINPUT118), .ZN(n677) );
  NOR2_X1 U749 ( .A1(n678), .A2(n677), .ZN(n691) );
  NOR2_X1 U750 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n687) );
  NOR2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U753 ( .A(KEYINPUT119), .B(n685), .Z(n686) );
  NOR2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n689) );
  NOR2_X1 U755 ( .A1(n689), .A2(n366), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U757 ( .A(n692), .B(KEYINPUT52), .ZN(n693) );
  NOR2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U759 ( .A1(n695), .A2(G952), .ZN(n698) );
  NAND2_X1 U760 ( .A1(n696), .A2(n688), .ZN(n697) );
  NAND2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U762 ( .A1(G953), .A2(n699), .ZN(n707) );
  NOR2_X1 U763 ( .A1(n620), .A2(KEYINPUT85), .ZN(n700) );
  XNOR2_X1 U764 ( .A(n700), .B(KEYINPUT2), .ZN(n705) );
  INV_X1 U765 ( .A(n702), .ZN(n728) );
  NAND2_X1 U766 ( .A1(n701), .A2(n728), .ZN(n703) );
  NAND2_X1 U767 ( .A1(n703), .A2(KEYINPUT85), .ZN(n704) );
  NAND2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U770 ( .A(n709), .B(n708), .ZN(G75) );
  XNOR2_X1 U771 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n711) );
  XOR2_X1 U772 ( .A(n711), .B(KEYINPUT57), .Z(n712) );
  XNOR2_X1 U773 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U774 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U775 ( .A1(n727), .A2(n716), .ZN(G54) );
  XOR2_X1 U776 ( .A(n718), .B(KEYINPUT59), .Z(n719) );
  NAND2_X1 U777 ( .A1(n723), .A2(G478), .ZN(n721) );
  NAND2_X1 U778 ( .A1(n723), .A2(G217), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U780 ( .A1(n727), .A2(n726), .ZN(G66) );
  XNOR2_X1 U781 ( .A(KEYINPUT124), .B(KEYINPUT123), .ZN(n742) );
  NAND2_X1 U782 ( .A1(n728), .A2(n750), .ZN(n733) );
  NAND2_X1 U783 ( .A1(G224), .A2(G953), .ZN(n729) );
  XNOR2_X1 U784 ( .A(n729), .B(KEYINPUT122), .ZN(n730) );
  XNOR2_X1 U785 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U786 ( .A1(G898), .A2(n731), .ZN(n732) );
  NAND2_X1 U787 ( .A1(n733), .A2(n732), .ZN(n740) );
  XNOR2_X1 U788 ( .A(n734), .B(G101), .ZN(n735) );
  XNOR2_X1 U789 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U790 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U791 ( .A(n740), .B(n739), .Z(n741) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(G69) );
  XNOR2_X1 U793 ( .A(n743), .B(n744), .ZN(n745) );
  XNOR2_X1 U794 ( .A(n746), .B(n745), .ZN(n748) );
  XNOR2_X1 U795 ( .A(n748), .B(n701), .ZN(n747) );
  NAND2_X1 U796 ( .A1(n747), .A2(n750), .ZN(n753) );
  XNOR2_X1 U797 ( .A(n748), .B(G227), .ZN(n749) );
  NOR2_X1 U798 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U799 ( .A1(G900), .A2(n751), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U801 ( .A(KEYINPUT125), .B(n754), .ZN(G72) );
  XOR2_X1 U802 ( .A(G134), .B(KEYINPUT116), .Z(n755) );
  XNOR2_X1 U803 ( .A(n756), .B(n755), .ZN(G36) );
  XNOR2_X1 U804 ( .A(G137), .B(n757), .ZN(n758) );
  XNOR2_X1 U805 ( .A(n758), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U806 ( .A(n759), .B(G131), .Z(G33) );
  XOR2_X1 U807 ( .A(G101), .B(n760), .Z(G3) );
endmodule

