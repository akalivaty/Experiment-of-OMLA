//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT86), .B(G469), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n190), .B(KEYINPUT11), .C1(new_n191), .C2(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G134), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n189), .B1(new_n196), .B2(new_n200), .ZN(new_n201));
  AOI211_X1 g015(.A(KEYINPUT66), .B(new_n199), .C1(new_n194), .C2(new_n195), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n198), .A2(G134), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n203), .B1(new_n194), .B2(new_n195), .ZN(new_n204));
  OAI22_X1  g018(.A1(new_n201), .A2(new_n202), .B1(new_n197), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n206), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n209));
  XNOR2_X1  g023(.A(G143), .B(G146), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT84), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT84), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n216), .B1(G143), .B2(new_n207), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n214), .B(new_n215), .C1(new_n206), .C2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n208), .A2(new_n213), .A3(new_n216), .A4(G128), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT83), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n210), .A2(KEYINPUT83), .A3(new_n216), .A4(G128), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n211), .A2(new_n218), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  INV_X1    g038(.A(G107), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G104), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G107), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT3), .B1(new_n227), .B2(G107), .ZN(new_n230));
  AOI21_X1  g044(.A(G101), .B1(new_n227), .B2(G107), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n225), .A3(G104), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT81), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT81), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n230), .A2(new_n231), .A3(new_n233), .A4(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n229), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n223), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT69), .A2(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT69), .A2(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n214), .B1(new_n242), .B2(new_n217), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n219), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n205), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT12), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT12), .B(new_n205), .C1(new_n239), .C2(new_n245), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n223), .A2(new_n238), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT10), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n235), .A2(new_n237), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n230), .A2(new_n233), .A3(new_n228), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(G101), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n208), .A2(new_n213), .A3(KEYINPUT0), .A4(G128), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT0), .B(G128), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n210), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n255), .A2(G101), .ZN(new_n261));
  XOR2_X1   g075(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n251), .A2(new_n252), .B1(new_n257), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n191), .A2(G137), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n197), .B1(new_n196), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n195), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n198), .A2(G134), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT11), .B1(new_n268), .B2(new_n190), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n200), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT66), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n196), .A2(new_n189), .A3(new_n200), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n266), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n252), .B1(new_n243), .B2(new_n219), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT85), .B1(new_n238), .B2(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n238), .A2(KEYINPUT85), .A3(new_n274), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n264), .B(new_n273), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  XOR2_X1   g091(.A(G110), .B(G140), .Z(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(KEYINPUT80), .ZN(new_n279));
  AND2_X1   g093(.A1(KEYINPUT72), .A2(G953), .ZN(new_n280));
  NOR2_X1   g094(.A1(KEYINPUT72), .A2(G953), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G227), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n279), .B(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n250), .A2(new_n277), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n257), .A2(new_n263), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n239), .B2(KEYINPUT10), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n276), .A2(new_n275), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n205), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n284), .B1(new_n289), .B2(new_n277), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT87), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n285), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI211_X1 g106(.A(KEYINPUT87), .B(new_n284), .C1(new_n289), .C2(new_n277), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n187), .B(new_n188), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n284), .B1(new_n250), .B2(new_n277), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n289), .A2(new_n277), .A3(new_n284), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n187), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G469), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT9), .B(G234), .ZN(new_n300));
  OAI21_X1  g114(.A(G221), .B1(new_n300), .B2(G902), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G214), .B1(G237), .B2(G902), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(G110), .B(G122), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n305), .B(KEYINPUT88), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n255), .A2(G101), .A3(new_n262), .ZN(new_n308));
  OR2_X1    g122(.A1(KEYINPUT70), .A2(G119), .ZN(new_n309));
  NAND2_X1  g123(.A1(KEYINPUT70), .A2(G119), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(G116), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G116), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G119), .ZN(new_n313));
  INV_X1    g127(.A(G113), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G113), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n311), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n311), .B2(new_n313), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n308), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n253), .B2(new_n256), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n311), .A2(new_n313), .A3(new_n318), .ZN(new_n323));
  AND2_X1   g137(.A1(KEYINPUT70), .A2(G119), .ZN(new_n324));
  NOR2_X1   g138(.A1(KEYINPUT70), .A2(G119), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n324), .A2(new_n325), .A3(new_n312), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT5), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n314), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n311), .A2(KEYINPUT5), .A3(new_n313), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n238), .A2(new_n323), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n307), .B1(new_n322), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n318), .ZN(new_n333));
  INV_X1    g147(.A(new_n313), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(new_n326), .B2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n261), .A2(new_n262), .B1(new_n335), .B2(new_n323), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n257), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n324), .A2(new_n325), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n334), .B1(new_n338), .B2(G116), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n328), .A2(new_n329), .B1(new_n339), .B2(new_n318), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n238), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n341), .A3(new_n306), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n332), .A2(KEYINPUT6), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n260), .A2(G125), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(G125), .B2(new_n244), .ZN(new_n345));
  INV_X1    g159(.A(G224), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n346), .A2(G953), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT90), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n345), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT89), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n306), .B1(new_n337), .B2(new_n341), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n336), .A2(new_n257), .B1(new_n340), .B2(new_n238), .ZN(new_n354));
  NOR4_X1   g168(.A1(new_n354), .A2(KEYINPUT89), .A3(KEYINPUT6), .A4(new_n306), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n343), .B(new_n349), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n347), .A2(KEYINPUT7), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n345), .A2(new_n357), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n345), .A2(new_n357), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n342), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n306), .B(KEYINPUT8), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n340), .A2(new_n238), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n361), .B1(new_n331), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(G902), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n356), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G210), .B1(G237), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n356), .A2(new_n364), .A3(new_n366), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n304), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G475), .A2(G902), .ZN(new_n371));
  OR2_X1    g185(.A1(KEYINPUT72), .A2(G953), .ZN(new_n372));
  INV_X1    g186(.A(G237), .ZN(new_n373));
  NAND2_X1  g187(.A1(KEYINPUT72), .A2(G953), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n372), .A2(G214), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n212), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n282), .A2(G143), .A3(G214), .A4(new_n373), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G131), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT92), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT17), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n382), .A3(G131), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n376), .A2(new_n377), .A3(new_n197), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n380), .A2(new_n381), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(G125), .B(G140), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT16), .ZN(new_n387));
  INV_X1    g201(.A(G125), .ZN(new_n388));
  OR3_X1    g202(.A1(new_n388), .A2(KEYINPUT16), .A3(G140), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n207), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(G146), .A3(new_n389), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n382), .B1(new_n378), .B2(G131), .ZN(new_n395));
  AOI211_X1 g209(.A(KEYINPUT92), .B(new_n197), .C1(new_n376), .C2(new_n377), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT17), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n385), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G113), .B(G122), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(new_n227), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n378), .A2(KEYINPUT18), .A3(G131), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n386), .A2(KEYINPUT76), .A3(new_n207), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT76), .B1(new_n386), .B2(new_n207), .ZN(new_n403));
  OAI22_X1  g217(.A1(new_n402), .A2(new_n403), .B1(new_n207), .B2(new_n386), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT18), .A2(G131), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n376), .A2(new_n377), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT91), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT91), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n401), .A2(new_n404), .A3(new_n409), .A4(new_n406), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n398), .A2(new_n400), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n380), .A2(new_n383), .A3(new_n384), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n386), .B(KEYINPUT19), .Z(new_n414));
  MUX2_X1   g228(.A(new_n390), .B(new_n414), .S(new_n207), .Z(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n400), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n371), .B1(new_n412), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT20), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n411), .A2(new_n416), .ZN(new_n420));
  INV_X1    g234(.A(new_n400), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n398), .A2(new_n400), .A3(new_n411), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n371), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n400), .B1(new_n398), .B2(new_n411), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n187), .B1(new_n412), .B2(new_n427), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n419), .A2(new_n426), .B1(G475), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT93), .ZN(new_n430));
  INV_X1    g244(.A(G122), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n430), .B1(new_n431), .B2(G116), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n312), .A2(KEYINPUT93), .A3(G122), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(G116), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n434), .A2(new_n225), .A3(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n240), .A2(new_n241), .A3(new_n212), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n206), .A2(G143), .ZN(new_n438));
  OAI21_X1  g252(.A(G134), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n242), .A2(G143), .ZN(new_n440));
  INV_X1    g254(.A(new_n438), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n191), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n436), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n434), .A2(KEYINPUT14), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n435), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n434), .A2(KEYINPUT14), .ZN(new_n446));
  OAI21_X1  g260(.A(G107), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT13), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n440), .B(new_n441), .C1(new_n449), .C2(new_n191), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n437), .A2(KEYINPUT13), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n225), .B1(new_n434), .B2(new_n435), .ZN(new_n452));
  OAI221_X1 g266(.A(new_n450), .B1(new_n439), .B2(new_n451), .C1(new_n452), .C2(new_n436), .ZN(new_n453));
  INV_X1    g267(.A(G217), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n300), .A2(new_n454), .A3(G953), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT94), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n448), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n456), .B1(new_n448), .B2(new_n453), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n187), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT95), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(KEYINPUT95), .B(new_n187), .C1(new_n458), .C2(new_n459), .ZN(new_n463));
  INV_X1    g277(.A(G478), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n460), .A2(new_n465), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G952), .ZN(new_n469));
  AOI211_X1 g283(.A(G953), .B(new_n469), .C1(G234), .C2(G237), .ZN(new_n470));
  AOI211_X1 g284(.A(new_n187), .B(new_n282), .C1(G234), .C2(G237), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(G898), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n370), .A2(new_n429), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n302), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n392), .B1(new_n403), .B2(new_n402), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT23), .ZN(new_n478));
  OR2_X1    g292(.A1(KEYINPUT69), .A2(G128), .ZN(new_n479));
  NAND2_X1  g293(.A1(KEYINPUT69), .A2(G128), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(G119), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n309), .A2(G128), .A3(new_n310), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n309), .A2(new_n310), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT23), .B1(new_n484), .B2(new_n206), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n483), .A2(new_n485), .A3(G110), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n481), .A2(new_n482), .ZN(new_n487));
  XOR2_X1   g301(.A(KEYINPUT24), .B(G110), .Z(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT75), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G110), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n478), .B1(new_n338), .B2(G128), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n491), .B(new_n492), .C1(new_n487), .C2(new_n478), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n487), .A2(new_n488), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT75), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n477), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G110), .B1(new_n483), .B2(new_n485), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n487), .A2(new_n488), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n393), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT22), .B(G137), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT77), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT78), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n502), .A2(KEYINPUT77), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT78), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(KEYINPUT77), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n282), .A2(G221), .A3(G234), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n504), .B2(new_n508), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n497), .A2(new_n501), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n477), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n495), .B1(new_n493), .B2(new_n494), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n486), .A2(new_n489), .A3(KEYINPUT75), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n510), .A2(new_n511), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n500), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n512), .A2(new_n518), .A3(new_n187), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT25), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n512), .A2(new_n518), .A3(new_n521), .A4(new_n187), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n454), .B1(G234), .B2(new_n187), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(G902), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n512), .A2(new_n518), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT79), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n526), .A2(KEYINPUT79), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G472), .A2(G902), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT67), .B1(new_n191), .B2(G137), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n532), .A2(new_n203), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT67), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n191), .A3(G137), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G131), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT68), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n268), .A2(new_n265), .A3(KEYINPUT67), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT68), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n538), .A2(new_n539), .A3(G131), .A4(new_n535), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n541), .B(new_n244), .C1(new_n201), .C2(new_n202), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n542), .B(KEYINPUT30), .C1(new_n273), .C2(new_n260), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n319), .A2(new_n320), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n260), .B(KEYINPUT64), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n271), .A2(new_n272), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n537), .A2(new_n540), .B1(new_n219), .B2(new_n243), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n205), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n543), .B(new_n545), .C1(new_n549), .C2(KEYINPUT30), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n542), .B(new_n544), .C1(new_n273), .C2(new_n260), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n260), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n205), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n555), .A2(KEYINPUT71), .A3(new_n544), .A4(new_n542), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n282), .A2(G210), .A3(new_n373), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT27), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT26), .B(G101), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n550), .A2(new_n553), .A3(new_n556), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT31), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n553), .A2(new_n556), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT31), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n560), .A4(new_n550), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n551), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(KEYINPUT28), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT64), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n260), .B(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n542), .B1(new_n273), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n545), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n553), .A2(new_n572), .A3(new_n556), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n568), .B1(new_n573), .B2(KEYINPUT28), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(new_n560), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n531), .B1(new_n566), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT73), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT32), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n562), .B(new_n565), .C1(new_n574), .C2(new_n560), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(KEYINPUT73), .A3(new_n531), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G472), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n574), .A2(new_n560), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n550), .A2(new_n553), .A3(new_n556), .ZN(new_n585));
  INV_X1    g399(.A(new_n560), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT29), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n555), .A2(new_n542), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n545), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n553), .A3(new_n556), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n568), .B1(new_n591), .B2(KEYINPUT28), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n560), .A2(KEYINPUT29), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n583), .B1(new_n588), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n579), .A2(G472), .A3(G902), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n580), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT74), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT74), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n580), .A2(new_n600), .A3(new_n597), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n596), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n476), .B(new_n530), .C1(new_n582), .C2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NAND2_X1  g418(.A1(new_n580), .A2(new_n187), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(G472), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n606), .A2(new_n578), .A3(new_n581), .ZN(new_n607));
  INV_X1    g421(.A(new_n301), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n294), .B2(new_n298), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n530), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n428), .A2(G475), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n425), .B1(new_n424), .B2(new_n371), .ZN(new_n612));
  INV_X1    g426(.A(new_n371), .ZN(new_n613));
  AOI211_X1 g427(.A(KEYINPUT20), .B(new_n613), .C1(new_n422), .C2(new_n423), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n611), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n458), .A2(new_n459), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n457), .B2(new_n618), .ZN(new_n619));
  OR2_X1    g433(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n616), .A2(new_n619), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n620), .A2(G478), .A3(new_n187), .A4(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n615), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n368), .A2(KEYINPUT96), .A3(new_n369), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n366), .B1(new_n356), .B2(new_n364), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT96), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n304), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n625), .A2(new_n630), .A3(new_n473), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n610), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT98), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT99), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NAND3_X1  g451(.A1(new_n419), .A2(new_n426), .A3(KEYINPUT100), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n612), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n638), .A2(new_n611), .A3(new_n468), .A4(new_n640), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n641), .A2(new_n630), .A3(new_n473), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n610), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT35), .B(G107), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NAND2_X1  g460(.A1(new_n516), .A2(new_n500), .ZN(new_n647));
  OR3_X1    g461(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT36), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(new_n525), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n524), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n429), .A2(new_n474), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n607), .A2(new_n609), .A3(new_n370), .A4(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NAND3_X1  g471(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n580), .A2(new_n600), .A3(new_n597), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n600), .B1(new_n580), .B2(new_n597), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n658), .A2(new_n661), .A3(new_n596), .ZN(new_n662));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n470), .B1(new_n471), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n641), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n626), .A2(new_n652), .A3(new_n629), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n302), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n662), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G128), .ZN(G30));
  NAND2_X1  g483(.A1(new_n615), .A2(new_n468), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n670), .A2(new_n304), .A3(new_n652), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n368), .A2(new_n369), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n664), .B(KEYINPUT39), .Z(new_n677));
  AND2_X1   g491(.A1(new_n609), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n675), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n585), .A2(new_n560), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n680), .B(new_n187), .C1(new_n560), .C2(new_n591), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G472), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n599), .A2(new_n601), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n658), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n679), .B(new_n685), .C1(new_n676), .C2(new_n678), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  INV_X1    g501(.A(new_n664), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n615), .A2(new_n624), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n667), .B(new_n690), .C1(new_n582), .C2(new_n602), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  OAI21_X1  g506(.A(new_n187), .B1(new_n292), .B2(new_n293), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G469), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n301), .A3(new_n294), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n662), .A2(new_n530), .A3(new_n631), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND4_X1  g513(.A1(new_n662), .A2(new_n530), .A3(new_n642), .A4(new_n696), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT102), .B(G116), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G18));
  NOR3_X1   g516(.A1(new_n695), .A2(new_n653), .A3(new_n630), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n662), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  INV_X1    g519(.A(new_n473), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n694), .A2(new_n301), .A3(new_n294), .A4(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n615), .A2(new_n626), .A3(new_n468), .A4(new_n629), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT103), .B(G472), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n605), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n592), .A2(new_n560), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n531), .B1(new_n566), .B2(new_n712), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n711), .A2(new_n530), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  NAND3_X1  g530(.A1(new_n711), .A2(new_n652), .A3(new_n713), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n695), .A2(new_n630), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n719), .A3(new_n690), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT104), .B(G125), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G27));
  NOR3_X1   g536(.A1(new_n659), .A2(new_n660), .A3(new_n595), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n529), .B1(new_n723), .B2(new_n658), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n368), .A2(new_n303), .A3(new_n369), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n368), .A2(KEYINPUT105), .A3(new_n303), .A4(new_n369), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n609), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT106), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n609), .A2(new_n727), .A3(new_n731), .A4(new_n728), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n724), .A2(new_n690), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n730), .A2(new_n732), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n580), .A2(new_n597), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n595), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n576), .A2(new_n579), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n529), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n689), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n733), .A2(new_n734), .B1(new_n735), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n197), .ZN(G33));
  NAND3_X1  g558(.A1(new_n735), .A2(new_n724), .A3(new_n665), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  NAND2_X1  g560(.A1(new_n429), .A2(new_n624), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(KEYINPUT43), .Z(new_n748));
  INV_X1    g562(.A(new_n607), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n652), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(G469), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n295), .A2(new_n296), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n756), .B1(new_n755), .B2(new_n754), .ZN(new_n757));
  NAND2_X1  g571(.A1(G469), .A2(G902), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT46), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n294), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n758), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n608), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(new_n677), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n750), .A2(new_n751), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n727), .A2(new_n728), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT108), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n752), .A2(new_n764), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n763), .A2(new_n771), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n763), .B1(new_n773), .B2(new_n771), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n662), .A2(new_n530), .A3(new_n689), .A4(new_n766), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  AND2_X1   g591(.A1(new_n748), .A2(new_n470), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(new_n714), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n674), .A2(new_n303), .A3(new_n695), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT50), .Z(new_n782));
  NAND2_X1  g596(.A1(new_n772), .A2(new_n774), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n694), .A2(new_n294), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n608), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n767), .A3(new_n779), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n766), .A2(new_n695), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n778), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n685), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n530), .A2(new_n791), .A3(new_n470), .A4(new_n788), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n615), .A2(new_n624), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n790), .A2(new_n718), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n782), .A2(new_n787), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n790), .A2(new_n739), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT48), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n798), .A2(KEYINPUT116), .A3(new_n799), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n469), .B(G953), .C1(new_n779), .C2(new_n719), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n792), .A2(new_n615), .A3(new_n624), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n800), .B(new_n803), .C1(new_n798), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n795), .A2(new_n796), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n797), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n672), .A2(new_n303), .A3(new_n706), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n429), .A2(new_n468), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n808), .B1(new_n809), .B2(new_n625), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n607), .A2(new_n810), .A3(new_n530), .A4(new_n609), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n603), .A2(new_n655), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n717), .A2(new_n689), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n730), .A3(new_n732), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n609), .A2(new_n727), .A3(new_n728), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n611), .A2(new_n467), .A3(new_n466), .A4(new_n688), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n640), .A2(new_n816), .A3(new_n638), .A4(new_n652), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n815), .B(new_n817), .C1(new_n582), .C2(new_n602), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n812), .A2(new_n819), .A3(new_n745), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n662), .A2(new_n703), .B1(new_n709), .B2(new_n714), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n697), .A3(new_n700), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n820), .A2(new_n743), .A3(KEYINPUT112), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n733), .A2(new_n734), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n742), .A2(new_n735), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n662), .A2(new_n730), .A3(new_n530), .A4(new_n732), .ZN(new_n828));
  INV_X1    g642(.A(new_n665), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n814), .B(new_n818), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n603), .A2(new_n811), .A3(new_n655), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n824), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n823), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n664), .B(KEYINPUT113), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n524), .A2(new_n651), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n302), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n708), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n837), .B(new_n838), .C1(new_n582), .C2(new_n683), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n668), .A2(new_n691), .A3(new_n839), .A4(new_n720), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n662), .B(new_n667), .C1(new_n665), .C2(new_n690), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(KEYINPUT52), .A3(new_n720), .A4(new_n839), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT53), .B1(new_n834), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n842), .B2(new_n844), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n823), .A2(new_n833), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT54), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n827), .A2(new_n832), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT112), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n827), .A2(new_n832), .A3(new_n824), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n845), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n847), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n812), .A2(new_n819), .A3(new_n745), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n827), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT114), .B1(new_n830), .B2(new_n831), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n848), .A4(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n848), .A2(new_n827), .A3(new_n861), .A4(new_n858), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT115), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n856), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n851), .A2(new_n867), .ZN(new_n868));
  OAI22_X1  g682(.A1(new_n807), .A2(new_n868), .B1(G952), .B2(G953), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT49), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n784), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT110), .Z(new_n872));
  NOR2_X1   g686(.A1(new_n784), .A2(new_n870), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n530), .A2(new_n301), .A3(new_n303), .ZN(new_n874));
  NOR4_X1   g688(.A1(new_n873), .A2(new_n747), .A3(new_n674), .A4(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n875), .A3(new_n791), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT111), .Z(new_n877));
  NAND2_X1  g691(.A1(new_n869), .A2(new_n877), .ZN(G75));
  NOR2_X1   g692(.A1(new_n282), .A2(G952), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n187), .B1(new_n856), .B2(new_n865), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT56), .B1(new_n881), .B2(G210), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n343), .B1(new_n353), .B2(new_n355), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(new_n349), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT55), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n880), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n863), .B(new_n860), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n846), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n889), .B2(new_n187), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n881), .A2(KEYINPUT117), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n367), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n886), .B1(new_n892), .B2(new_n894), .ZN(G51));
  OAI21_X1  g709(.A(KEYINPUT54), .B1(new_n888), .B2(new_n846), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(KEYINPUT118), .A3(new_n867), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n898), .B(KEYINPUT54), .C1(new_n888), .C2(new_n846), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n758), .B(KEYINPUT57), .Z(new_n900));
  NAND3_X1  g714(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n293), .B2(new_n292), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n757), .B(KEYINPUT119), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n890), .A2(new_n891), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n879), .B1(new_n902), .B2(new_n904), .ZN(G54));
  AND2_X1   g719(.A1(KEYINPUT58), .A2(G475), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n890), .A2(new_n891), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n422), .A3(new_n423), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n890), .A2(new_n424), .A3(new_n891), .A4(new_n906), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n908), .A2(new_n880), .A3(new_n909), .ZN(G60));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n620), .A2(new_n621), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(G478), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT59), .Z(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n897), .A2(new_n899), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n851), .B2(new_n867), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n880), .B1(new_n918), .B2(new_n912), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n911), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n851), .A2(new_n867), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n913), .B1(new_n921), .B2(new_n915), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n897), .A2(new_n899), .A3(new_n916), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT120), .A4(new_n880), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n920), .A2(new_n924), .ZN(G63));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT60), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n889), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n928), .A2(new_n649), .A3(new_n650), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n512), .A2(new_n518), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT121), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n889), .B2(new_n927), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n929), .A2(new_n880), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n929), .A2(KEYINPUT61), .A3(new_n880), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(G66));
  NOR2_X1   g751(.A1(new_n822), .A2(new_n831), .ZN(new_n938));
  INV_X1    g752(.A(new_n282), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT122), .Z(new_n941));
  OAI21_X1  g755(.A(G953), .B1(new_n472), .B2(new_n346), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n883), .B1(G898), .B2(new_n282), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n768), .A2(new_n776), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n766), .B1(new_n625), .B2(new_n809), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n724), .A2(new_n678), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n843), .A2(new_n720), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n686), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(KEYINPUT62), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT123), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(KEYINPUT62), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n950), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  MUX2_X1   g770(.A(new_n549), .B(new_n589), .S(KEYINPUT30), .Z(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(new_n414), .Z(new_n958));
  NOR3_X1   g772(.A1(new_n956), .A2(new_n939), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(G227), .B2(new_n282), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n764), .A2(new_n838), .A3(new_n739), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n961), .A2(new_n745), .A3(new_n951), .ZN(new_n962));
  INV_X1    g776(.A(new_n743), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n947), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n960), .B1(new_n964), .B2(new_n282), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n946), .B1(new_n959), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(G227), .B1(new_n958), .B2(new_n946), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n939), .B1(new_n967), .B2(new_n663), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(G72));
  XNOR2_X1  g783(.A(new_n585), .B(new_n560), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  XOR2_X1   g785(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n972));
  NOR2_X1   g786(.A1(new_n583), .A2(new_n187), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n880), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n950), .A2(new_n954), .A3(new_n955), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n563), .A2(new_n586), .A3(new_n550), .ZN(new_n977));
  OAI22_X1  g791(.A1(new_n976), .A2(new_n680), .B1(new_n964), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n975), .B1(new_n978), .B2(new_n938), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n846), .A2(new_n850), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT126), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n971), .A2(new_n974), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n980), .B2(new_n982), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT127), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT127), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n979), .B(new_n987), .C1(new_n983), .C2(new_n984), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n988), .ZN(G57));
endmodule


