//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1169, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  OR2_X1    g0003(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n205));
  NAND3_X1  g0005(.A1(new_n204), .A2(G50), .A3(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  NOR3_X1   g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(new_n207), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G58), .B2(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  XOR2_X1   g0022(.A(KEYINPUT65), .B(G77), .Z(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n212), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n212), .A2(G13), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(KEYINPUT0), .ZN(new_n233));
  OR2_X1    g0033(.A1(new_n232), .A2(KEYINPUT0), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n209), .B(new_n230), .C1(new_n233), .C2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G226), .B(G232), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n217), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G222), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n252), .B(new_n254), .C1(new_n255), .C2(new_n253), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n256), .B(new_n260), .C1(new_n223), .C2(new_n252), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n262), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n261), .B(new_n265), .C1(new_n215), .C2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT67), .ZN(new_n268));
  INV_X1    g0068(.A(G200), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g0070(.A(new_n270), .B(KEYINPUT70), .Z(new_n271));
  INV_X1    g0071(.A(new_n203), .ZN(new_n272));
  OAI21_X1  g0072(.A(G20), .B1(new_n272), .B2(G50), .ZN(new_n273));
  INV_X1    g0073(.A(G150), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  XOR2_X1   g0076(.A(KEYINPUT8), .B(G58), .Z(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n257), .A2(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n273), .B1(new_n274), .B2(new_n276), .C1(new_n278), .C2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n208), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT68), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n210), .A2(G20), .ZN(new_n287));
  INV_X1    g0087(.A(G13), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n281), .A2(new_n286), .B1(new_n214), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n285), .A2(G50), .A3(new_n287), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n295));
  AOI211_X1 g0095(.A(new_n294), .B(new_n295), .C1(G190), .C2(new_n268), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT69), .B(KEYINPUT10), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n271), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n270), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n268), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n303), .B(new_n292), .C1(G169), .C2(new_n268), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n215), .A2(new_n253), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n252), .B(new_n305), .C1(G232), .C2(new_n253), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G97), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n259), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n266), .A2(new_n221), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n308), .A2(new_n264), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT13), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT71), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n311), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT72), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(G190), .A3(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n279), .A2(G77), .B1(new_n275), .B2(G50), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n207), .B2(G68), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n286), .A2(new_n318), .ZN(new_n319));
  XOR2_X1   g0119(.A(new_n319), .B(KEYINPUT11), .Z(new_n320));
  NOR2_X1   g0120(.A1(new_n289), .A2(new_n283), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(G68), .A3(new_n287), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT73), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n321), .A2(KEYINPUT73), .A3(G68), .A4(new_n287), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT12), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n288), .A2(G1), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(G20), .A3(new_n220), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n324), .A2(new_n325), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n326), .B2(new_n328), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n320), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n310), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(KEYINPUT13), .ZN(new_n333));
  OAI21_X1  g0133(.A(G200), .B1(new_n333), .B2(new_n312), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n316), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n331), .B(KEYINPUT74), .ZN(new_n336));
  OAI21_X1  g0136(.A(G169), .B1(new_n333), .B2(new_n312), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n337), .A2(KEYINPUT14), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n313), .A2(G179), .A3(new_n315), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(KEYINPUT14), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n335), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G238), .A2(G1698), .ZN(new_n343));
  INV_X1    g0143(.A(G232), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n252), .B(new_n343), .C1(new_n344), .C2(G1698), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n260), .C1(G107), .C2(new_n252), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(new_n265), .C1(new_n222), .C2(new_n266), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n347), .A2(G179), .ZN(new_n348));
  AOI22_X1  g0148(.A1(G20), .A2(new_n223), .B1(new_n277), .B2(new_n275), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT15), .B(G87), .Z(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n349), .B1(new_n280), .B2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(new_n283), .B1(new_n224), .B2(new_n289), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n321), .A2(G77), .A3(new_n287), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n347), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n348), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n301), .A2(new_n304), .A3(new_n342), .A4(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n283), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(new_n207), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT3), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n257), .ZN(new_n366));
  NAND2_X1  g0166(.A1(KEYINPUT3), .A2(G33), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G68), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G58), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(new_n220), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n372), .B2(new_n203), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n275), .A2(G159), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT76), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n373), .A2(KEYINPUT76), .A3(new_n374), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n370), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n360), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n373), .A2(KEYINPUT76), .A3(new_n374), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT76), .B1(new_n373), .B2(new_n374), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n366), .A2(new_n207), .A3(new_n367), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n368), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT75), .B1(new_n388), .B2(G68), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT75), .ZN(new_n390));
  AOI211_X1 g0190(.A(new_n390), .B(new_n220), .C1(new_n387), .C2(new_n368), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT16), .B(new_n384), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n381), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n255), .A2(new_n253), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n252), .B(new_n394), .C1(G226), .C2(new_n253), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n259), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n265), .B1(new_n266), .B2(new_n344), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G200), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(G190), .ZN(new_n402));
  INV_X1    g0202(.A(new_n287), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n277), .B1(new_n286), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n289), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n278), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n393), .A2(new_n401), .A3(new_n402), .A4(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT17), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n381), .A2(new_n392), .B1(new_n404), .B2(new_n406), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n411), .A2(KEYINPUT17), .A3(new_n401), .A4(new_n402), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G190), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n347), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n347), .A2(G200), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n416), .A2(new_n353), .A3(new_n354), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n393), .A2(new_n407), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n397), .A2(new_n302), .A3(new_n398), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n400), .B2(G169), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT18), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n411), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n414), .B(new_n418), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n359), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n207), .B(G87), .C1(new_n361), .C2(new_n362), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT22), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT22), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n252), .A2(new_n430), .A3(new_n207), .A4(G87), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT82), .B(G116), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n279), .ZN(new_n434));
  INV_X1    g0234(.A(G107), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G20), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT23), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n432), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT24), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n432), .A2(KEYINPUT24), .A3(new_n434), .A4(new_n438), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n283), .A3(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n285), .B(new_n405), .C1(G1), .C2(new_n257), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G107), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  OR2_X1    g0247(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n448));
  NAND2_X1  g0248(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n289), .A2(new_n435), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(KEYINPUT87), .B(KEYINPUT25), .C1(new_n405), .C2(G107), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n252), .A2(G257), .A3(G1698), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n252), .A2(G250), .A3(new_n253), .ZN(new_n453));
  XOR2_X1   g0253(.A(KEYINPUT88), .B(G294), .Z(new_n454));
  OAI211_X1 g0254(.A(new_n452), .B(new_n453), .C1(new_n257), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n260), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT79), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(new_n258), .A3(KEYINPUT5), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT5), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(KEYINPUT79), .B2(G41), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n458), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n263), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n463), .A2(new_n259), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G264), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n456), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n269), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n455), .A2(new_n260), .B1(G264), .B2(new_n466), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(new_n415), .A3(new_n465), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n447), .A2(new_n450), .A3(new_n451), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n405), .A2(G97), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n444), .B2(new_n226), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT6), .ZN(new_n477));
  AND2_X1   g0277(.A1(G97), .A2(G107), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n435), .A2(KEYINPUT6), .A3(G97), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G20), .ZN(new_n483));
  INV_X1    g0283(.A(G77), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n276), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n435), .B1(new_n387), .B2(new_n368), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n283), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT77), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n388), .A2(G107), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n482), .A2(G20), .B1(G77), .B2(new_n275), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n360), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT77), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n476), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G250), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n363), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT4), .ZN(new_n497));
  OAI21_X1  g0297(.A(G1698), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT78), .ZN(new_n499));
  OAI21_X1  g0299(.A(G244), .B1(new_n361), .B2(new_n362), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(new_n497), .B1(G33), .B2(G283), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n253), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n498), .A2(new_n499), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(new_n497), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n252), .A2(G250), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n253), .B1(new_n507), .B2(KEYINPUT4), .ZN(new_n508));
  OAI21_X1  g0308(.A(KEYINPUT78), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n260), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n466), .A2(KEYINPUT80), .A3(G257), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT80), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n463), .A2(new_n259), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n227), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n464), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n511), .A2(G190), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n259), .B1(new_n503), .B2(new_n509), .ZN(new_n518));
  INV_X1    g0318(.A(new_n516), .ZN(new_n519));
  OAI21_X1  g0319(.A(G200), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n494), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n511), .A2(new_n302), .A3(new_n516), .ZN(new_n522));
  INV_X1    g0322(.A(new_n476), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n491), .A2(new_n492), .ZN(new_n524));
  AOI211_X1 g0324(.A(KEYINPUT77), .B(new_n360), .C1(new_n489), .C2(new_n490), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n356), .B1(new_n518), .B2(new_n519), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n473), .A2(new_n521), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(G116), .B1(new_n257), .B2(G1), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n289), .A2(new_n283), .A3(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n505), .B(new_n207), .C1(G33), .C2(new_n226), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n283), .B(new_n532), .C1(new_n433), .C2(new_n207), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT20), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n216), .A2(KEYINPUT82), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT82), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G116), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G20), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n540), .A2(KEYINPUT20), .A3(new_n283), .A4(new_n532), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n531), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(G20), .A3(new_n327), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(G264), .A2(G1698), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n361), .B2(new_n362), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT85), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n252), .A2(G257), .A3(new_n253), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n363), .A2(G303), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT85), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n550), .B(new_n545), .C1(new_n361), .C2(new_n362), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n260), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n464), .B1(new_n466), .B2(G270), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT86), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT86), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(G200), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n558), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n557), .B1(new_n553), .B2(new_n554), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n544), .B(new_n559), .C1(new_n562), .C2(new_n415), .ZN(new_n563));
  OR3_X1    g0363(.A1(new_n544), .A2(new_n302), .A3(new_n555), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n356), .B1(new_n542), .B2(new_n543), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n556), .A2(new_n565), .A3(KEYINPUT21), .A4(new_n558), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n556), .A2(new_n565), .A3(new_n558), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n563), .A2(new_n564), .A3(new_n566), .A4(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n443), .A2(new_n450), .A3(new_n451), .A4(new_n446), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n470), .A2(new_n302), .A3(new_n465), .ZN(new_n572));
  AOI21_X1  g0372(.A(G169), .B1(new_n470), .B2(new_n465), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n529), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT84), .ZN(new_n577));
  OAI211_X1 g0377(.A(G244), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT81), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT81), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n252), .A2(new_n580), .A3(G244), .A4(G1698), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n252), .A2(G238), .A3(new_n253), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n433), .A2(G33), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n260), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n462), .A2(new_n263), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n495), .B1(new_n461), .B2(G1), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n259), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n589), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n579), .A2(new_n581), .A3(new_n584), .A4(new_n583), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(new_n260), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT83), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n269), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n252), .A2(new_n207), .A3(G68), .ZN(new_n598));
  INV_X1    g0398(.A(G87), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n479), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n307), .A2(new_n207), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(KEYINPUT19), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n307), .A2(G20), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n598), .B(new_n602), .C1(KEYINPUT19), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n283), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n351), .A2(new_n289), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n599), .B2(new_n444), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n577), .B1(new_n597), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n592), .A2(G190), .A3(new_n596), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n607), .B1(G87), .B2(new_n445), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT83), .B1(new_n586), .B2(new_n589), .ZN(new_n613));
  AOI211_X1 g0413(.A(new_n591), .B(new_n593), .C1(new_n594), .C2(new_n260), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(KEYINPUT84), .B(new_n612), .C1(new_n615), .C2(new_n269), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n610), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n302), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n608), .B1(new_n444), .B2(new_n351), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n618), .B(new_n619), .C1(G169), .C2(new_n615), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n427), .A2(new_n576), .A3(new_n621), .ZN(G372));
  NAND2_X1  g0422(.A1(new_n341), .A2(new_n336), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n335), .B2(new_n358), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n624), .A2(new_n414), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n423), .A2(new_n425), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n301), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n304), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n569), .A2(new_n566), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT89), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n571), .A2(new_n574), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n564), .A4(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n473), .A2(new_n521), .A3(new_n528), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n569), .A2(new_n564), .A3(new_n566), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT89), .B1(new_n635), .B2(new_n575), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n590), .A2(new_n356), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n618), .A2(new_n619), .A3(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n611), .B(new_n612), .C1(new_n269), .C2(new_n595), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n633), .A2(new_n634), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n617), .A2(new_n642), .A3(new_n620), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT26), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n642), .A2(new_n645), .A3(new_n638), .A4(new_n639), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n646), .A2(new_n638), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n641), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n427), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n629), .A2(new_n649), .ZN(G369));
  INV_X1    g0450(.A(new_n473), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n327), .A2(new_n207), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(G213), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n571), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n632), .B1(new_n651), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n657), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n575), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n635), .A2(new_n660), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(new_n661), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n544), .A2(new_n660), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n635), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n570), .B2(new_n666), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n662), .A2(G330), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(new_n231), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n600), .A2(G116), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n206), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(new_n638), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n640), .A2(new_n642), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(KEYINPUT26), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n634), .B(new_n640), .C1(new_n635), .C2(new_n575), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n680), .B(new_n681), .C1(KEYINPUT26), .C2(new_n643), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(KEYINPUT29), .A3(new_n660), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT91), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n648), .A2(new_n660), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n685), .B1(new_n683), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n511), .A2(new_n516), .A3(new_n470), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n555), .A2(new_n302), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n592), .A3(new_n596), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n691), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT30), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n691), .B(new_n697), .C1(new_n692), .C2(new_n694), .ZN(new_n698));
  AOI21_X1  g0498(.A(G179), .B1(new_n511), .B2(new_n516), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(new_n468), .A3(new_n562), .A4(new_n590), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n696), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n576), .A2(new_n621), .A3(new_n660), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n703), .A2(KEYINPUT31), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n701), .A2(new_n657), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n690), .B1(G330), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n677), .B1(new_n707), .B2(G1), .ZN(G364));
  OR2_X1    g0508(.A1(new_n668), .A2(G330), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n668), .A2(G330), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n288), .A2(G20), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G45), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n673), .A2(G1), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT92), .Z(new_n715));
  AOI21_X1  g0515(.A(new_n208), .B1(G20), .B2(new_n356), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n207), .A2(G190), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(new_n302), .A3(new_n269), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT94), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(KEYINPUT94), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n207), .A2(new_n302), .A3(new_n269), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G190), .ZN(new_n726));
  XNOR2_X1  g0526(.A(KEYINPUT33), .B(G317), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n723), .A2(G329), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G303), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n302), .A2(G200), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT95), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n207), .A2(new_n415), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n415), .A2(G179), .A3(G200), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n207), .ZN(new_n736));
  OAI221_X1 g0536(.A(new_n728), .B1(new_n729), .B2(new_n734), .C1(new_n454), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n731), .A2(new_n718), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n737), .B1(G283), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n725), .A2(new_n415), .ZN(new_n741));
  XOR2_X1   g0541(.A(KEYINPUT96), .B(G326), .Z(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n302), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n732), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G322), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(new_n718), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n252), .B1(new_n749), .B2(G311), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n740), .A2(new_n743), .A3(new_n747), .A4(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n741), .A2(G50), .B1(new_n223), .B2(new_n749), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n371), .B2(new_n745), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT93), .Z(new_n754));
  INV_X1    g0554(.A(G159), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n722), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT32), .ZN(new_n757));
  INV_X1    g0557(.A(new_n726), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n734), .A2(new_n599), .B1(new_n220), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n736), .A2(new_n226), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n738), .A2(new_n435), .ZN(new_n761));
  NOR4_X1   g0561(.A1(new_n759), .A2(new_n363), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n754), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n717), .B1(new_n751), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n668), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n231), .A2(G355), .A3(new_n252), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n671), .A2(new_n252), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(G45), .B2(new_n206), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n247), .A2(new_n461), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n770), .B1(G116), .B2(new_n231), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n767), .A2(new_n716), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n713), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n769), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n715), .B1(new_n764), .B2(new_n778), .ZN(G396));
  NAND2_X1  g0579(.A1(new_n706), .A2(G330), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n355), .A2(new_n657), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n418), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n358), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n358), .A2(new_n657), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n686), .B(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n780), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n713), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G68), .A2(new_n739), .B1(new_n733), .B2(G50), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G137), .A2(new_n741), .B1(new_n726), .B2(G150), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT97), .ZN(new_n793));
  INV_X1    g0593(.A(G143), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n793), .B1(new_n794), .B2(new_n745), .C1(new_n755), .C2(new_n748), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT34), .ZN(new_n796));
  INV_X1    g0596(.A(new_n736), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n790), .A2(KEYINPUT98), .B1(G58), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n796), .A2(new_n252), .A3(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n791), .B(new_n799), .C1(G132), .C2(new_n723), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n363), .B1(new_n599), .B2(new_n738), .C1(new_n734), .C2(new_n435), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  INV_X1    g0602(.A(new_n741), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n722), .A2(new_n802), .B1(new_n803), .B2(new_n729), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n801), .A2(new_n760), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n726), .A2(G283), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n805), .B(new_n806), .C1(new_n539), .C2(new_n748), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(G294), .B2(new_n746), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n716), .B1(new_n800), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n716), .A2(new_n765), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n484), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n785), .A2(new_n765), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n809), .A2(new_n777), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n789), .A2(new_n813), .ZN(G384));
  INV_X1    g0614(.A(new_n655), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n384), .B1(new_n389), .B2(new_n391), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n380), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n817), .A2(new_n286), .A3(new_n392), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n407), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n815), .B(new_n819), .C1(new_n626), .C2(new_n413), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n815), .B(new_n420), .C1(G169), .C2(new_n400), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n407), .B2(new_n818), .ZN(new_n822));
  INV_X1    g0622(.A(new_n408), .ZN(new_n823));
  OAI21_X1  g0623(.A(KEYINPUT37), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT37), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n408), .B(new_n825), .C1(new_n411), .C2(new_n821), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n820), .A2(new_n827), .A3(KEYINPUT38), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n419), .B(new_n815), .C1(new_n626), .C2(new_n413), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n408), .B1(new_n411), .B2(new_n821), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(KEYINPUT37), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n826), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT38), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n820), .A2(new_n827), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n828), .ZN(new_n839));
  MUX2_X1   g0639(.A(new_n835), .B(new_n839), .S(KEYINPUT39), .Z(new_n840));
  NOR2_X1   g0640(.A1(new_n623), .A2(new_n657), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n840), .A2(new_n841), .B1(new_n626), .B2(new_n655), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n648), .A2(new_n660), .A3(new_n786), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n784), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT101), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n843), .A2(KEYINPUT101), .A3(new_n784), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n316), .A2(new_n331), .A3(new_n334), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n336), .A2(new_n657), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n623), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n336), .B(new_n657), .C1(new_n335), .C2(new_n341), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n848), .A2(new_n839), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n842), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n628), .B1(new_n690), .B2(new_n427), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n705), .B1(new_n703), .B2(KEYINPUT31), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n702), .A2(KEYINPUT102), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT102), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n701), .A2(new_n860), .A3(KEYINPUT31), .A4(new_n657), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n835), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n785), .B1(new_n851), .B2(new_n852), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n863), .A2(KEYINPUT40), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n839), .B(new_n865), .C1(new_n858), .C2(new_n862), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT40), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT103), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT103), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n868), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n867), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(new_n427), .A3(new_n863), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n868), .A2(new_n872), .A3(new_n869), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n872), .B1(new_n868), .B2(new_n869), .ZN(new_n877));
  OAI211_X1 g0677(.A(G330), .B(new_n866), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n427), .A2(G330), .A3(new_n863), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n857), .B(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n210), .B2(new_n711), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n223), .B1(new_n371), .B2(new_n220), .ZN(new_n884));
  OAI22_X1  g0684(.A1(new_n884), .A2(new_n206), .B1(G50), .B2(new_n220), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(G1), .A3(new_n288), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT100), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n216), .B1(new_n482), .B2(KEYINPUT35), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n208), .A2(new_n207), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n888), .B(new_n889), .C1(KEYINPUT35), .C2(new_n482), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT99), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT36), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n883), .A2(new_n887), .A3(new_n892), .ZN(G367));
  OAI211_X1 g0693(.A(new_n521), .B(new_n528), .C1(new_n494), .C2(new_n660), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n664), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT42), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n528), .B1(new_n894), .B2(new_n632), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n660), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n640), .B1(new_n612), .B2(new_n660), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n678), .A2(new_n609), .A3(new_n657), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n896), .A2(new_n898), .B1(KEYINPUT43), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n669), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n894), .B1(new_n528), .B2(new_n660), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n904), .B(new_n907), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n672), .B(KEYINPUT41), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n662), .B(new_n663), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n905), .B1(new_n911), .B2(new_n710), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n707), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT104), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n665), .A2(new_n906), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT45), .Z(new_n916));
  NOR2_X1   g0716(.A1(new_n665), .A2(new_n906), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT44), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n913), .A2(new_n914), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n910), .B1(new_n920), .B2(new_n707), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n712), .A2(G1), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n908), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n901), .A2(new_n768), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n723), .A2(G137), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n797), .A2(G68), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n739), .A2(new_n223), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n726), .A2(G159), .B1(G50), .B2(new_n749), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT107), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n252), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n928), .B(new_n931), .C1(G143), .C2(new_n741), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n932), .B1(new_n371), .B2(new_n734), .C1(new_n274), .C2(new_n745), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n733), .A2(KEYINPUT46), .A3(G116), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT105), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n797), .A2(G107), .B1(new_n749), .B2(G283), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n934), .A2(KEYINPUT106), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(G317), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n937), .B1(new_n935), .B2(new_n936), .C1(new_n938), .C2(new_n722), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT46), .B1(new_n733), .B2(new_n433), .ZN(new_n940));
  INV_X1    g0740(.A(new_n454), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n726), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n741), .A2(G311), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n746), .A2(G303), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n942), .A2(new_n943), .A3(new_n363), .A4(new_n944), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n939), .A2(new_n940), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n226), .B2(new_n738), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n934), .A2(KEYINPUT106), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n933), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT47), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n716), .ZN(new_n951));
  INV_X1    g0751(.A(new_n771), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n775), .B1(new_n231), .B2(new_n351), .C1(new_n243), .C2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n951), .A2(new_n777), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n923), .B1(new_n924), .B2(new_n954), .ZN(G387));
  NOR2_X1   g0755(.A1(new_n734), .A2(new_n454), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n726), .A2(G311), .B1(G303), .B2(new_n749), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n938), .B2(new_n745), .ZN(new_n958));
  XNOR2_X1  g0758(.A(KEYINPUT108), .B(G322), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n741), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT48), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n956), .B(new_n961), .C1(G283), .C2(new_n797), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(KEYINPUT49), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n962), .A2(KEYINPUT49), .B1(new_n433), .B2(new_n739), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n723), .A2(new_n742), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n963), .A2(new_n964), .A3(new_n363), .A4(new_n965), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n803), .A2(new_n755), .B1(new_n220), .B2(new_n748), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n734), .A2(new_n224), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(new_n350), .C2(new_n797), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n738), .A2(new_n226), .B1(new_n214), .B2(new_n745), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n363), .B(new_n970), .C1(new_n277), .C2(new_n726), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n969), .B(new_n971), .C1(new_n274), .C2(new_n722), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n717), .B1(new_n966), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n662), .A2(new_n768), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n240), .A2(G45), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n231), .A2(new_n252), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n975), .A2(new_n952), .B1(new_n674), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n277), .A2(new_n214), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT50), .Z(new_n979));
  NAND2_X1  g0779(.A1(G68), .A2(G77), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n979), .A2(new_n461), .A3(new_n980), .A4(new_n674), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n977), .A2(new_n981), .B1(new_n435), .B2(new_n671), .ZN(new_n982));
  INV_X1    g0782(.A(new_n775), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n777), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n973), .A2(new_n974), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n912), .B2(new_n922), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n672), .B1(new_n707), .B2(new_n912), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n986), .B1(new_n913), .B2(new_n987), .ZN(G393));
  XNOR2_X1  g0788(.A(new_n919), .B(new_n669), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n920), .B(new_n672), .C1(new_n913), .C2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n922), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n734), .A2(new_n220), .B1(new_n722), .B2(new_n794), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT109), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n363), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n993), .B2(new_n992), .C1(new_n599), .C2(new_n738), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT110), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n741), .A2(G150), .B1(G159), .B2(new_n746), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT51), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n797), .A2(G77), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n749), .A2(new_n277), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G50), .B2(new_n726), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n741), .A2(G317), .B1(G311), .B2(new_n746), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT52), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G303), .B2(new_n726), .ZN(new_n1006));
  INV_X1    g0806(.A(G294), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n363), .B1(new_n748), .B2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1008), .B(new_n761), .C1(new_n723), .C2(new_n959), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1006), .B(new_n1009), .C1(new_n539), .C2(new_n736), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G283), .B2(new_n733), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n716), .B1(new_n1003), .B2(new_n1011), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n775), .B1(new_n226), .B2(new_n231), .C1(new_n952), .C2(new_n250), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n906), .A2(new_n768), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1012), .A2(new_n777), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n990), .A2(new_n991), .A3(new_n1015), .ZN(G390));
  NAND3_X1  g0816(.A1(new_n863), .A2(G330), .A3(new_n865), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AND3_X1   g0818(.A1(new_n843), .A2(KEYINPUT101), .A3(new_n784), .ZN(new_n1019));
  AOI21_X1  g0819(.A(KEYINPUT101), .B1(new_n843), .B2(new_n784), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n853), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n841), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n840), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n682), .A2(new_n660), .A3(new_n783), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n784), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n835), .B(new_n841), .C1(new_n1025), .C2(new_n853), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1018), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n706), .A2(new_n853), .A3(G330), .A4(new_n786), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1025), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n853), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n864), .B(new_n1022), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n841), .B1(new_n848), .B2(new_n853), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1028), .B(new_n1031), .C1(new_n1032), .C2(new_n840), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1027), .A2(new_n1033), .A3(KEYINPUT111), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT111), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n1018), .C1(new_n1023), .C2(new_n1026), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n706), .A2(G330), .A3(new_n786), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n1030), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1038), .B1(new_n1040), .B2(new_n1017), .ZN(new_n1041));
  OAI211_X1 g0841(.A(G330), .B(new_n786), .C1(new_n858), .C2(new_n862), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n1030), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1028), .A2(new_n1029), .A3(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n856), .B(new_n879), .C1(new_n1041), .C2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1037), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1034), .A2(new_n1045), .A3(new_n1036), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n672), .A3(new_n1048), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n840), .A2(new_n766), .ZN(new_n1050));
  INV_X1    g0850(.A(G125), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n722), .A2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(KEYINPUT54), .B(G143), .Z(new_n1053));
  AOI22_X1  g0853(.A1(new_n797), .A2(G159), .B1(new_n749), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(G137), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n758), .B2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT112), .Z(new_n1057));
  NAND2_X1  g0857(.A1(new_n733), .A2(G150), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT53), .Z(new_n1059));
  OAI21_X1  g0859(.A(new_n252), .B1(new_n738), .B2(new_n214), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT113), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1060), .A2(KEYINPUT113), .B1(G132), .B2(new_n746), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1057), .A2(new_n1059), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1052), .B(new_n1063), .C1(G128), .C2(new_n741), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n363), .B1(new_n758), .B2(new_n435), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n723), .A2(G294), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n739), .A2(G68), .B1(G283), .B2(new_n741), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n733), .A2(G87), .B1(G97), .B2(new_n749), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1000), .A4(new_n1068), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1065), .B(new_n1069), .C1(G116), .C2(new_n746), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT114), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n716), .B1(new_n1064), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n713), .B1(new_n278), .B2(new_n810), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1050), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1037), .B2(new_n922), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(KEYINPUT115), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT115), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1077), .B(new_n1074), .C1(new_n1037), .C2(new_n922), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1049), .B1(new_n1076), .B2(new_n1078), .ZN(G378));
  INV_X1    g0879(.A(KEYINPUT118), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n878), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n871), .A2(new_n873), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1082), .A2(KEYINPUT118), .A3(G330), .A4(new_n866), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n301), .A2(new_n304), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1085));
  XNOR2_X1  g0885(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n293), .A2(new_n655), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1086), .B(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1081), .A2(new_n1083), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1087), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1086), .B(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n874), .A2(new_n1091), .A3(KEYINPUT118), .A4(G330), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n1089), .A2(new_n855), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n855), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g0894(.A(KEYINPUT119), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1089), .A2(new_n855), .A3(new_n1092), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT119), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n922), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1045), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n856), .A2(new_n879), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT57), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n672), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1100), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1099), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n351), .A2(new_n748), .ZN(new_n1108));
  AOI21_X1  g0908(.A(G41), .B1(new_n723), .B2(G283), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1109), .B1(new_n435), .B2(new_n745), .C1(new_n216), .C2(new_n803), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1108), .B(new_n1110), .C1(G97), .C2(new_n726), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n252), .B(new_n968), .C1(G58), .C2(new_n739), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n926), .A3(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT58), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n214), .B1(new_n361), .B2(G41), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n803), .A2(new_n1051), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n733), .A2(new_n1053), .B1(G128), .B2(new_n746), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT116), .Z(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n1055), .B2(new_n748), .C1(new_n274), .C2(new_n736), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1116), .B(new_n1119), .C1(G132), .C2(new_n726), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT59), .ZN(new_n1121));
  AOI21_X1  g0921(.A(G33), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(G41), .B1(new_n723), .B2(G124), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(new_n755), .C2(new_n738), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1114), .B(new_n1115), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT117), .Z(new_n1127));
  NOR2_X1   g0927(.A1(new_n1127), .A2(new_n717), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1088), .A2(new_n766), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n810), .A2(new_n214), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NOR4_X1   g0931(.A1(new_n1128), .A2(new_n1129), .A3(new_n713), .A4(new_n1131), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1093), .A2(new_n1094), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n673), .A2(new_n1104), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1107), .A2(new_n1135), .ZN(G375));
  OR2_X1    g0936(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1030), .A2(new_n765), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n738), .A2(new_n371), .B1(new_n274), .B2(new_n748), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n734), .A2(new_n755), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(G128), .C2(new_n723), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n797), .A2(G50), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n741), .A2(G132), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n745), .A2(new_n1055), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n363), .B(new_n1144), .C1(new_n726), .C2(new_n1053), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n722), .A2(new_n729), .B1(new_n803), .B2(new_n1007), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n252), .B(new_n1147), .C1(G283), .C2(new_n746), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n733), .A2(G97), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n726), .A2(new_n433), .B1(G107), .B2(new_n749), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT120), .Z(new_n1151));
  AOI22_X1  g0951(.A1(new_n739), .A2(G77), .B1(new_n350), .B2(new_n797), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1148), .A2(new_n1149), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n717), .B1(new_n1146), .B2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n713), .B(new_n1154), .C1(new_n220), .C2(new_n810), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT121), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1137), .A2(new_n922), .B1(new_n1138), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n690), .A2(new_n427), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1158), .A2(new_n629), .A3(new_n879), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n909), .B1(new_n1137), .B2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1157), .B1(new_n1160), .B2(new_n1046), .ZN(G381));
  NOR2_X1   g0961(.A1(G387), .A2(G390), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OR2_X1    g0963(.A1(G381), .A2(G384), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1163), .A2(G396), .A3(G393), .A4(new_n1164), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1049), .A2(new_n1075), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1107), .A2(new_n1135), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(G407));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n1165), .B2(new_n656), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(G213), .ZN(G409));
  NAND2_X1  g0970(.A1(new_n656), .A2(G213), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1107), .A2(G378), .A3(new_n1135), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n909), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n922), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1132), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1166), .B(KEYINPUT122), .C1(new_n1174), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1172), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n910), .B1(new_n1047), .B2(new_n1159), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n855), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1097), .B1(new_n1183), .B2(new_n1096), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1098), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1180), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1096), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1132), .B1(new_n1187), .B2(new_n922), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT122), .B1(new_n1189), .B2(new_n1166), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1171), .B1(new_n1179), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n656), .A2(G213), .A3(G2897), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1137), .A2(new_n1159), .ZN(new_n1194));
  OAI211_X1 g0994(.A(KEYINPUT123), .B(new_n1045), .C1(new_n1194), .C2(KEYINPUT60), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT123), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1197));
  AOI21_X1  g0997(.A(KEYINPUT60), .B1(new_n1197), .B2(new_n1102), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1196), .B1(new_n1198), .B2(new_n1046), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1194), .A2(KEYINPUT60), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1195), .A2(new_n1199), .A3(new_n672), .A4(new_n1200), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1201), .A2(G384), .A3(new_n1157), .ZN(new_n1202));
  AOI21_X1  g1002(.A(G384), .B1(new_n1201), .B2(new_n1157), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1193), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1157), .ZN(new_n1205));
  INV_X1    g1005(.A(G384), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1201), .A2(G384), .A3(new_n1157), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n1208), .A3(new_n1192), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1204), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1191), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT61), .B1(new_n1212), .B2(KEYINPUT124), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(G393), .B(G396), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G387), .A2(G390), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1215), .B1(new_n1217), .B2(new_n1162), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1163), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1166), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT122), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(new_n1178), .A3(new_n1172), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1210), .B1(new_n1224), .B2(new_n1171), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT124), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1220), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1171), .B(new_n1228), .C1(new_n1179), .C2(new_n1190), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(KEYINPUT63), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT63), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1224), .A2(new_n1231), .A3(new_n1171), .A4(new_n1228), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1213), .A2(new_n1227), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT125), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT125), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1213), .A2(new_n1227), .A3(new_n1233), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT126), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1220), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1218), .A2(new_n1219), .A3(KEYINPUT126), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1229), .A2(KEYINPUT62), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1229), .A2(KEYINPUT62), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1242), .B1(new_n1246), .B2(new_n1225), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1238), .A2(new_n1247), .ZN(G405));
  NAND2_X1  g1048(.A1(G375), .A2(new_n1166), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1242), .A2(new_n1249), .A3(new_n1172), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1172), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1240), .A2(new_n1241), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1228), .A2(KEYINPUT127), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1250), .A2(KEYINPUT127), .A3(new_n1228), .A4(new_n1252), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(G402));
endmodule


