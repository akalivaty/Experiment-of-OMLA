

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728;

  XNOR2_X1 U371 ( .A(n361), .B(G107), .ZN(n464) );
  INV_X1 U372 ( .A(G122), .ZN(n361) );
  XNOR2_X1 U373 ( .A(n703), .B(n407), .ZN(n667) );
  INV_X1 U374 ( .A(G953), .ZN(n717) );
  XNOR2_X2 U375 ( .A(n468), .B(KEYINPUT22), .ZN(n505) );
  XNOR2_X2 U376 ( .A(n710), .B(G146), .ZN(n482) );
  XNOR2_X2 U377 ( .A(n477), .B(n476), .ZN(n710) );
  XNOR2_X2 U378 ( .A(n479), .B(G469), .ZN(n563) );
  XNOR2_X2 U379 ( .A(n502), .B(KEYINPUT100), .ZN(n724) );
  AND2_X2 U380 ( .A1(n501), .A2(n553), .ZN(n502) );
  XNOR2_X1 U381 ( .A(n385), .B(n384), .ZN(n624) );
  NAND2_X1 U382 ( .A1(n517), .A2(n554), .ZN(n385) );
  INV_X1 U383 ( .A(G125), .ZN(n398) );
  INV_X1 U384 ( .A(G143), .ZN(n377) );
  XNOR2_X1 U385 ( .A(n381), .B(n380), .ZN(n531) );
  NOR2_X1 U386 ( .A1(n392), .A2(n390), .ZN(n389) );
  AND2_X1 U387 ( .A1(n578), .A2(n577), .ZN(n414) );
  XNOR2_X1 U388 ( .A(n373), .B(KEYINPUT77), .ZN(n651) );
  INV_X1 U389 ( .A(n350), .ZN(n518) );
  NOR2_X1 U390 ( .A1(n565), .A2(n564), .ZN(n575) );
  XNOR2_X1 U391 ( .A(n434), .B(KEYINPUT19), .ZN(n574) );
  XNOR2_X1 U392 ( .A(n375), .B(KEYINPUT98), .ZN(n374) );
  AND2_X1 U393 ( .A1(n547), .A2(n546), .ZN(n569) );
  NOR2_X1 U394 ( .A1(n595), .A2(n551), .ZN(n375) );
  XNOR2_X1 U395 ( .A(n605), .B(n503), .ZN(n554) );
  XNOR2_X1 U396 ( .A(n431), .B(n430), .ZN(n535) );
  XNOR2_X1 U397 ( .A(n500), .B(n499), .ZN(n602) );
  XNOR2_X1 U398 ( .A(n378), .B(G478), .ZN(n523) );
  OR2_X1 U399 ( .A1(n688), .A2(G902), .ZN(n378) );
  XNOR2_X1 U400 ( .A(n369), .B(n495), .ZN(n690) );
  XNOR2_X1 U401 ( .A(n379), .B(n465), .ZN(n688) );
  XNOR2_X1 U402 ( .A(n356), .B(n352), .ZN(n477) );
  XNOR2_X1 U403 ( .A(n475), .B(KEYINPUT4), .ZN(n356) );
  XNOR2_X1 U404 ( .A(n377), .B(G128), .ZN(n463) );
  XNOR2_X1 U405 ( .A(n398), .B(G146), .ZN(n446) );
  XNOR2_X2 U406 ( .A(n441), .B(n351), .ZN(n350) );
  XOR2_X1 U407 ( .A(n440), .B(KEYINPUT0), .Z(n351) );
  NAND2_X1 U408 ( .A1(n421), .A2(n420), .ZN(n480) );
  INV_X2 U409 ( .A(n664), .ZN(n665) );
  XNOR2_X1 U410 ( .A(n423), .B(n452), .ZN(n411) );
  INV_X1 U411 ( .A(KEYINPUT71), .ZN(n419) );
  XNOR2_X1 U412 ( .A(n429), .B(KEYINPUT78), .ZN(n430) );
  NOR2_X1 U413 ( .A1(G953), .A2(G237), .ZN(n483) );
  NOR2_X1 U414 ( .A1(n662), .A2(n579), .ZN(n586) );
  XNOR2_X1 U415 ( .A(n389), .B(n399), .ZN(n579) );
  INV_X1 U416 ( .A(KEYINPUT48), .ZN(n399) );
  XNOR2_X1 U417 ( .A(n368), .B(KEYINPUT70), .ZN(n562) );
  NAND2_X1 U418 ( .A1(n553), .A2(n552), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n563), .B(KEYINPUT1), .ZN(n607) );
  XNOR2_X1 U420 ( .A(n422), .B(n464), .ZN(n423) );
  XNOR2_X1 U421 ( .A(n660), .B(n391), .ZN(n390) );
  INV_X1 U422 ( .A(KEYINPUT82), .ZN(n391) );
  XNOR2_X1 U423 ( .A(n484), .B(G113), .ZN(n388) );
  NAND2_X1 U424 ( .A1(G234), .A2(G237), .ZN(n435) );
  NAND2_X1 U425 ( .A1(n605), .A2(n593), .ZN(n536) );
  NOR2_X1 U426 ( .A1(n562), .A2(n561), .ZN(n367) );
  XNOR2_X1 U427 ( .A(G119), .B(G128), .ZN(n488) );
  XNOR2_X1 U428 ( .A(n446), .B(n397), .ZN(n709) );
  XNOR2_X1 U429 ( .A(G140), .B(KEYINPUT10), .ZN(n397) );
  XNOR2_X1 U430 ( .A(G116), .B(KEYINPUT7), .ZN(n460) );
  XOR2_X1 U431 ( .A(KEYINPUT9), .B(KEYINPUT96), .Z(n461) );
  XNOR2_X1 U432 ( .A(n463), .B(n376), .ZN(n476) );
  INV_X1 U433 ( .A(G134), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n409), .B(n408), .ZN(n407) );
  XNOR2_X1 U435 ( .A(n427), .B(n472), .ZN(n408) );
  INV_X1 U436 ( .A(KEYINPUT33), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n548), .B(n401), .ZN(n558) );
  XNOR2_X1 U438 ( .A(n549), .B(KEYINPUT39), .ZN(n401) );
  INV_X1 U439 ( .A(KEYINPUT83), .ZN(n549) );
  NAND2_X1 U440 ( .A1(n650), .A2(n394), .ZN(n580) );
  AND2_X1 U441 ( .A1(n554), .A2(n395), .ZN(n394) );
  NOR2_X1 U442 ( .A1(n562), .A2(n396), .ZN(n395) );
  INV_X1 U443 ( .A(n593), .ZN(n396) );
  NOR2_X1 U444 ( .A1(n690), .A2(G902), .ZN(n500) );
  BUF_X1 U445 ( .A(n535), .Z(n585) );
  XNOR2_X1 U446 ( .A(n457), .B(n393), .ZN(n522) );
  XNOR2_X1 U447 ( .A(n456), .B(G475), .ZN(n393) );
  NOR2_X1 U448 ( .A1(n523), .A2(n522), .ZN(n557) );
  INV_X1 U449 ( .A(KEYINPUT44), .ZN(n508) );
  NAND2_X1 U450 ( .A1(n382), .A2(n530), .ZN(n381) );
  INV_X1 U451 ( .A(KEYINPUT84), .ZN(n380) );
  XNOR2_X1 U452 ( .A(G122), .B(G143), .ZN(n447) );
  XOR2_X1 U453 ( .A(KEYINPUT94), .B(KEYINPUT11), .Z(n450) );
  XNOR2_X1 U454 ( .A(G104), .B(G107), .ZN(n469) );
  XOR2_X1 U455 ( .A(G140), .B(G101), .Z(n470) );
  NAND2_X1 U456 ( .A1(n509), .A2(n522), .ZN(n595) );
  XNOR2_X1 U457 ( .A(n482), .B(n386), .ZN(n633) );
  XNOR2_X1 U458 ( .A(n480), .B(n387), .ZN(n386) );
  XNOR2_X1 U459 ( .A(n388), .B(n481), .ZN(n387) );
  NOR2_X1 U460 ( .A1(n588), .A2(n587), .ZN(n591) );
  XNOR2_X1 U461 ( .A(n363), .B(n362), .ZN(n616) );
  INV_X1 U462 ( .A(KEYINPUT41), .ZN(n362) );
  NOR2_X1 U463 ( .A1(n596), .A2(n595), .ZN(n363) );
  INV_X1 U464 ( .A(n550), .ZN(n544) );
  XNOR2_X1 U465 ( .A(n367), .B(n366), .ZN(n565) );
  INV_X1 U466 ( .A(KEYINPUT28), .ZN(n366) );
  INV_X1 U467 ( .A(KEYINPUT6), .ZN(n503) );
  XNOR2_X1 U468 ( .A(n370), .B(n494), .ZN(n369) );
  XNOR2_X1 U469 ( .A(n466), .B(n467), .ZN(n379) );
  XNOR2_X1 U470 ( .A(n667), .B(n412), .ZN(n668) );
  XNOR2_X1 U471 ( .A(n400), .B(n560), .ZN(n722) );
  NOR2_X1 U472 ( .A1(n580), .A2(n585), .ZN(n555) );
  XNOR2_X1 U473 ( .A(n557), .B(KEYINPUT101), .ZN(n653) );
  INV_X1 U474 ( .A(n695), .ZN(n358) );
  INV_X1 U475 ( .A(KEYINPUT53), .ZN(n404) );
  XNOR2_X1 U476 ( .A(G137), .B(KEYINPUT69), .ZN(n352) );
  XOR2_X1 U477 ( .A(G119), .B(KEYINPUT3), .Z(n353) );
  XOR2_X1 U478 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n354) );
  XNOR2_X1 U479 ( .A(n410), .B(n426), .ZN(n409) );
  NAND2_X1 U480 ( .A1(n355), .A2(n531), .ZN(n357) );
  NAND2_X1 U481 ( .A1(n515), .A2(n514), .ZN(n355) );
  NAND2_X1 U482 ( .A1(n728), .A2(n722), .ZN(n365) );
  XNOR2_X1 U483 ( .A(n365), .B(n354), .ZN(n364) );
  NAND2_X1 U484 ( .A1(n558), .A2(n557), .ZN(n400) );
  XNOR2_X2 U485 ( .A(n357), .B(n532), .ZN(n700) );
  AND2_X1 U486 ( .A1(n359), .A2(n358), .ZN(G54) );
  XNOR2_X1 U487 ( .A(n676), .B(n677), .ZN(n359) );
  NAND2_X1 U488 ( .A1(n360), .A2(n568), .ZN(n512) );
  XNOR2_X1 U489 ( .A(n510), .B(n511), .ZN(n360) );
  NAND2_X1 U490 ( .A1(n723), .A2(KEYINPUT44), .ZN(n382) );
  NAND2_X1 U491 ( .A1(n575), .A2(n616), .ZN(n566) );
  NAND2_X1 U492 ( .A1(n592), .A2(n593), .ZN(n596) );
  NAND2_X1 U493 ( .A1(n414), .A2(n364), .ZN(n392) );
  NAND2_X1 U494 ( .A1(n493), .A2(G221), .ZN(n370) );
  NAND2_X1 U495 ( .A1(n576), .A2(n371), .ZN(n577) );
  XNOR2_X1 U496 ( .A(n651), .B(n372), .ZN(n371) );
  INV_X1 U497 ( .A(KEYINPUT47), .ZN(n372) );
  NAND2_X1 U498 ( .A1(n575), .A2(n574), .ZN(n373) );
  NAND2_X1 U499 ( .A1(n350), .A2(n374), .ZN(n468) );
  XNOR2_X2 U500 ( .A(n512), .B(KEYINPUT35), .ZN(n723) );
  NAND2_X1 U501 ( .A1(n383), .A2(n350), .ZN(n510) );
  INV_X1 U502 ( .A(n624), .ZN(n383) );
  XNOR2_X1 U503 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X1 U504 ( .A1(n505), .A2(n581), .ZN(n527) );
  NAND2_X1 U505 ( .A1(n403), .A2(n402), .ZN(n487) );
  NOR2_X1 U506 ( .A1(n581), .A2(n605), .ZN(n402) );
  INV_X1 U507 ( .A(n505), .ZN(n403) );
  XNOR2_X1 U508 ( .A(n405), .B(n404), .ZN(G75) );
  NAND2_X1 U509 ( .A1(n406), .A2(n717), .ZN(n405) );
  XNOR2_X1 U510 ( .A(n629), .B(KEYINPUT117), .ZN(n406) );
  XNOR2_X1 U511 ( .A(n446), .B(n463), .ZN(n410) );
  XNOR2_X2 U512 ( .A(n411), .B(n480), .ZN(n703) );
  XNOR2_X1 U513 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n412) );
  XNOR2_X1 U514 ( .A(KEYINPUT59), .B(KEYINPUT85), .ZN(n413) );
  OR2_X1 U515 ( .A1(n625), .A2(n624), .ZN(n415) );
  INV_X1 U516 ( .A(KEYINPUT67), .ZN(n440) );
  AND2_X1 U517 ( .A1(n626), .A2(n415), .ZN(n627) );
  AND2_X1 U518 ( .A1(n545), .A2(n544), .ZN(n546) );
  INV_X1 U519 ( .A(KEYINPUT31), .ZN(n519) );
  XNOR2_X1 U520 ( .A(n680), .B(n413), .ZN(n681) );
  XNOR2_X1 U521 ( .A(n519), .B(KEYINPUT93), .ZN(n520) );
  XNOR2_X1 U522 ( .A(n521), .B(n520), .ZN(n655) );
  NOR2_X1 U523 ( .A1(G952), .A2(n717), .ZN(n695) );
  XNOR2_X1 U524 ( .A(G116), .B(G101), .ZN(n416) );
  XNOR2_X1 U525 ( .A(n353), .B(n416), .ZN(n418) );
  INV_X1 U526 ( .A(n418), .ZN(n417) );
  NAND2_X1 U527 ( .A1(n417), .A2(KEYINPUT71), .ZN(n421) );
  NAND2_X1 U528 ( .A1(n419), .A2(n418), .ZN(n420) );
  XOR2_X1 U529 ( .A(KEYINPUT16), .B(KEYINPUT74), .Z(n422) );
  XNOR2_X1 U530 ( .A(G113), .B(G104), .ZN(n452) );
  XOR2_X1 U531 ( .A(KEYINPUT72), .B(G110), .Z(n472) );
  XOR2_X1 U532 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n425) );
  XNOR2_X1 U533 ( .A(KEYINPUT4), .B(KEYINPUT86), .ZN(n424) );
  XNOR2_X1 U534 ( .A(n425), .B(n424), .ZN(n426) );
  NAND2_X1 U535 ( .A1(G224), .A2(n717), .ZN(n427) );
  XNOR2_X1 U536 ( .A(G902), .B(KEYINPUT15), .ZN(n630) );
  NAND2_X1 U537 ( .A1(n667), .A2(n630), .ZN(n431) );
  NOR2_X1 U538 ( .A1(G237), .A2(G902), .ZN(n428) );
  XNOR2_X1 U539 ( .A(n428), .B(KEYINPUT75), .ZN(n432) );
  NAND2_X1 U540 ( .A1(n432), .A2(G210), .ZN(n429) );
  INV_X1 U541 ( .A(n535), .ZN(n433) );
  NAND2_X1 U542 ( .A1(G214), .A2(n432), .ZN(n593) );
  NAND2_X1 U543 ( .A1(n433), .A2(n593), .ZN(n434) );
  XOR2_X1 U544 ( .A(KEYINPUT14), .B(n435), .Z(n622) );
  NAND2_X1 U545 ( .A1(G952), .A2(n717), .ZN(n541) );
  INV_X1 U546 ( .A(n541), .ZN(n437) );
  NAND2_X1 U547 ( .A1(G953), .A2(G902), .ZN(n538) );
  NOR2_X1 U548 ( .A1(G898), .A2(n538), .ZN(n436) );
  NOR2_X1 U549 ( .A1(n437), .A2(n436), .ZN(n438) );
  NOR2_X1 U550 ( .A1(n622), .A2(n438), .ZN(n439) );
  NAND2_X1 U551 ( .A1(n574), .A2(n439), .ZN(n441) );
  XOR2_X1 U552 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n443) );
  NAND2_X1 U553 ( .A1(G234), .A2(n630), .ZN(n442) );
  XNOR2_X1 U554 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U555 ( .A(KEYINPUT90), .B(n444), .ZN(n496) );
  NAND2_X1 U556 ( .A1(n496), .A2(G221), .ZN(n445) );
  XOR2_X1 U557 ( .A(KEYINPUT21), .B(n445), .Z(n601) );
  INV_X1 U558 ( .A(n601), .ZN(n551) );
  XOR2_X2 U559 ( .A(KEYINPUT68), .B(G131), .Z(n475) );
  XNOR2_X1 U560 ( .A(n475), .B(n447), .ZN(n448) );
  XNOR2_X1 U561 ( .A(n709), .B(n448), .ZN(n455) );
  NAND2_X1 U562 ( .A1(G214), .A2(n483), .ZN(n449) );
  XNOR2_X1 U563 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U564 ( .A(KEYINPUT12), .B(n451), .ZN(n453) );
  XNOR2_X1 U565 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U566 ( .A(n455), .B(n454), .ZN(n680) );
  NOR2_X1 U567 ( .A1(G902), .A2(n680), .ZN(n457) );
  XNOR2_X1 U568 ( .A(KEYINPUT95), .B(KEYINPUT13), .ZN(n456) );
  XOR2_X1 U569 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n459) );
  NAND2_X1 U570 ( .A1(G234), .A2(n717), .ZN(n458) );
  XNOR2_X1 U571 ( .A(n459), .B(n458), .ZN(n493) );
  NAND2_X1 U572 ( .A1(G217), .A2(n493), .ZN(n467) );
  XNOR2_X1 U573 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U574 ( .A(n462), .B(KEYINPUT97), .Z(n466) );
  XNOR2_X1 U575 ( .A(n464), .B(n476), .ZN(n465) );
  INV_X1 U576 ( .A(n523), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U578 ( .A(n472), .B(n471), .Z(n474) );
  NAND2_X1 U579 ( .A1(G227), .A2(n717), .ZN(n473) );
  XNOR2_X1 U580 ( .A(n474), .B(n473), .ZN(n478) );
  XNOR2_X1 U581 ( .A(n478), .B(n482), .ZN(n673) );
  NOR2_X1 U582 ( .A1(G902), .A2(n673), .ZN(n479) );
  INV_X1 U583 ( .A(n607), .ZN(n581) );
  XOR2_X1 U584 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n481) );
  NAND2_X1 U585 ( .A1(n483), .A2(G210), .ZN(n484) );
  NOR2_X1 U586 ( .A1(G902), .A2(n633), .ZN(n486) );
  XNOR2_X1 U587 ( .A(KEYINPUT73), .B(G472), .ZN(n485) );
  XNOR2_X2 U588 ( .A(n486), .B(n485), .ZN(n605) );
  INV_X1 U589 ( .A(n605), .ZN(n561) );
  XNOR2_X1 U590 ( .A(n487), .B(KEYINPUT65), .ZN(n501) );
  XOR2_X1 U591 ( .A(G137), .B(G110), .Z(n489) );
  XNOR2_X1 U592 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U593 ( .A(n709), .B(n490), .ZN(n495) );
  XNOR2_X1 U594 ( .A(KEYINPUT88), .B(KEYINPUT24), .ZN(n491) );
  XNOR2_X1 U595 ( .A(n491), .B(KEYINPUT87), .ZN(n492) );
  XOR2_X1 U596 ( .A(KEYINPUT23), .B(n492), .Z(n494) );
  XOR2_X1 U597 ( .A(KEYINPUT89), .B(KEYINPUT25), .Z(n498) );
  NAND2_X1 U598 ( .A1(G217), .A2(n496), .ZN(n497) );
  XNOR2_X1 U599 ( .A(n498), .B(n497), .ZN(n499) );
  NOR2_X1 U600 ( .A1(n554), .A2(n602), .ZN(n504) );
  NAND2_X1 U601 ( .A1(n504), .A2(n581), .ZN(n506) );
  NOR2_X1 U602 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U603 ( .A(n507), .B(KEYINPUT32), .ZN(n725) );
  NOR2_X2 U604 ( .A1(n724), .A2(n725), .ZN(n513) );
  XNOR2_X1 U605 ( .A(n513), .B(n508), .ZN(n515) );
  NOR2_X1 U606 ( .A1(n522), .A2(n509), .ZN(n568) );
  XOR2_X1 U607 ( .A(KEYINPUT34), .B(KEYINPUT76), .Z(n511) );
  NAND2_X1 U608 ( .A1(n602), .A2(n601), .ZN(n608) );
  NOR2_X1 U609 ( .A1(n607), .A2(n608), .ZN(n517) );
  NAND2_X1 U610 ( .A1(n513), .A2(n723), .ZN(n514) );
  NOR2_X1 U611 ( .A1(n563), .A2(n608), .ZN(n545) );
  NOR2_X1 U612 ( .A1(n605), .A2(n518), .ZN(n516) );
  NAND2_X1 U613 ( .A1(n545), .A2(n516), .ZN(n642) );
  NAND2_X1 U614 ( .A1(n605), .A2(n517), .ZN(n614) );
  NOR2_X1 U615 ( .A1(n518), .A2(n614), .ZN(n521) );
  NAND2_X1 U616 ( .A1(n642), .A2(n655), .ZN(n525) );
  NAND2_X1 U617 ( .A1(n523), .A2(n522), .ZN(n656) );
  INV_X1 U618 ( .A(n656), .ZN(n646) );
  NOR2_X1 U619 ( .A1(n557), .A2(n646), .ZN(n597) );
  INV_X1 U620 ( .A(n597), .ZN(n524) );
  NAND2_X1 U621 ( .A1(n525), .A2(n524), .ZN(n528) );
  INV_X1 U622 ( .A(n602), .ZN(n553) );
  NOR2_X1 U623 ( .A1(n554), .A2(n553), .ZN(n526) );
  NAND2_X1 U624 ( .A1(n527), .A2(n526), .ZN(n639) );
  NAND2_X1 U625 ( .A1(n528), .A2(n639), .ZN(n529) );
  XNOR2_X1 U626 ( .A(n529), .B(KEYINPUT99), .ZN(n530) );
  INV_X1 U627 ( .A(KEYINPUT45), .ZN(n532) );
  INV_X1 U628 ( .A(KEYINPUT2), .ZN(n533) );
  NAND2_X1 U629 ( .A1(n700), .A2(n533), .ZN(n534) );
  XNOR2_X1 U630 ( .A(n534), .B(KEYINPUT81), .ZN(n588) );
  XNOR2_X1 U631 ( .A(n585), .B(KEYINPUT38), .ZN(n592) );
  XOR2_X1 U632 ( .A(KEYINPUT104), .B(KEYINPUT30), .Z(n537) );
  XNOR2_X1 U633 ( .A(n537), .B(n536), .ZN(n547) );
  NOR2_X1 U634 ( .A1(n622), .A2(n538), .ZN(n539) );
  XOR2_X1 U635 ( .A(KEYINPUT102), .B(n539), .Z(n540) );
  NOR2_X1 U636 ( .A1(G900), .A2(n540), .ZN(n543) );
  NOR2_X1 U637 ( .A1(n622), .A2(n541), .ZN(n542) );
  NOR2_X1 U638 ( .A1(n543), .A2(n542), .ZN(n550) );
  NAND2_X1 U639 ( .A1(n592), .A2(n569), .ZN(n548) );
  AND2_X1 U640 ( .A1(n558), .A2(n646), .ZN(n662) );
  NOR2_X1 U641 ( .A1(n551), .A2(n550), .ZN(n552) );
  INV_X1 U642 ( .A(n653), .ZN(n650) );
  XNOR2_X1 U643 ( .A(n555), .B(KEYINPUT36), .ZN(n556) );
  NAND2_X1 U644 ( .A1(n556), .A2(n581), .ZN(n660) );
  XOR2_X1 U645 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n559) );
  XNOR2_X1 U646 ( .A(KEYINPUT107), .B(n559), .ZN(n560) );
  XOR2_X1 U647 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n567) );
  XNOR2_X1 U648 ( .A(n563), .B(KEYINPUT106), .ZN(n564) );
  XNOR2_X1 U649 ( .A(n567), .B(n566), .ZN(n728) );
  NAND2_X1 U650 ( .A1(n597), .A2(KEYINPUT47), .ZN(n572) );
  NAND2_X1 U651 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U652 ( .A1(n570), .A2(n585), .ZN(n571) );
  XNOR2_X1 U653 ( .A(n571), .B(KEYINPUT105), .ZN(n726) );
  NAND2_X1 U654 ( .A1(n572), .A2(n726), .ZN(n573) );
  XNOR2_X1 U655 ( .A(n573), .B(KEYINPUT79), .ZN(n578) );
  NAND2_X1 U656 ( .A1(n651), .A2(n597), .ZN(n576) );
  NOR2_X1 U657 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U658 ( .A(KEYINPUT43), .B(KEYINPUT103), .ZN(n582) );
  XNOR2_X1 U659 ( .A(n583), .B(n582), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n663) );
  NAND2_X1 U661 ( .A1(n586), .A2(n663), .ZN(n589) );
  INV_X1 U662 ( .A(n589), .ZN(n715) );
  NOR2_X1 U663 ( .A1(n715), .A2(KEYINPUT2), .ZN(n587) );
  NOR2_X2 U664 ( .A1(n589), .A2(n700), .ZN(n631) );
  NAND2_X1 U665 ( .A1(n631), .A2(KEYINPUT2), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n628) );
  NOR2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U668 ( .A1(n595), .A2(n594), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n624), .A2(n600), .ZN(n619) );
  NOR2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U673 ( .A(KEYINPUT49), .B(n603), .Z(n604) );
  NOR2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U675 ( .A(KEYINPUT115), .B(n606), .Z(n612) );
  NAND2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U677 ( .A(n609), .B(KEYINPUT116), .ZN(n610) );
  XNOR2_X1 U678 ( .A(KEYINPUT50), .B(n610), .ZN(n611) );
  NAND2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U680 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U681 ( .A(KEYINPUT51), .B(n615), .ZN(n617) );
  INV_X1 U682 ( .A(n616), .ZN(n625) );
  NOR2_X1 U683 ( .A1(n617), .A2(n625), .ZN(n618) );
  NOR2_X1 U684 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U685 ( .A(n620), .B(KEYINPUT52), .ZN(n621) );
  NOR2_X1 U686 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U687 ( .A1(G952), .A2(n623), .ZN(n626) );
  NAND2_X1 U688 ( .A1(n628), .A2(n627), .ZN(n629) );
  INV_X1 U689 ( .A(n630), .ZN(n678) );
  AND2_X1 U690 ( .A1(n678), .A2(G472), .ZN(n632) );
  XNOR2_X1 U691 ( .A(n631), .B(KEYINPUT2), .ZN(n664) );
  NAND2_X1 U692 ( .A1(n632), .A2(n665), .ZN(n635) );
  XNOR2_X1 U693 ( .A(n633), .B(KEYINPUT62), .ZN(n634) );
  XNOR2_X1 U694 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X1 U695 ( .A1(n695), .A2(n636), .ZN(n638) );
  INV_X1 U696 ( .A(KEYINPUT63), .ZN(n637) );
  XNOR2_X1 U697 ( .A(n638), .B(n637), .ZN(G57) );
  XNOR2_X1 U698 ( .A(G101), .B(KEYINPUT110), .ZN(n640) );
  XNOR2_X1 U699 ( .A(n640), .B(n639), .ZN(G3) );
  NOR2_X1 U700 ( .A1(n653), .A2(n642), .ZN(n641) );
  XOR2_X1 U701 ( .A(G104), .B(n641), .Z(G6) );
  NOR2_X1 U702 ( .A1(n656), .A2(n642), .ZN(n644) );
  XNOR2_X1 U703 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n643) );
  XNOR2_X1 U704 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U705 ( .A(G107), .B(n645), .ZN(G9) );
  XOR2_X1 U706 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n648) );
  NAND2_X1 U707 ( .A1(n651), .A2(n646), .ZN(n647) );
  XNOR2_X1 U708 ( .A(n648), .B(n647), .ZN(n649) );
  XOR2_X1 U709 ( .A(G128), .B(n649), .Z(G30) );
  NAND2_X1 U710 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U711 ( .A(n652), .B(G146), .ZN(G48) );
  NOR2_X1 U712 ( .A1(n653), .A2(n655), .ZN(n654) );
  XOR2_X1 U713 ( .A(G113), .B(n654), .Z(G15) );
  NOR2_X1 U714 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U715 ( .A(G116), .B(n657), .Z(G18) );
  XOR2_X1 U716 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n659) );
  XNOR2_X1 U717 ( .A(G125), .B(KEYINPUT37), .ZN(n658) );
  XNOR2_X1 U718 ( .A(n659), .B(n658), .ZN(n661) );
  XOR2_X1 U719 ( .A(n661), .B(n660), .Z(G27) );
  XOR2_X1 U720 ( .A(G134), .B(n662), .Z(G36) );
  XNOR2_X1 U721 ( .A(G140), .B(n663), .ZN(G42) );
  AND2_X1 U722 ( .A1(n678), .A2(G210), .ZN(n666) );
  NAND2_X1 U723 ( .A1(n666), .A2(n665), .ZN(n669) );
  NOR2_X1 U724 ( .A1(n695), .A2(n670), .ZN(n672) );
  XNOR2_X1 U725 ( .A(KEYINPUT56), .B(KEYINPUT118), .ZN(n671) );
  XNOR2_X1 U726 ( .A(n672), .B(n671), .ZN(G51) );
  XOR2_X1 U727 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n675) );
  XNOR2_X1 U728 ( .A(n673), .B(KEYINPUT119), .ZN(n674) );
  XNOR2_X1 U729 ( .A(n675), .B(n674), .ZN(n677) );
  AND2_X2 U730 ( .A1(n678), .A2(n665), .ZN(n691) );
  NAND2_X1 U731 ( .A1(n691), .A2(G469), .ZN(n676) );
  AND2_X1 U732 ( .A1(n678), .A2(G475), .ZN(n679) );
  NAND2_X1 U733 ( .A1(n679), .A2(n665), .ZN(n682) );
  XNOR2_X1 U734 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U735 ( .A1(n695), .A2(n683), .ZN(n686) );
  XNOR2_X1 U736 ( .A(KEYINPUT120), .B(KEYINPUT60), .ZN(n684) );
  XNOR2_X1 U737 ( .A(n684), .B(KEYINPUT66), .ZN(n685) );
  XNOR2_X1 U738 ( .A(n686), .B(n685), .ZN(G60) );
  NAND2_X1 U739 ( .A1(G478), .A2(n691), .ZN(n687) );
  XNOR2_X1 U740 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X1 U741 ( .A1(n695), .A2(n689), .ZN(G63) );
  XOR2_X1 U742 ( .A(n690), .B(KEYINPUT121), .Z(n693) );
  NAND2_X1 U743 ( .A1(n691), .A2(G217), .ZN(n692) );
  XNOR2_X1 U744 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U745 ( .A1(n695), .A2(n694), .ZN(G66) );
  NAND2_X1 U746 ( .A1(G224), .A2(G953), .ZN(n696) );
  XNOR2_X1 U747 ( .A(n696), .B(KEYINPUT61), .ZN(n697) );
  XNOR2_X1 U748 ( .A(KEYINPUT122), .B(n697), .ZN(n698) );
  NAND2_X1 U749 ( .A1(n698), .A2(G898), .ZN(n699) );
  XNOR2_X1 U750 ( .A(n699), .B(KEYINPUT123), .ZN(n702) );
  NOR2_X1 U751 ( .A1(n700), .A2(G953), .ZN(n701) );
  NOR2_X1 U752 ( .A1(n702), .A2(n701), .ZN(n708) );
  NOR2_X1 U753 ( .A1(G898), .A2(n717), .ZN(n705) );
  XOR2_X1 U754 ( .A(n703), .B(G110), .Z(n704) );
  NOR2_X1 U755 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U756 ( .A(KEYINPUT124), .B(n706), .Z(n707) );
  XNOR2_X1 U757 ( .A(n708), .B(n707), .ZN(G69) );
  XOR2_X1 U758 ( .A(n710), .B(n709), .Z(n711) );
  XOR2_X1 U759 ( .A(KEYINPUT125), .B(n711), .Z(n716) );
  XOR2_X1 U760 ( .A(KEYINPUT126), .B(n716), .Z(n712) );
  XNOR2_X1 U761 ( .A(G227), .B(n712), .ZN(n713) );
  NAND2_X1 U762 ( .A1(n713), .A2(G900), .ZN(n714) );
  NAND2_X1 U763 ( .A1(n714), .A2(G953), .ZN(n720) );
  XNOR2_X1 U764 ( .A(n716), .B(n715), .ZN(n718) );
  NAND2_X1 U765 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U766 ( .A1(n720), .A2(n719), .ZN(G72) );
  XOR2_X1 U767 ( .A(G131), .B(KEYINPUT127), .Z(n721) );
  XNOR2_X1 U768 ( .A(n722), .B(n721), .ZN(G33) );
  XOR2_X1 U769 ( .A(G122), .B(n723), .Z(G24) );
  XOR2_X1 U770 ( .A(G110), .B(n724), .Z(G12) );
  XOR2_X1 U771 ( .A(G119), .B(n725), .Z(G21) );
  XNOR2_X1 U772 ( .A(G143), .B(KEYINPUT112), .ZN(n727) );
  XNOR2_X1 U773 ( .A(n727), .B(n726), .ZN(G45) );
  XNOR2_X1 U774 ( .A(G137), .B(n728), .ZN(G39) );
endmodule

