

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737;

  XNOR2_X1 U380 ( .A(n669), .B(KEYINPUT6), .ZN(n557) );
  INV_X1 U381 ( .A(G953), .ZN(n716) );
  XOR2_X1 U382 ( .A(n363), .B(n423), .Z(n358) );
  XNOR2_X2 U383 ( .A(n398), .B(KEYINPUT0), .ZN(n520) );
  NOR2_X2 U384 ( .A1(n569), .A2(n441), .ZN(n398) );
  XNOR2_X1 U385 ( .A(n448), .B(n416), .ZN(n712) );
  NOR2_X2 U386 ( .A1(n557), .A2(n536), .ZN(n480) );
  XNOR2_X2 U387 ( .A(n454), .B(n453), .ZN(n669) );
  XNOR2_X2 U388 ( .A(n474), .B(n403), .ZN(n723) );
  XNOR2_X2 U389 ( .A(n385), .B(n449), .ZN(n474) );
  NOR2_X1 U390 ( .A1(n698), .A2(G902), .ZN(n478) );
  NOR2_X1 U391 ( .A1(n614), .A2(n706), .ZN(n616) );
  NOR2_X1 U392 ( .A1(n610), .A2(n706), .ZN(n612) );
  NOR2_X1 U393 ( .A1(n696), .A2(n706), .ZN(n697) );
  NAND2_X1 U394 ( .A1(n361), .A2(n359), .ZN(n374) );
  OR2_X1 U395 ( .A1(n414), .A2(KEYINPUT32), .ZN(n412) );
  XNOR2_X1 U396 ( .A(n472), .B(n381), .ZN(n665) );
  XNOR2_X1 U397 ( .A(n400), .B(n713), .ZN(n475) );
  XNOR2_X1 U398 ( .A(n425), .B(n417), .ZN(n448) );
  XNOR2_X1 U399 ( .A(n418), .B(G119), .ZN(n417) );
  XNOR2_X1 U400 ( .A(n444), .B(n430), .ZN(n400) );
  XNOR2_X1 U401 ( .A(n426), .B(G122), .ZN(n416) );
  XNOR2_X1 U402 ( .A(G131), .B(G134), .ZN(n449) );
  XNOR2_X1 U403 ( .A(n429), .B(G107), .ZN(n713) );
  XNOR2_X1 U404 ( .A(G104), .B(G110), .ZN(n429) );
  XNOR2_X1 U405 ( .A(n473), .B(KEYINPUT88), .ZN(n403) );
  XOR2_X1 U406 ( .A(G137), .B(G140), .Z(n473) );
  XNOR2_X1 U407 ( .A(G146), .B(G125), .ZN(n459) );
  INV_X1 U408 ( .A(KEYINPUT3), .ZN(n418) );
  NOR2_X1 U409 ( .A1(n693), .A2(n600), .ZN(n433) );
  XNOR2_X1 U410 ( .A(n452), .B(KEYINPUT72), .ZN(n453) );
  INV_X1 U411 ( .A(G472), .ZN(n452) );
  XNOR2_X1 U412 ( .A(KEYINPUT10), .B(n459), .ZN(n722) );
  XOR2_X1 U413 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n430) );
  INV_X1 U414 ( .A(G469), .ZN(n477) );
  XNOR2_X1 U415 ( .A(G113), .B(G131), .ZN(n489) );
  NAND2_X1 U416 ( .A1(n386), .A2(n380), .ZN(n379) );
  AND2_X1 U417 ( .A1(n364), .A2(n387), .ZN(n386) );
  AND2_X1 U418 ( .A1(n599), .A2(n370), .ZN(n380) );
  OR2_X1 U419 ( .A1(n662), .A2(KEYINPUT84), .ZN(n387) );
  NOR2_X1 U420 ( .A1(n530), .A2(n528), .ZN(n529) );
  XNOR2_X1 U421 ( .A(n428), .B(n427), .ZN(n498) );
  XNOR2_X1 U422 ( .A(G143), .B(G128), .ZN(n428) );
  XNOR2_X1 U423 ( .A(n677), .B(KEYINPUT117), .ZN(n408) );
  XNOR2_X1 U424 ( .A(n401), .B(KEYINPUT51), .ZN(n675) );
  XNOR2_X1 U425 ( .A(G119), .B(G110), .ZN(n460) );
  XNOR2_X1 U426 ( .A(n488), .B(n376), .ZN(n613) );
  XNOR2_X1 U427 ( .A(n495), .B(n487), .ZN(n376) );
  XNOR2_X1 U428 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n423) );
  XNOR2_X1 U429 ( .A(n498), .B(KEYINPUT4), .ZN(n385) );
  XOR2_X1 U430 ( .A(KEYINPUT74), .B(KEYINPUT16), .Z(n426) );
  XNOR2_X1 U431 ( .A(n409), .B(n435), .ZN(n586) );
  NOR2_X1 U432 ( .A1(n527), .A2(n415), .ZN(n414) );
  INV_X1 U433 ( .A(n557), .ZN(n415) );
  XNOR2_X1 U434 ( .A(n586), .B(KEYINPUT19), .ZN(n569) );
  XNOR2_X1 U435 ( .A(n567), .B(n568), .ZN(n384) );
  NOR2_X1 U436 ( .A1(n704), .A2(G902), .ZN(n381) );
  XNOR2_X1 U437 ( .A(KEYINPUT22), .B(KEYINPUT73), .ZN(n521) );
  NAND2_X1 U438 ( .A1(n699), .A2(G475), .ZN(n397) );
  XNOR2_X1 U439 ( .A(n404), .B(n723), .ZN(n698) );
  XNOR2_X1 U440 ( .A(n476), .B(G146), .ZN(n404) );
  XNOR2_X1 U441 ( .A(n475), .B(n421), .ZN(n476) );
  NOR2_X1 U442 ( .A1(G952), .A2(n716), .ZN(n706) );
  INV_X1 U443 ( .A(KEYINPUT84), .ZN(n390) );
  XOR2_X1 U444 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n484) );
  XNOR2_X1 U445 ( .A(KEYINPUT94), .B(KEYINPUT96), .ZN(n483) );
  XNOR2_X1 U446 ( .A(G143), .B(G140), .ZN(n491) );
  AND2_X1 U447 ( .A1(n377), .A2(n369), .ZN(n727) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n377) );
  INV_X1 U449 ( .A(KEYINPUT48), .ZN(n378) );
  XNOR2_X1 U450 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n545) );
  XOR2_X1 U451 ( .A(G122), .B(G107), .Z(n500) );
  XNOR2_X1 U452 ( .A(n407), .B(n405), .ZN(n678) );
  XNOR2_X1 U453 ( .A(n406), .B(KEYINPUT120), .ZN(n405) );
  NAND2_X1 U454 ( .A1(n408), .A2(n362), .ZN(n407) );
  INV_X1 U455 ( .A(KEYINPUT52), .ZN(n406) );
  XNOR2_X1 U456 ( .A(n556), .B(n555), .ZN(n596) );
  XNOR2_X1 U457 ( .A(n554), .B(KEYINPUT39), .ZN(n555) );
  NOR2_X1 U458 ( .A1(n565), .A2(n396), .ZN(n585) );
  OR2_X1 U459 ( .A1(n557), .A2(n636), .ZN(n396) );
  NOR2_X1 U460 ( .A1(n536), .A2(n566), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n497), .B(n496), .ZN(n538) );
  INV_X1 U462 ( .A(n669), .ZN(n566) );
  XNOR2_X1 U463 ( .A(n467), .B(n382), .ZN(n704) );
  XNOR2_X1 U464 ( .A(n466), .B(n722), .ZN(n382) );
  XNOR2_X1 U465 ( .A(n712), .B(n375), .ZN(n431) );
  XNOR2_X1 U466 ( .A(n424), .B(n358), .ZN(n375) );
  OR2_X1 U467 ( .A1(n525), .A2(KEYINPUT32), .ZN(n411) );
  NAND2_X1 U468 ( .A1(n384), .A2(n367), .ZN(n634) );
  INV_X1 U469 ( .A(n569), .ZN(n383) );
  INV_X1 U470 ( .A(n634), .ZN(n629) );
  XNOR2_X1 U471 ( .A(n397), .B(n372), .ZN(n614) );
  INV_X1 U472 ( .A(n706), .ZN(n392) );
  XNOR2_X1 U473 ( .A(n698), .B(n373), .ZN(n394) );
  NOR2_X1 U474 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U475 ( .A1(n544), .A2(n365), .ZN(n359) );
  NAND2_X1 U476 ( .A1(n557), .A2(KEYINPUT32), .ZN(n360) );
  NAND2_X2 U477 ( .A1(n606), .A2(n605), .ZN(n699) );
  AND2_X1 U478 ( .A1(n533), .A2(n532), .ZN(n361) );
  OR2_X1 U479 ( .A1(n661), .A2(n660), .ZN(n362) );
  XOR2_X1 U480 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n363) );
  AND2_X1 U481 ( .A1(n584), .A2(n583), .ZN(n364) );
  AND2_X1 U482 ( .A1(n543), .A2(n617), .ZN(n365) );
  AND2_X1 U483 ( .A1(n410), .A2(n412), .ZN(n366) );
  AND2_X1 U484 ( .A1(n383), .A2(n534), .ZN(n367) );
  XOR2_X1 U485 ( .A(n432), .B(KEYINPUT79), .Z(n368) );
  AND2_X1 U486 ( .A1(n645), .A2(n646), .ZN(n369) );
  AND2_X1 U487 ( .A1(n389), .A2(n388), .ZN(n370) );
  AND2_X1 U488 ( .A1(n662), .A2(KEYINPUT84), .ZN(n371) );
  XOR2_X1 U489 ( .A(n613), .B(KEYINPUT59), .Z(n372) );
  XNOR2_X1 U490 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n373) );
  XNOR2_X2 U491 ( .A(n374), .B(n545), .ZN(n707) );
  NAND2_X1 U492 ( .A1(n525), .A2(n413), .ZN(n410) );
  XNOR2_X2 U493 ( .A(n522), .B(n521), .ZN(n525) );
  INV_X1 U494 ( .A(n459), .ZN(n458) );
  XOR2_X2 U495 ( .A(KEYINPUT67), .B(G101), .Z(n444) );
  XNOR2_X1 U496 ( .A(n431), .B(n399), .ZN(n693) );
  NOR2_X1 U497 ( .A1(n653), .A2(n666), .ZN(n518) );
  XNOR2_X1 U498 ( .A(n517), .B(KEYINPUT99), .ZN(n653) );
  NAND2_X1 U499 ( .A1(n366), .A2(n411), .ZN(n735) );
  NAND2_X1 U500 ( .A1(n384), .A2(n534), .ZN(n594) );
  XNOR2_X1 U501 ( .A(n475), .B(n385), .ZN(n399) );
  NAND2_X1 U502 ( .A1(n590), .A2(n662), .ZN(n644) );
  NAND2_X1 U503 ( .A1(n590), .A2(n371), .ZN(n388) );
  NAND2_X1 U504 ( .A1(n391), .A2(n390), .ZN(n389) );
  INV_X1 U505 ( .A(n590), .ZN(n391) );
  AND2_X1 U506 ( .A1(n393), .A2(n392), .ZN(G54) );
  XNOR2_X1 U507 ( .A(n395), .B(n394), .ZN(n393) );
  NAND2_X1 U508 ( .A1(n699), .A2(G469), .ZN(n395) );
  INV_X1 U509 ( .A(n520), .ZN(n515) );
  NAND2_X1 U510 ( .A1(n673), .A2(n674), .ZN(n401) );
  XNOR2_X1 U511 ( .A(n402), .B(KEYINPUT93), .ZN(n674) );
  NAND2_X1 U512 ( .A1(n553), .A2(n650), .ZN(n409) );
  XNOR2_X1 U513 ( .A(n433), .B(n368), .ZN(n553) );
  NOR2_X1 U514 ( .A1(n527), .A2(n360), .ZN(n413) );
  NAND2_X1 U515 ( .A1(n525), .A2(n557), .ZN(n541) );
  NAND2_X1 U516 ( .A1(n727), .A2(n707), .ZN(n648) );
  XNOR2_X1 U517 ( .A(n609), .B(n608), .ZN(n610) );
  AND2_X1 U518 ( .A1(G224), .A2(n716), .ZN(n419) );
  XNOR2_X1 U519 ( .A(KEYINPUT62), .B(KEYINPUT108), .ZN(n420) );
  AND2_X1 U520 ( .A1(G227), .A2(n716), .ZN(n421) );
  AND2_X1 U521 ( .A1(n530), .A2(n528), .ZN(n422) );
  XNOR2_X1 U522 ( .A(G113), .B(G116), .ZN(n425) );
  XNOR2_X1 U523 ( .A(n458), .B(n419), .ZN(n424) );
  INV_X1 U524 ( .A(KEYINPUT64), .ZN(n427) );
  INV_X1 U525 ( .A(KEYINPUT85), .ZN(n554) );
  XNOR2_X1 U526 ( .A(n607), .B(n420), .ZN(n608) );
  XNOR2_X1 U527 ( .A(KEYINPUT36), .B(KEYINPUT107), .ZN(n588) );
  INV_X1 U528 ( .A(KEYINPUT63), .ZN(n611) );
  XNOR2_X1 U529 ( .A(KEYINPUT60), .B(KEYINPUT66), .ZN(n615) );
  INV_X1 U530 ( .A(KEYINPUT34), .ZN(n482) );
  XOR2_X1 U531 ( .A(KEYINPUT15), .B(G902), .Z(n600) );
  OR2_X1 U532 ( .A1(G237), .A2(G902), .ZN(n434) );
  NAND2_X1 U533 ( .A1(n434), .A2(G210), .ZN(n432) );
  NAND2_X1 U534 ( .A1(G214), .A2(n434), .ZN(n650) );
  INV_X1 U535 ( .A(KEYINPUT86), .ZN(n435) );
  NAND2_X1 U536 ( .A1(G234), .A2(G237), .ZN(n436) );
  XNOR2_X1 U537 ( .A(n436), .B(KEYINPUT14), .ZN(n649) );
  OR2_X1 U538 ( .A1(n716), .A2(G902), .ZN(n437) );
  NAND2_X1 U539 ( .A1(n649), .A2(n437), .ZN(n439) );
  NOR2_X1 U540 ( .A1(G953), .A2(G952), .ZN(n438) );
  NOR2_X1 U541 ( .A1(n439), .A2(n438), .ZN(n549) );
  NAND2_X1 U542 ( .A1(G953), .A2(G898), .ZN(n440) );
  NAND2_X1 U543 ( .A1(n549), .A2(n440), .ZN(n441) );
  XOR2_X1 U544 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n443) );
  NOR2_X1 U545 ( .A1(G953), .A2(G237), .ZN(n486) );
  NAND2_X1 U546 ( .A1(n486), .A2(G210), .ZN(n442) );
  XNOR2_X1 U547 ( .A(n443), .B(n442), .ZN(n447) );
  XNOR2_X1 U548 ( .A(n444), .B(G146), .ZN(n445) );
  XNOR2_X1 U549 ( .A(n445), .B(G137), .ZN(n446) );
  XOR2_X1 U550 ( .A(n447), .B(n446), .Z(n451) );
  XNOR2_X1 U551 ( .A(n448), .B(n474), .ZN(n450) );
  XNOR2_X1 U552 ( .A(n451), .B(n450), .ZN(n607) );
  NOR2_X1 U553 ( .A1(n607), .A2(G902), .ZN(n454) );
  XOR2_X1 U554 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n457) );
  INV_X1 U555 ( .A(n600), .ZN(n602) );
  NAND2_X1 U556 ( .A1(n602), .A2(G234), .ZN(n455) );
  XNOR2_X1 U557 ( .A(n455), .B(KEYINPUT20), .ZN(n468) );
  NAND2_X1 U558 ( .A1(G221), .A2(n468), .ZN(n456) );
  XNOR2_X1 U559 ( .A(n457), .B(n456), .ZN(n666) );
  XNOR2_X1 U560 ( .A(n460), .B(n473), .ZN(n464) );
  XOR2_X1 U561 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n462) );
  XNOR2_X1 U562 ( .A(G128), .B(KEYINPUT23), .ZN(n461) );
  XNOR2_X1 U563 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U564 ( .A(n464), .B(n463), .Z(n467) );
  NAND2_X1 U565 ( .A1(G234), .A2(n716), .ZN(n465) );
  XOR2_X1 U566 ( .A(KEYINPUT8), .B(n465), .Z(n503) );
  NAND2_X1 U567 ( .A1(G221), .A2(n503), .ZN(n466) );
  XOR2_X1 U568 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n470) );
  NAND2_X1 U569 ( .A1(G217), .A2(n468), .ZN(n469) );
  XNOR2_X1 U570 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U571 ( .A(KEYINPUT90), .B(n471), .ZN(n472) );
  NOR2_X1 U572 ( .A1(n666), .A2(n665), .ZN(n663) );
  XNOR2_X2 U573 ( .A(n478), .B(n477), .ZN(n534) );
  XNOR2_X2 U574 ( .A(n534), .B(KEYINPUT1), .ZN(n662) );
  NAND2_X1 U575 ( .A1(n663), .A2(n662), .ZN(n536) );
  XOR2_X1 U576 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n479) );
  XNOR2_X1 U577 ( .A(n480), .B(n479), .ZN(n661) );
  NOR2_X1 U578 ( .A1(n515), .A2(n661), .ZN(n481) );
  XNOR2_X1 U579 ( .A(n482), .B(n481), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U581 ( .A(n722), .B(n485), .Z(n488) );
  NAND2_X1 U582 ( .A1(G214), .A2(n486), .ZN(n487) );
  XOR2_X1 U583 ( .A(G122), .B(G104), .Z(n490) );
  XNOR2_X1 U584 ( .A(n490), .B(n489), .ZN(n494) );
  XOR2_X1 U585 ( .A(KEYINPUT95), .B(KEYINPUT11), .Z(n492) );
  XNOR2_X1 U586 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U587 ( .A(n494), .B(n493), .Z(n495) );
  NOR2_X1 U588 ( .A1(G902), .A2(n613), .ZN(n497) );
  XNOR2_X1 U589 ( .A(KEYINPUT13), .B(G475), .ZN(n496) );
  INV_X1 U590 ( .A(n498), .ZN(n502) );
  XNOR2_X1 U591 ( .A(G116), .B(G134), .ZN(n499) );
  XNOR2_X1 U592 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U593 ( .A(n502), .B(n501), .ZN(n507) );
  XOR2_X1 U594 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n505) );
  NAND2_X1 U595 ( .A1(G217), .A2(n503), .ZN(n504) );
  XNOR2_X1 U596 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U597 ( .A(n507), .B(n506), .ZN(n701) );
  NOR2_X1 U598 ( .A1(G902), .A2(n701), .ZN(n509) );
  XNOR2_X1 U599 ( .A(KEYINPUT98), .B(G478), .ZN(n508) );
  XNOR2_X1 U600 ( .A(n509), .B(n508), .ZN(n539) );
  INV_X1 U601 ( .A(n539), .ZN(n516) );
  NAND2_X1 U602 ( .A1(n538), .A2(n516), .ZN(n510) );
  XOR2_X1 U603 ( .A(KEYINPUT102), .B(n510), .Z(n574) );
  INV_X1 U604 ( .A(n574), .ZN(n511) );
  NOR2_X2 U605 ( .A1(n512), .A2(n511), .ZN(n514) );
  XNOR2_X1 U606 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n513) );
  XNOR2_X2 U607 ( .A(n514), .B(n513), .ZN(n734) );
  NAND2_X1 U608 ( .A1(KEYINPUT44), .A2(n734), .ZN(n544) );
  NOR2_X1 U609 ( .A1(n538), .A2(n516), .ZN(n517) );
  XNOR2_X1 U610 ( .A(KEYINPUT100), .B(n518), .ZN(n519) );
  NAND2_X1 U611 ( .A1(n520), .A2(n519), .ZN(n522) );
  INV_X1 U612 ( .A(n662), .ZN(n561) );
  NAND2_X1 U613 ( .A1(n525), .A2(n561), .ZN(n524) );
  NAND2_X1 U614 ( .A1(n665), .A2(n566), .ZN(n523) );
  NOR2_X1 U615 ( .A1(n524), .A2(n523), .ZN(n627) );
  NAND2_X1 U616 ( .A1(n665), .A2(n662), .ZN(n526) );
  XOR2_X1 U617 ( .A(KEYINPUT101), .B(n526), .Z(n527) );
  NOR2_X1 U618 ( .A1(n627), .A2(n735), .ZN(n530) );
  INV_X1 U619 ( .A(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U620 ( .A(n529), .B(KEYINPUT65), .ZN(n533) );
  INV_X1 U621 ( .A(n734), .ZN(n531) );
  NAND2_X1 U622 ( .A1(n422), .A2(n531), .ZN(n532) );
  NAND2_X1 U623 ( .A1(n663), .A2(n534), .ZN(n550) );
  NOR2_X1 U624 ( .A1(n515), .A2(n550), .ZN(n535) );
  NAND2_X1 U625 ( .A1(n566), .A2(n535), .ZN(n622) );
  NOR2_X1 U626 ( .A1(n674), .A2(n515), .ZN(n537) );
  XNOR2_X1 U627 ( .A(n537), .B(KEYINPUT31), .ZN(n639) );
  NAND2_X1 U628 ( .A1(n622), .A2(n639), .ZN(n540) );
  NOR2_X1 U629 ( .A1(n539), .A2(n538), .ZN(n628) );
  INV_X1 U630 ( .A(n628), .ZN(n640) );
  NAND2_X1 U631 ( .A1(n539), .A2(n538), .ZN(n636) );
  NAND2_X1 U632 ( .A1(n640), .A2(n636), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n540), .A2(n576), .ZN(n543) );
  NOR2_X1 U634 ( .A1(n665), .A2(n541), .ZN(n542) );
  NAND2_X1 U635 ( .A1(n561), .A2(n542), .ZN(n617) );
  NAND2_X1 U636 ( .A1(n650), .A2(n669), .ZN(n547) );
  XNOR2_X1 U637 ( .A(KEYINPUT103), .B(KEYINPUT30), .ZN(n546) );
  XNOR2_X1 U638 ( .A(n547), .B(n546), .ZN(n552) );
  NAND2_X1 U639 ( .A1(G953), .A2(G900), .ZN(n548) );
  NAND2_X1 U640 ( .A1(n549), .A2(n548), .ZN(n558) );
  NOR2_X1 U641 ( .A1(n550), .A2(n558), .ZN(n551) );
  NAND2_X1 U642 ( .A1(n552), .A2(n551), .ZN(n572) );
  INV_X1 U643 ( .A(n553), .ZN(n573) );
  XOR2_X1 U644 ( .A(KEYINPUT38), .B(n573), .Z(n591) );
  NOR2_X1 U645 ( .A1(n572), .A2(n591), .ZN(n556) );
  OR2_X1 U646 ( .A1(n596), .A2(n640), .ZN(n645) );
  NOR2_X1 U647 ( .A1(n666), .A2(n558), .ZN(n559) );
  NAND2_X1 U648 ( .A1(n559), .A2(n665), .ZN(n560) );
  XNOR2_X1 U649 ( .A(KEYINPUT68), .B(n560), .ZN(n565) );
  AND2_X1 U650 ( .A1(n585), .A2(n561), .ZN(n562) );
  NAND2_X1 U651 ( .A1(n562), .A2(n650), .ZN(n563) );
  XNOR2_X1 U652 ( .A(n563), .B(KEYINPUT43), .ZN(n564) );
  NAND2_X1 U653 ( .A1(n564), .A2(n573), .ZN(n646) );
  XNOR2_X1 U654 ( .A(KEYINPUT104), .B(KEYINPUT28), .ZN(n568) );
  NOR2_X1 U655 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U656 ( .A1(KEYINPUT80), .A2(n634), .ZN(n570) );
  NAND2_X1 U657 ( .A1(n570), .A2(n576), .ZN(n571) );
  NAND2_X1 U658 ( .A1(n571), .A2(KEYINPUT47), .ZN(n584) );
  NOR2_X1 U659 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U660 ( .A1(n575), .A2(n574), .ZN(n633) );
  INV_X1 U661 ( .A(n576), .ZN(n655) );
  NOR2_X1 U662 ( .A1(KEYINPUT47), .A2(n655), .ZN(n577) );
  XNOR2_X1 U663 ( .A(KEYINPUT75), .B(n577), .ZN(n578) );
  NAND2_X1 U664 ( .A1(n578), .A2(KEYINPUT80), .ZN(n579) );
  NAND2_X1 U665 ( .A1(n579), .A2(n629), .ZN(n580) );
  NAND2_X1 U666 ( .A1(n633), .A2(n580), .ZN(n582) );
  NOR2_X1 U667 ( .A1(KEYINPUT47), .A2(KEYINPUT80), .ZN(n581) );
  NOR2_X1 U668 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U669 ( .A(n585), .B(KEYINPUT106), .ZN(n587) );
  NAND2_X1 U670 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U671 ( .A(n589), .B(n588), .ZN(n590) );
  INV_X1 U672 ( .A(n591), .ZN(n651) );
  NAND2_X1 U673 ( .A1(n651), .A2(n650), .ZN(n656) );
  NOR2_X1 U674 ( .A1(n656), .A2(n653), .ZN(n593) );
  XOR2_X1 U675 ( .A(KEYINPUT105), .B(KEYINPUT41), .Z(n592) );
  XNOR2_X1 U676 ( .A(n593), .B(n592), .ZN(n676) );
  NOR2_X1 U677 ( .A1(n676), .A2(n594), .ZN(n595) );
  XNOR2_X1 U678 ( .A(KEYINPUT42), .B(n595), .ZN(n736) );
  NOR2_X1 U679 ( .A1(n636), .A2(n596), .ZN(n597) );
  XNOR2_X1 U680 ( .A(n597), .B(KEYINPUT40), .ZN(n737) );
  NOR2_X1 U681 ( .A1(n736), .A2(n737), .ZN(n598) );
  XNOR2_X1 U682 ( .A(n598), .B(KEYINPUT46), .ZN(n599) );
  INV_X1 U683 ( .A(n648), .ZN(n686) );
  INV_X1 U684 ( .A(KEYINPUT2), .ZN(n685) );
  AND2_X1 U685 ( .A1(n685), .A2(n600), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n686), .A2(n601), .ZN(n606) );
  XNOR2_X1 U687 ( .A(n602), .B(KEYINPUT81), .ZN(n603) );
  AND2_X1 U688 ( .A1(KEYINPUT2), .A2(n603), .ZN(n604) );
  NAND2_X1 U689 ( .A1(n648), .A2(n604), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n699), .A2(G472), .ZN(n609) );
  XNOR2_X1 U691 ( .A(n612), .B(n611), .ZN(G57) );
  XNOR2_X1 U692 ( .A(n616), .B(n615), .ZN(G60) );
  XNOR2_X1 U693 ( .A(G101), .B(n617), .ZN(G3) );
  NOR2_X1 U694 ( .A1(n636), .A2(n622), .ZN(n619) );
  XNOR2_X1 U695 ( .A(G104), .B(KEYINPUT109), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n619), .B(n618), .ZN(G6) );
  XOR2_X1 U697 ( .A(KEYINPUT112), .B(KEYINPUT27), .Z(n621) );
  XNOR2_X1 U698 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n621), .B(n620), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n640), .A2(n622), .ZN(n624) );
  XNOR2_X1 U701 ( .A(G107), .B(KEYINPUT26), .ZN(n623) );
  XNOR2_X1 U702 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n626), .B(n625), .ZN(G9) );
  XOR2_X1 U704 ( .A(G110), .B(n627), .Z(G12) );
  XOR2_X1 U705 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n631) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n631), .B(n630), .ZN(n632) );
  XOR2_X1 U708 ( .A(G128), .B(n632), .Z(G30) );
  XNOR2_X1 U709 ( .A(G143), .B(n633), .ZN(G45) );
  OR2_X1 U710 ( .A1(n634), .A2(n636), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(G146), .ZN(G48) );
  NOR2_X1 U712 ( .A1(n636), .A2(n639), .ZN(n637) );
  XOR2_X1 U713 ( .A(KEYINPUT114), .B(n637), .Z(n638) );
  XNOR2_X1 U714 ( .A(G113), .B(n638), .ZN(G15) );
  NOR2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n642) );
  XNOR2_X1 U716 ( .A(G116), .B(KEYINPUT115), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n642), .B(n641), .ZN(G18) );
  XOR2_X1 U718 ( .A(G125), .B(KEYINPUT37), .Z(n643) );
  XNOR2_X1 U719 ( .A(n644), .B(n643), .ZN(G27) );
  XNOR2_X1 U720 ( .A(G134), .B(n645), .ZN(G36) );
  XNOR2_X1 U721 ( .A(G140), .B(n646), .ZN(G42) );
  NOR2_X1 U722 ( .A1(n676), .A2(n661), .ZN(n647) );
  NOR2_X1 U723 ( .A1(G953), .A2(n647), .ZN(n684) );
  AND2_X1 U724 ( .A1(KEYINPUT2), .A2(n648), .ZN(n682) );
  NAND2_X1 U725 ( .A1(G952), .A2(n649), .ZN(n679) );
  NOR2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U728 ( .A(n654), .B(KEYINPUT118), .ZN(n658) );
  NOR2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U731 ( .A(KEYINPUT119), .B(n659), .Z(n660) );
  NOR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U733 ( .A(KEYINPUT50), .B(n664), .Z(n672) );
  NAND2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(KEYINPUT49), .B(n667), .ZN(n668) );
  NOR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U737 ( .A(KEYINPUT116), .B(n670), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U740 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U741 ( .A(KEYINPUT121), .B(n680), .Z(n681) );
  NOR2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n688) );
  AND2_X1 U744 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U745 ( .A(n689), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U746 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n691) );
  XNOR2_X1 U747 ( .A(KEYINPUT87), .B(KEYINPUT55), .ZN(n690) );
  XNOR2_X1 U748 ( .A(n691), .B(n690), .ZN(n692) );
  XOR2_X1 U749 ( .A(n693), .B(n692), .Z(n695) );
  NAND2_X1 U750 ( .A1(n699), .A2(G210), .ZN(n694) );
  XNOR2_X1 U751 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U752 ( .A(n697), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U753 ( .A1(G478), .A2(n699), .ZN(n700) );
  XNOR2_X1 U754 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n706), .A2(n702), .ZN(G63) );
  NAND2_X1 U756 ( .A1(G217), .A2(n699), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U758 ( .A1(n706), .A2(n705), .ZN(G66) );
  NAND2_X1 U759 ( .A1(n716), .A2(n707), .ZN(n711) );
  NAND2_X1 U760 ( .A1(G953), .A2(G224), .ZN(n708) );
  XNOR2_X1 U761 ( .A(KEYINPUT61), .B(n708), .ZN(n709) );
  NAND2_X1 U762 ( .A1(n709), .A2(G898), .ZN(n710) );
  NAND2_X1 U763 ( .A1(n711), .A2(n710), .ZN(n720) );
  XOR2_X1 U764 ( .A(KEYINPUT123), .B(n712), .Z(n715) );
  XNOR2_X1 U765 ( .A(G101), .B(n713), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n715), .B(n714), .ZN(n718) );
  NOR2_X1 U767 ( .A1(G898), .A2(n716), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U769 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U770 ( .A(KEYINPUT124), .B(n721), .ZN(G69) );
  XOR2_X1 U771 ( .A(n723), .B(n722), .Z(n728) );
  XNOR2_X1 U772 ( .A(G227), .B(n728), .ZN(n724) );
  NAND2_X1 U773 ( .A1(n724), .A2(G900), .ZN(n725) );
  NAND2_X1 U774 ( .A1(n725), .A2(G953), .ZN(n726) );
  XOR2_X1 U775 ( .A(KEYINPUT126), .B(n726), .Z(n732) );
  XNOR2_X1 U776 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U777 ( .A1(G953), .A2(n729), .ZN(n730) );
  XOR2_X1 U778 ( .A(KEYINPUT125), .B(n730), .Z(n731) );
  NOR2_X1 U779 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U780 ( .A(KEYINPUT127), .B(n733), .ZN(G72) );
  XOR2_X1 U781 ( .A(n734), .B(G122), .Z(G24) );
  XOR2_X1 U782 ( .A(n735), .B(G119), .Z(G21) );
  XOR2_X1 U783 ( .A(G137), .B(n736), .Z(G39) );
  XOR2_X1 U784 ( .A(G131), .B(n737), .Z(G33) );
endmodule

