//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  NAND2_X1  g0006(.A1(G97), .A2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G116), .ZN(new_n211));
  INV_X1    g0011(.A(G270), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AND2_X1   g0013(.A1(G68), .A2(G238), .ZN(new_n214));
  AND2_X1   g0014(.A1(G107), .A2(G264), .ZN(new_n215));
  NOR4_X1   g0015(.A1(new_n210), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n203), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT64), .Z(new_n231));
  AOI211_X1 g0031(.A(new_n206), .B(new_n226), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n212), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G222), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G223), .A2(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n256), .B(new_n257), .C1(G77), .C2(new_n252), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n259), .B(G274), .C1(G41), .C2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  OAI211_X1 g0061(.A(G1), .B(G13), .C1(new_n249), .C2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G226), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n258), .A2(new_n260), .A3(new_n265), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n266), .A2(G179), .ZN(new_n267));
  INV_X1    g0067(.A(G169), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G50), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n273), .A2(new_n227), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n270), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n259), .A2(G20), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(KEYINPUT66), .A3(G50), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(KEYINPUT66), .B1(new_n276), .B2(G50), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n275), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n273), .A2(new_n227), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G150), .ZN(new_n284));
  NOR3_X1   g0084(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(new_n228), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n228), .A2(G33), .ZN(new_n287));
  AND2_X1   g0087(.A1(KEYINPUT8), .A2(G58), .ZN(new_n288));
  NOR2_X1   g0088(.A1(KEYINPUT8), .A2(G58), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n282), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(KEYINPUT65), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT65), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G58), .A2(G68), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n217), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G20), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n249), .A2(G20), .ZN(new_n297));
  OR2_X1    g0097(.A1(KEYINPUT8), .A2(G58), .ZN(new_n298));
  NAND2_X1  g0098(.A1(KEYINPUT8), .A2(G58), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n296), .A2(new_n300), .A3(new_n284), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n293), .B1(new_n301), .B2(new_n282), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n272), .B(new_n281), .C1(new_n292), .C2(new_n302), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n267), .A2(new_n269), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n266), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n291), .A2(KEYINPUT65), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n293), .A3(new_n282), .ZN(new_n308));
  AOI211_X1 g0108(.A(new_n271), .B(new_n280), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n306), .B1(new_n309), .B2(KEYINPUT9), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n266), .A2(G200), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT69), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT9), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n303), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n312), .B1(new_n303), .B2(new_n313), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n310), .B(new_n311), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT10), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT69), .B1(new_n309), .B2(KEYINPUT9), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n303), .A2(new_n312), .A3(new_n313), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT10), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(new_n311), .A4(new_n310), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n304), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT13), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n223), .A2(G1698), .ZN(new_n325));
  AND2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n325), .B1(G226), .B2(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  AND3_X1   g0128(.A1(KEYINPUT70), .A2(G33), .A3(G97), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT70), .B1(G33), .B2(G97), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n262), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n262), .A2(G238), .A3(new_n263), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n260), .B(KEYINPUT71), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n324), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NOR4_X1   g0137(.A1(new_n332), .A2(new_n335), .A3(new_n333), .A4(KEYINPUT13), .ZN(new_n338));
  OAI21_X1  g0138(.A(G169), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n340));
  INV_X1    g0140(.A(new_n337), .ZN(new_n341));
  INV_X1    g0141(.A(new_n338), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(G179), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(G169), .C1(new_n337), .C2(new_n338), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n340), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n283), .A2(G50), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT72), .ZN(new_n348));
  INV_X1    g0148(.A(G68), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G20), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n297), .A2(G77), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT72), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n283), .A2(new_n352), .A3(G50), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n348), .A2(new_n350), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n282), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT11), .ZN(new_n356));
  INV_X1    g0156(.A(new_n270), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT67), .B1(new_n357), .B2(new_n282), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT67), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n270), .A2(new_n359), .A3(new_n227), .A4(new_n273), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(G68), .A3(new_n276), .ZN(new_n362));
  INV_X1    g0162(.A(G13), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(G1), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n350), .ZN(new_n366));
  XOR2_X1   g0166(.A(new_n366), .B(KEYINPUT12), .Z(new_n367));
  NAND3_X1  g0167(.A1(new_n356), .A2(new_n362), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT73), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n356), .A2(new_n370), .A3(new_n362), .A4(new_n367), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n346), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n298), .A2(new_n299), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(new_n283), .B1(G20), .B2(G77), .ZN(new_n376));
  XOR2_X1   g0176(.A(KEYINPUT15), .B(G87), .Z(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n376), .B1(new_n287), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n282), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n357), .A2(new_n219), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n361), .A2(G77), .A3(new_n276), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G238), .A2(G1698), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n252), .B(new_n384), .C1(new_n223), .C2(G1698), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n385), .B(new_n257), .C1(G107), .C2(new_n252), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n264), .A2(G244), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n260), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n383), .B1(G190), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G200), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n388), .A2(new_n268), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n383), .A2(KEYINPUT68), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT68), .B1(new_n383), .B2(new_n395), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n388), .A2(G179), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n323), .A2(new_n373), .A3(new_n394), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G283), .ZN(new_n403));
  INV_X1    g0203(.A(G97), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n228), .C1(G33), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n211), .A2(G20), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n282), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT20), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n405), .A2(KEYINPUT20), .A3(new_n282), .A4(new_n406), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT80), .B1(new_n270), .B2(G116), .ZN(new_n411));
  OR3_X1    g0211(.A1(new_n270), .A2(KEYINPUT80), .A3(G116), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n409), .A2(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT79), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n259), .A2(G33), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G116), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n414), .B1(new_n361), .B2(new_n417), .ZN(new_n418));
  AOI211_X1 g0218(.A(KEYINPUT79), .B(new_n416), .C1(new_n358), .C2(new_n360), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n413), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n253), .A2(G257), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G264), .A2(G1698), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n421), .B(new_n422), .C1(new_n326), .C2(new_n327), .ZN(new_n423));
  INV_X1    g0223(.A(G303), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n250), .A2(new_n424), .A3(new_n251), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n257), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G45), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(G1), .ZN(new_n428));
  NAND2_X1  g0228(.A1(KEYINPUT5), .A2(G41), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(KEYINPUT5), .A2(G41), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(G270), .A3(new_n262), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n259), .A2(G45), .ZN(new_n434));
  OR2_X1    g0234(.A1(KEYINPUT5), .A2(G41), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(new_n429), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G274), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n426), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n420), .A2(G169), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT21), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AND4_X1   g0241(.A1(G179), .A2(new_n426), .A3(new_n433), .A4(new_n437), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n420), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n420), .A2(KEYINPUT21), .A3(G169), .A4(new_n438), .ZN(new_n444));
  INV_X1    g0244(.A(new_n420), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n438), .A2(new_n305), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(G200), .B2(new_n438), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n441), .A2(new_n443), .A3(new_n444), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n297), .A2(G116), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n228), .A2(G107), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT23), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n208), .A2(KEYINPUT81), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(new_n228), .C1(new_n327), .C2(new_n326), .ZN(new_n454));
  XOR2_X1   g0254(.A(KEYINPUT82), .B(KEYINPUT22), .Z(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n457));
  AOI21_X1  g0257(.A(G20), .B1(new_n250), .B2(new_n251), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n450), .B(new_n452), .C1(new_n456), .C2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT24), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n454), .B(new_n455), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n463), .A2(KEYINPUT24), .A3(new_n450), .A4(new_n452), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n464), .A3(new_n282), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n357), .A2(new_n282), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n415), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G107), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n364), .A2(new_n451), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n470), .B(KEYINPUT25), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n465), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(G257), .A2(G1698), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n326), .B2(new_n327), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT83), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G294), .ZN(new_n477));
  OAI211_X1 g0277(.A(G250), .B(new_n253), .C1(new_n326), .C2(new_n327), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT83), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n479), .B(new_n474), .C1(new_n326), .C2(new_n327), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n476), .A2(new_n477), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n257), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n436), .A2(new_n257), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G264), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n437), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n268), .ZN(new_n486));
  INV_X1    g0286(.A(new_n485), .ZN(new_n487));
  INV_X1    g0287(.A(G179), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n473), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n487), .A2(new_n391), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n485), .A2(new_n305), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n473), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT4), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G1698), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n496), .B(G244), .C1(new_n327), .C2(new_n326), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n220), .B1(new_n250), .B2(new_n251), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n497), .B(new_n403), .C1(new_n498), .C2(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g0299(.A(G250), .B1(new_n326), .B2(new_n327), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n253), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n257), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n432), .A2(G257), .A3(new_n262), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n437), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT77), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT77), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n502), .A2(new_n508), .A3(new_n505), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(G200), .A3(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n467), .A2(new_n404), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n357), .A2(new_n404), .ZN(new_n512));
  XOR2_X1   g0312(.A(new_n512), .B(KEYINPUT76), .Z(new_n513));
  NAND3_X1  g0313(.A1(new_n250), .A2(new_n228), .A3(new_n251), .ZN(new_n514));
  XNOR2_X1  g0314(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n228), .A4(new_n251), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G107), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n283), .A2(G77), .ZN(new_n520));
  INV_X1    g0320(.A(G107), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(KEYINPUT6), .A3(G97), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n404), .A2(new_n521), .ZN(new_n523));
  NOR2_X1   g0323(.A1(G97), .A2(G107), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n522), .B1(new_n525), .B2(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G20), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n519), .A2(new_n520), .A3(new_n527), .ZN(new_n528));
  AOI211_X1 g0328(.A(new_n511), .B(new_n513), .C1(new_n528), .C2(new_n282), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT78), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n506), .B2(new_n305), .ZN(new_n531));
  OAI21_X1  g0331(.A(G244), .B1(new_n326), .B2(new_n327), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(new_n495), .B1(G33), .B2(G283), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n495), .B1(new_n252), .B2(G250), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n497), .C1(new_n253), .C2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n504), .B1(new_n535), .B2(new_n257), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(KEYINPUT78), .A3(G190), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n510), .A2(new_n529), .A3(new_n531), .A4(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n511), .B1(new_n528), .B2(new_n282), .ZN(new_n539));
  INV_X1    g0339(.A(new_n513), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n506), .A2(new_n268), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n488), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n377), .A2(new_n270), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n458), .A2(G68), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n287), .B2(new_n404), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n329), .A2(new_n330), .ZN(new_n549));
  AOI21_X1  g0349(.A(G20), .B1(new_n549), .B2(KEYINPUT19), .ZN(new_n550));
  NOR3_X1   g0350(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n546), .B(new_n548), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n545), .B1(new_n552), .B2(new_n282), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n468), .A2(new_n377), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n434), .A2(new_n209), .ZN(new_n555));
  INV_X1    g0355(.A(G274), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n259), .A2(new_n556), .A3(G45), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n262), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n220), .A2(G1698), .ZN(new_n559));
  OAI221_X1 g0359(.A(new_n559), .B1(G238), .B2(G1698), .C1(new_n326), .C2(new_n327), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G116), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n558), .B1(new_n562), .B2(new_n257), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n553), .A2(new_n554), .B1(new_n268), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n488), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n467), .A2(new_n208), .ZN(new_n567));
  AOI211_X1 g0367(.A(new_n545), .B(new_n567), .C1(new_n552), .C2(new_n282), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(G190), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n262), .B1(new_n560), .B2(new_n561), .ZN(new_n570));
  OAI21_X1  g0370(.A(G200), .B1(new_n570), .B2(new_n558), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n565), .A2(new_n566), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n538), .A2(new_n544), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n494), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n262), .A2(G232), .A3(new_n263), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n250), .A2(new_n251), .B1(new_n218), .B2(G1698), .ZN(new_n577));
  OR2_X1    g0377(.A1(G223), .A2(G1698), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n577), .A2(new_n578), .B1(G33), .B2(G87), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n576), .B(new_n260), .C1(new_n579), .C2(new_n262), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n391), .ZN(new_n581));
  OAI221_X1 g0381(.A(new_n578), .B1(G226), .B2(new_n253), .C1(new_n326), .C2(new_n327), .ZN(new_n582));
  NAND2_X1  g0382(.A1(G33), .A2(G87), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n257), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n585), .A2(new_n305), .A3(new_n576), .A4(new_n260), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(G58), .A2(G68), .ZN(new_n588));
  OAI21_X1  g0388(.A(G20), .B1(new_n588), .B2(new_n294), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT75), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(KEYINPUT75), .B(G20), .C1(new_n588), .C2(new_n294), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n326), .A2(new_n327), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n515), .A3(new_n228), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n514), .A2(KEYINPUT7), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(G68), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n283), .A2(G159), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n593), .A2(new_n597), .A3(KEYINPUT16), .A4(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT16), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n349), .B1(new_n516), .B2(new_n517), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n591), .A2(new_n598), .A3(new_n592), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(new_n603), .A3(new_n282), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n375), .A2(new_n274), .A3(new_n276), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n357), .B2(new_n374), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n587), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT17), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n587), .A2(KEYINPUT17), .A3(new_n604), .A4(new_n606), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT18), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n580), .A2(G169), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n585), .A2(G179), .A3(new_n576), .A4(new_n260), .ZN(new_n613));
  AOI221_X4 g0413(.A(new_n611), .B1(new_n612), .B2(new_n613), .C1(new_n604), .C2(new_n606), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n604), .A2(new_n606), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n613), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT18), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n609), .B(new_n610), .C1(new_n614), .C2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n368), .ZN(new_n620));
  OAI21_X1  g0420(.A(G200), .B1(new_n337), .B2(new_n338), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n341), .A2(G190), .A3(new_n342), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NOR4_X1   g0424(.A1(new_n402), .A2(new_n449), .A3(new_n575), .A4(new_n624), .ZN(G372));
  INV_X1    g0425(.A(new_n623), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n401), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n372), .B2(new_n346), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n609), .A2(new_n610), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n628), .A2(new_n629), .B1(new_n617), .B2(new_n614), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n317), .A2(new_n322), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n304), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n402), .A2(new_n624), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n538), .A2(new_n544), .A3(new_n573), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(new_n493), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT84), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n473), .A2(new_n486), .A3(new_n489), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT84), .B1(new_n490), .B2(new_n636), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n635), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  INV_X1    g0443(.A(new_n573), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n643), .B1(new_n644), .B2(new_n544), .ZN(new_n645));
  INV_X1    g0445(.A(new_n544), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(KEYINPUT26), .A3(new_n573), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n645), .A2(new_n647), .B1(new_n566), .B2(new_n565), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n633), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n632), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g0451(.A(new_n651), .B(KEYINPUT85), .Z(G369));
  XOR2_X1   g0452(.A(new_n449), .B(KEYINPUT86), .Z(new_n653));
  OR3_X1    g0453(.A1(new_n365), .A2(KEYINPUT27), .A3(G20), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT27), .B1(new_n365), .B2(G20), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n445), .A2(new_n659), .ZN(new_n660));
  MUX2_X1   g0460(.A(new_n653), .B(new_n636), .S(new_n660), .Z(new_n661));
  AND2_X1   g0461(.A1(new_n473), .A2(new_n658), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n639), .B1(new_n662), .B2(new_n493), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n490), .A2(new_n659), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n661), .A2(G330), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT87), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n666), .B(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n636), .A2(new_n659), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n494), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n664), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT88), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n668), .A2(new_n673), .ZN(G399));
  NAND2_X1  g0474(.A1(new_n551), .A2(new_n211), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n204), .A2(new_n261), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G1), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n230), .B2(new_n677), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n637), .A2(KEYINPUT90), .A3(new_n639), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT90), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n490), .B2(new_n636), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n635), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n658), .B1(new_n684), .B2(new_n648), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT29), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI211_X1 g0487(.A(KEYINPUT29), .B(new_n658), .C1(new_n642), .C2(new_n648), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT31), .ZN(new_n690));
  AND4_X1   g0490(.A1(new_n488), .A2(new_n485), .A3(new_n438), .A4(new_n564), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n482), .A2(new_n563), .A3(new_n484), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(new_n442), .A4(new_n536), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n442), .A2(new_n502), .A3(new_n505), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n482), .A2(new_n563), .A3(new_n484), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT30), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n506), .A2(new_n691), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n658), .B1(new_n698), .B2(KEYINPUT89), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n481), .A2(new_n257), .B1(G264), .B2(new_n483), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n563), .B1(new_n700), .B2(new_n437), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(new_n488), .A3(new_n438), .A4(new_n506), .ZN(new_n702));
  INV_X1    g0502(.A(new_n697), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n695), .A2(new_n696), .A3(KEYINPUT30), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT89), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n690), .B1(new_n699), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n449), .A2(new_n658), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n494), .A2(new_n574), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n689), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n680), .B1(new_n715), .B2(G1), .ZN(G364));
  NAND2_X1  g0516(.A1(new_n661), .A2(G330), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n363), .A2(G20), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G45), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n677), .A2(G1), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(G330), .B2(new_n661), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n722), .B1(new_n661), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n227), .B1(G20), .B2(new_n268), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n231), .A2(new_n427), .ZN(new_n732));
  INV_X1    g0532(.A(new_n204), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n252), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n732), .B(new_n734), .C1(new_n243), .C2(new_n427), .ZN(new_n735));
  INV_X1    g0535(.A(G355), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n252), .A2(new_n204), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n735), .B1(G116), .B2(new_n204), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n729), .B1(new_n731), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n228), .A2(G179), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G190), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT92), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G329), .ZN(new_n744));
  INV_X1    g0544(.A(G294), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n305), .A2(G179), .A3(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n228), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n744), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n228), .A2(new_n488), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n750), .A2(new_n305), .A3(G200), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n252), .B(new_n748), .C1(G322), .C2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n305), .A2(new_n391), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n740), .ZN(new_n754));
  INV_X1    g0554(.A(G326), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n749), .A2(new_n753), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n752), .B1(new_n424), .B2(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n749), .A2(new_n741), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n391), .A2(G190), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n740), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT33), .B(G317), .Z(new_n765));
  NAND2_X1  g0565(.A1(new_n749), .A2(new_n761), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n757), .A2(new_n760), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n758), .ZN(new_n769));
  INV_X1    g0569(.A(new_n762), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G77), .A2(new_n769), .B1(new_n770), .B2(G107), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n771), .B(new_n252), .C1(new_n349), .C2(new_n766), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n747), .B(KEYINPUT91), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G97), .ZN(new_n775));
  INV_X1    g0575(.A(G159), .ZN(new_n776));
  OR3_X1    g0576(.A1(new_n742), .A2(KEYINPUT32), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(KEYINPUT32), .B1(new_n742), .B2(new_n776), .ZN(new_n778));
  INV_X1    g0578(.A(new_n756), .ZN(new_n779));
  INV_X1    g0579(.A(new_n754), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G50), .A2(new_n779), .B1(new_n780), .B2(G87), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n775), .A2(new_n777), .A3(new_n778), .A4(new_n781), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n772), .B(new_n782), .C1(G58), .C2(new_n751), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n730), .B1(new_n768), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n739), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n724), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(G396));
  NAND2_X1  g0587(.A1(new_n743), .A2(G311), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n770), .A2(G87), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n252), .B1(new_n780), .B2(G107), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n775), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n758), .A2(new_n211), .ZN(new_n792));
  INV_X1    g0592(.A(new_n751), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n745), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n756), .A2(new_n424), .B1(new_n766), .B2(new_n763), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n791), .A2(new_n792), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n766), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G137), .A2(new_n779), .B1(new_n797), .B2(G150), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT93), .Z(new_n799));
  INV_X1    g0599(.A(G143), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n799), .B1(new_n800), .B2(new_n793), .C1(new_n776), .C2(new_n758), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT34), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n802), .B1(new_n217), .B2(new_n754), .C1(new_n349), .C2(new_n762), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G132), .B2(new_n743), .ZN(new_n804));
  INV_X1    g0604(.A(new_n747), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n594), .B1(new_n805), .B2(G58), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n796), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT94), .Z(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n730), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n730), .A2(new_n725), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n219), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n383), .A2(new_n658), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n398), .B2(new_n400), .ZN(new_n814));
  NOR4_X1   g0614(.A1(new_n396), .A2(new_n397), .A3(new_n399), .A4(new_n812), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n394), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n725), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n809), .A2(new_n722), .A3(new_n811), .A4(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n658), .B1(new_n642), .B2(new_n648), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(new_n816), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(new_n713), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n721), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n818), .A2(new_n822), .ZN(G384));
  INV_X1    g0623(.A(new_n656), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n615), .B1(new_n616), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n825), .A2(new_n607), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n599), .A2(new_n282), .ZN(new_n827));
  INV_X1    g0627(.A(new_n602), .ZN(new_n828));
  AOI21_X1  g0628(.A(KEYINPUT16), .B1(new_n828), .B2(new_n597), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n606), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n616), .B2(new_n824), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n607), .ZN(new_n832));
  MUX2_X1   g0632(.A(new_n826), .B(new_n832), .S(KEYINPUT37), .Z(new_n833));
  AND2_X1   g0633(.A1(new_n830), .A2(new_n824), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n618), .A2(KEYINPUT97), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT97), .B1(new_n618), .B2(new_n834), .ZN(new_n836));
  OAI211_X1 g0636(.A(KEYINPUT38), .B(new_n833), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT99), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n614), .A2(new_n617), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n834), .B1(new_n840), .B2(new_n629), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT97), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n618), .A2(KEYINPUT97), .A3(new_n834), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n845), .A2(KEYINPUT99), .A3(KEYINPUT38), .A4(new_n833), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n615), .A2(new_n824), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT37), .B1(new_n849), .B2(KEYINPUT98), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(new_n826), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n619), .B2(new_n848), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n839), .A2(new_n846), .B1(new_n847), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT101), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n372), .A2(new_n658), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT95), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n346), .A2(new_n372), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n346), .B2(new_n372), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n623), .B(new_n855), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n372), .B(new_n658), .C1(new_n626), .C2(new_n346), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n816), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT89), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n659), .B1(new_n710), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n707), .A2(new_n709), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n854), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT40), .B1(new_n853), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n816), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n859), .A2(new_n860), .ZN(new_n869));
  NAND2_X1  g0669(.A1(KEYINPUT101), .A2(KEYINPUT40), .ZN(new_n870));
  AND4_X1   g0670(.A1(new_n868), .A2(new_n869), .A3(new_n865), .A4(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n847), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT40), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n874), .A3(new_n837), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n867), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n633), .A2(new_n865), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(G330), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT100), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n633), .B1(new_n687), .B2(new_n688), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n632), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n881), .B(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n401), .A2(new_n658), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n885), .B1(new_n819), .B2(new_n868), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT96), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(new_n869), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n873), .A2(new_n837), .ZN(new_n890));
  INV_X1    g0690(.A(new_n869), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT96), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n840), .A2(new_n656), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n857), .A2(new_n858), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n658), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n873), .A2(KEYINPUT39), .A3(new_n837), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n896), .B(new_n897), .C1(new_n853), .C2(KEYINPUT39), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n893), .A2(new_n894), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n884), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n259), .B2(new_n719), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n211), .B1(new_n526), .B2(KEYINPUT35), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n902), .B(new_n229), .C1(KEYINPUT35), .C2(new_n526), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT36), .ZN(new_n904));
  OAI21_X1  g0704(.A(G77), .B1(new_n222), .B2(new_n349), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n905), .A2(new_n230), .B1(G50), .B2(new_n349), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(G1), .A3(new_n363), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n901), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT102), .Z(G367));
  OAI22_X1  g0709(.A1(new_n793), .A2(new_n424), .B1(new_n404), .B2(new_n762), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n252), .B(new_n910), .C1(G283), .C2(new_n769), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n805), .A2(G107), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n780), .A2(G116), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT46), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n756), .A2(new_n759), .B1(new_n766), .B2(new_n745), .ZN(new_n915));
  INV_X1    g0715(.A(new_n742), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(G317), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n911), .A2(new_n912), .A3(new_n914), .A4(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n774), .A2(G68), .B1(G50), .B2(new_n769), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n222), .B2(new_n754), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n756), .A2(new_n800), .B1(new_n762), .B2(new_n219), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n920), .A2(new_n594), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n916), .A2(G137), .ZN(new_n923));
  INV_X1    g0723(.A(G150), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n922), .B(new_n923), .C1(new_n924), .C2(new_n793), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n766), .A2(new_n776), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n918), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT47), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n730), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n573), .B1(new_n568), .B2(new_n659), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n568), .A2(new_n659), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n566), .A3(new_n565), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n727), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n734), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n731), .B1(new_n204), .B2(new_n378), .C1(new_n239), .C2(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n929), .A2(new_n722), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n720), .A2(G1), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n670), .B1(new_n665), .B2(new_n669), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n717), .B(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT106), .B1(new_n939), .B2(new_n714), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n718), .A2(new_n938), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n717), .B(new_n670), .C1(new_n665), .C2(new_n669), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT106), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(new_n944), .A3(new_n715), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n538), .B(new_n544), .C1(new_n529), .C2(new_n659), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT103), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n646), .A2(new_n658), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n948), .B1(new_n947), .B2(new_n949), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n673), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT45), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT44), .B1(new_n673), .B2(new_n953), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n671), .B(KEYINPUT88), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT44), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n958), .A2(new_n959), .A3(new_n952), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n956), .A2(new_n668), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n666), .B(KEYINPUT87), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n954), .B(KEYINPUT45), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n964), .B1(new_n965), .B2(new_n961), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n946), .A2(new_n963), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n715), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n677), .B(KEYINPUT41), .Z(new_n969));
  AOI21_X1  g0769(.A(new_n937), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n930), .A2(new_n932), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  XOR2_X1   g0772(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n952), .A2(new_n670), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n952), .B2(new_n670), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n646), .B1(new_n953), .B2(new_n490), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n975), .B(new_n976), .C1(new_n977), .C2(new_n658), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT105), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n979), .B1(new_n978), .B2(new_n980), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n972), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n983), .ZN(new_n985));
  INV_X1    g0785(.A(new_n972), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n985), .A2(new_n986), .A3(new_n981), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n668), .A2(new_n952), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n988), .B(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n936), .B1(new_n970), .B2(new_n991), .ZN(G387));
  NAND2_X1  g0792(.A1(new_n943), .A2(new_n715), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n939), .A2(new_n714), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n677), .B(KEYINPUT111), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n734), .B1(new_n236), .B2(new_n427), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n676), .B2(new_n737), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n375), .A2(new_n217), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT108), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n676), .B(new_n427), .C1(new_n349), .C2(new_n219), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n999), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n733), .A2(new_n521), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n730), .B(new_n727), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n722), .B1(new_n665), .B2(new_n728), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n774), .A2(new_n377), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n762), .A2(new_n404), .B1(new_n742), .B2(new_n924), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n594), .B(new_n1010), .C1(G68), .C2(new_n769), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n751), .A2(G50), .B1(new_n375), .B2(new_n797), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G159), .A2(new_n779), .B1(new_n780), .B2(G77), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G322), .A2(new_n779), .B1(new_n797), .B2(G311), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n424), .B2(new_n758), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G317), .B2(new_n751), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT48), .Z(new_n1018));
  AOI22_X1  g0818(.A1(new_n805), .A2(G283), .B1(new_n780), .B2(G294), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT109), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT49), .Z(new_n1024));
  OAI221_X1 g0824(.A(new_n594), .B1(new_n742), .B2(new_n755), .C1(new_n211), .C2(new_n762), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT110), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1014), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1007), .B(new_n1008), .C1(new_n1027), .C2(new_n730), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n943), .B2(new_n937), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n997), .A2(new_n1029), .ZN(G393));
  NOR3_X1   g0830(.A1(new_n965), .A2(new_n964), .A3(new_n961), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n668), .B1(new_n956), .B2(new_n962), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n937), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n773), .A2(new_n219), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n789), .A2(new_n252), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n754), .A2(new_n349), .B1(new_n742), .B2(new_n800), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n374), .B2(new_n758), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT51), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n793), .A2(new_n776), .B1(new_n756), .B2(new_n924), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1035), .B(new_n1039), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n1040), .B2(new_n1041), .C1(new_n217), .C2(new_n766), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n751), .A2(G311), .B1(new_n779), .B2(G317), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT52), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n252), .B1(new_n916), .B2(G322), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n521), .B2(new_n762), .C1(new_n763), .C2(new_n754), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT112), .Z(new_n1048));
  AOI211_X1 g0848(.A(new_n1045), .B(new_n1048), .C1(G116), .C2(new_n805), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n745), .B2(new_n758), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n766), .A2(new_n424), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1043), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n730), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n952), .A2(new_n727), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n731), .B1(new_n404), .B2(new_n204), .C1(new_n246), .C2(new_n934), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n722), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT113), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n995), .B1(new_n1033), .B2(new_n946), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n993), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AND4_X1   g0860(.A1(new_n1057), .A2(new_n967), .A3(new_n1059), .A4(new_n996), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1034), .B(new_n1056), .C1(new_n1060), .C2(new_n1061), .ZN(G390));
  INV_X1    g0862(.A(KEYINPUT53), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n780), .B2(G150), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n751), .A2(G132), .B1(G137), .B2(new_n797), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT54), .B(G143), .Z(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1065), .B(new_n252), .C1(new_n758), .C2(new_n1067), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1064), .B(new_n1068), .C1(G125), .C2(new_n743), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n754), .A2(KEYINPUT53), .A3(new_n924), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n774), .B2(G159), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(new_n217), .C2(new_n762), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G128), .B2(new_n779), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n594), .B1(new_n208), .B2(new_n754), .C1(new_n793), .C2(new_n211), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1035), .B(new_n1074), .C1(G294), .C2(new_n743), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G97), .A2(new_n769), .B1(new_n770), .B2(G68), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n763), .C2(new_n756), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G107), .B2(new_n797), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n730), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n873), .A2(KEYINPUT39), .A3(new_n837), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n839), .A2(new_n846), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n852), .A2(new_n847), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT39), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1080), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n722), .B(new_n1079), .C1(new_n1085), .C2(new_n726), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n374), .B2(new_n810), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n885), .B1(new_n685), .B2(new_n868), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(new_n891), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n896), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n1090), .A3(new_n1083), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n869), .A2(new_n712), .A3(G330), .A4(new_n868), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1090), .B1(new_n886), .B2(new_n891), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1091), .B(new_n1093), .C1(new_n1085), .C2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n861), .A2(G330), .A3(new_n865), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n897), .B1(new_n853), .B2(KEYINPUT39), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n853), .A2(new_n896), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1099), .A2(new_n1094), .B1(new_n1100), .B2(new_n1089), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1096), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1087), .B1(new_n937), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT114), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n865), .A2(G330), .A3(new_n868), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n891), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1106), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n712), .A2(G330), .A3(new_n868), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n891), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n886), .B1(new_n1109), .B2(new_n1097), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n633), .A2(G330), .A3(new_n865), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n882), .A2(new_n632), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1104), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n882), .A2(new_n1112), .A3(new_n632), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1106), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n865), .A2(G330), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1117), .A2(new_n861), .B1(new_n1108), .B2(new_n891), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1118), .B2(new_n886), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(KEYINPUT114), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1102), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1091), .B1(new_n1085), .B2(new_n1095), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1097), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1124), .A2(new_n1114), .A3(new_n1120), .A4(new_n1096), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1122), .B(new_n996), .C1(new_n1125), .C2(KEYINPUT115), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1125), .A2(KEYINPUT115), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1103), .B1(new_n1126), .B2(new_n1127), .ZN(G378));
  XNOR2_X1  g0928(.A(new_n1115), .B(KEYINPUT120), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1122), .A2(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n317), .A2(new_n322), .ZN(new_n1132));
  OAI21_X1  g0932(.A(KEYINPUT119), .B1(new_n1132), .B2(new_n304), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT119), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n323), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n309), .A2(new_n656), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n323), .A2(new_n1134), .ZN(new_n1139));
  AOI211_X1 g0939(.A(KEYINPUT119), .B(new_n304), .C1(new_n317), .C2(new_n322), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1138), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n871), .A2(new_n875), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n866), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1083), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1146), .B1(new_n1148), .B2(KEYINPUT40), .ZN(new_n1149));
  INV_X1    g0949(.A(G330), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1145), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n893), .A2(new_n894), .A3(new_n898), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1145), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n877), .A2(G330), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n877), .B2(G330), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1150), .B(new_n1145), .C1(new_n867), .C2(new_n876), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n899), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1131), .A2(KEYINPUT57), .A3(new_n1155), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1155), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1129), .B1(new_n1102), .B2(new_n1121), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1159), .A2(new_n996), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1158), .A2(new_n1155), .A3(new_n937), .ZN(new_n1165));
  INV_X1    g0965(.A(G124), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n249), .B1(new_n742), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n773), .A2(new_n924), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1067), .A2(new_n754), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT116), .ZN(new_n1170));
  INV_X1    g0970(.A(G125), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(new_n756), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1168), .B(new_n1172), .C1(G137), .C2(new_n769), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n797), .A2(G132), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n751), .A2(G128), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G41), .B(new_n1167), .C1(new_n1176), .C2(KEYINPUT59), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(KEYINPUT59), .B2(new_n1176), .C1(new_n776), .C2(new_n762), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n774), .A2(G68), .B1(G283), .B2(new_n743), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n219), .B2(new_n754), .C1(new_n404), .C2(new_n766), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G41), .B(new_n1180), .C1(G107), .C2(new_n751), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n252), .B1(new_n770), .B2(G58), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n769), .A2(new_n377), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n779), .A2(G116), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT58), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n217), .B1(new_n326), .B2(G41), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1178), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n730), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT117), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1153), .A2(new_n725), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n721), .B1(new_n217), .B2(new_n810), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(KEYINPUT118), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1192), .A2(KEYINPUT118), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1165), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1164), .A2(new_n1197), .ZN(G375));
  NOR2_X1   g0998(.A1(new_n869), .A2(new_n726), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT121), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n810), .A2(new_n349), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1009), .B1(new_n219), .B2(new_n762), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n252), .B1(new_n743), .B2(G303), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n521), .B2(new_n758), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n793), .A2(new_n763), .B1(new_n404), .B2(new_n754), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n211), .B2(new_n766), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n756), .A2(new_n745), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n773), .A2(new_n217), .B1(new_n924), .B2(new_n758), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n594), .B(new_n1209), .C1(G58), .C2(new_n770), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n797), .A2(new_n1066), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n743), .A2(G128), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n751), .A2(G137), .B1(new_n779), .B2(G132), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n754), .A2(new_n776), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n1207), .A2(new_n1208), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n721), .B1(new_n1216), .B2(new_n730), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1200), .A2(new_n1201), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n937), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1218), .B1(new_n1111), .B2(new_n1219), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT122), .Z(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n969), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1222), .B1(new_n1121), .B2(new_n1225), .ZN(G381));
  NOR2_X1   g1026(.A1(G375), .A2(G378), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(G387), .A2(G384), .A3(G381), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(G407));
  INV_X1    g1030(.A(G213), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1227), .B2(new_n657), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(G407), .ZN(G409));
  OR2_X1    g1033(.A1(new_n1125), .A2(KEYINPUT115), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1125), .A2(KEYINPUT115), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1234), .A2(new_n996), .A3(new_n1235), .A4(new_n1122), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1164), .A2(new_n1197), .B1(new_n1236), .B2(new_n1103), .ZN(new_n1237));
  INV_X1    g1037(.A(G384), .ZN(new_n1238));
  XOR2_X1   g1038(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n1239));
  NAND3_X1  g1039(.A1(new_n1114), .A2(new_n1120), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT124), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1240), .A2(new_n1241), .A3(new_n1224), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(new_n1240), .B2(new_n1224), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n995), .B1(new_n1223), .B2(KEYINPUT60), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1238), .B1(new_n1246), .B2(new_n1221), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1240), .A2(new_n1224), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT124), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1240), .A2(new_n1241), .A3(new_n1224), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(new_n1244), .A3(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(G384), .A3(new_n1222), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1247), .A2(new_n1252), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1124), .A2(new_n1096), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1155), .B(new_n1158), .C1(new_n1254), .C2(new_n1129), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n969), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1165), .B(new_n1195), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(G378), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1231), .A2(G343), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(new_n1237), .A2(new_n1253), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1259), .ZN(new_n1261));
  INV_X1    g1061(.A(G378), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1196), .B1(new_n969), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n995), .B1(new_n1263), .B2(KEYINPUT57), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1196), .B1(new_n1266), .B2(new_n1163), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1261), .B(new_n1265), .C1(new_n1267), .C2(new_n1262), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1252), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G384), .B1(new_n1251), .B2(new_n1222), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1259), .A2(G2897), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1272), .B1(new_n1247), .B2(new_n1252), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1268), .A2(new_n1273), .A3(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1260), .B1(new_n1276), .B2(KEYINPUT63), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n936), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n714), .B1(new_n1033), .B2(new_n946), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1219), .B1(new_n1279), .B2(new_n1256), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n988), .B(new_n989), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1278), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT126), .B1(G390), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G390), .A2(new_n1282), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(G393), .B(new_n786), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(G390), .A2(new_n1282), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1286), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1286), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT125), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1290), .B1(new_n1287), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1058), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n967), .A2(new_n1059), .A3(new_n996), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT113), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(G387), .A2(new_n1034), .A3(new_n1296), .A4(new_n1056), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(new_n1284), .A3(KEYINPUT125), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1285), .A2(new_n1289), .B1(new_n1292), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G375), .A2(G378), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1301), .A2(new_n1271), .A3(new_n1261), .A4(new_n1265), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1300), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(new_n1277), .A2(new_n1299), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1298), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1286), .B1(new_n1297), .B2(KEYINPUT125), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1290), .B1(new_n1297), .B2(KEYINPUT126), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1309));
  OAI22_X1  g1109(.A1(new_n1306), .A2(new_n1307), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1272), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1269), .A2(new_n1270), .A3(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1312), .A2(new_n1274), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(KEYINPUT62), .A2(new_n1302), .B1(new_n1313), .B2(new_n1268), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT62), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT61), .B1(new_n1260), .B2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1310), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(KEYINPUT127), .B1(new_n1305), .B2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1276), .B1(new_n1260), .B2(new_n1315), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1300), .B1(new_n1302), .B2(KEYINPUT62), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1299), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT127), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1303), .B1(new_n1313), .B2(new_n1268), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1310), .B1(new_n1323), .B2(new_n1260), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1321), .B(new_n1322), .C1(new_n1304), .C2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1318), .A2(new_n1325), .ZN(G405));
  OAI21_X1  g1126(.A(new_n1299), .B1(new_n1227), .B2(new_n1237), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1227), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1310), .A2(new_n1328), .A3(new_n1301), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1327), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1253), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1327), .A2(new_n1329), .A3(new_n1271), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(G402));
endmodule


