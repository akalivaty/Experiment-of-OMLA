//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1227, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n211), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  INV_X1    g0021(.A(new_n206), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n223), .A2(G50), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT65), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n231), .B1(new_n211), .B2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(G13), .ZN(new_n233));
  NAND4_X1  g0033(.A1(new_n233), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n235), .B(G250), .C1(G257), .C2(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT0), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n221), .A2(new_n230), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n238), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n252), .B(new_n253), .Z(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G222), .A3(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G77), .ZN(new_n262));
  OAI211_X1 g0062(.A(G223), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n258), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  OAI211_X1 g0068(.A(G1), .B(G13), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G1), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT69), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G45), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n278), .A3(new_n268), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n272), .A2(G226), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n266), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT70), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n266), .A2(KEYINPUT70), .A3(new_n280), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G200), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT75), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT10), .ZN(new_n288));
  INV_X1    g0088(.A(new_n284), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT70), .B1(new_n266), .B2(new_n280), .ZN(new_n290));
  OAI21_X1  g0090(.A(G190), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n283), .A2(KEYINPUT75), .A3(G200), .A4(new_n284), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n287), .A2(new_n288), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT71), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(new_n211), .B2(new_n267), .ZN(new_n296));
  NAND4_X1  g0096(.A1(KEYINPUT71), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n227), .A3(new_n297), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n233), .A2(new_n228), .A3(G1), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n270), .A2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G50), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n300), .A2(new_n303), .B1(new_n207), .B2(new_n299), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT8), .B(G58), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT72), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n228), .A2(G33), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT8), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n309), .A2(KEYINPUT72), .A3(G58), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n306), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G20), .A2(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G150), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT73), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n208), .A2(new_n316), .A3(G20), .ZN(new_n317));
  AOI21_X1  g0117(.A(G50), .B1(new_n204), .B2(new_n205), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT73), .B1(new_n318), .B2(new_n228), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n315), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n296), .A2(new_n227), .A3(new_n297), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n294), .B(new_n304), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n317), .A2(new_n319), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n310), .B1(new_n305), .B2(KEYINPUT72), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n308), .B1(G150), .B2(new_n313), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n321), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n304), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT9), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT74), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n322), .A2(new_n328), .A3(KEYINPUT74), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n293), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT76), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n322), .A2(new_n328), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n291), .A2(new_n285), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n332), .B(KEYINPUT10), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT10), .B1(new_n333), .B2(new_n334), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT76), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n331), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G97), .ZN(new_n340));
  OAI211_X1 g0140(.A(G226), .B(new_n257), .C1(new_n259), .C2(new_n260), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n265), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT13), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n272), .A2(G238), .B1(new_n274), .B2(new_n279), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g0148(.A(G200), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G77), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n307), .A2(new_n350), .B1(new_n228), .B2(G68), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT77), .ZN(new_n352));
  INV_X1    g0152(.A(new_n313), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n207), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n313), .A2(KEYINPUT77), .A3(G50), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT11), .ZN(new_n357));
  OR3_X1    g0157(.A1(new_n356), .A2(new_n357), .A3(new_n321), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n299), .A2(new_n203), .ZN(new_n359));
  NOR2_X1   g0159(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n360), .B2(new_n359), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n357), .B1(new_n356), .B2(new_n321), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n300), .A2(G68), .A3(new_n301), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n358), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n343), .A2(new_n345), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT13), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(G190), .A3(new_n346), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n349), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(G169), .B1(new_n347), .B2(new_n348), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT79), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT14), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  OAI221_X1 g0177(.A(G169), .B1(new_n374), .B2(new_n375), .C1(new_n347), .C2(new_n348), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n369), .A2(G179), .A3(new_n346), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n372), .B1(new_n380), .B2(new_n366), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  OR2_X1    g0182(.A1(KEYINPUT3), .A2(G33), .ZN(new_n383));
  NAND2_X1  g0183(.A1(KEYINPUT3), .A2(G33), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n228), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n383), .A2(KEYINPUT7), .A3(new_n228), .A4(new_n384), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n203), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G58), .A2(G68), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n204), .A2(new_n205), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G20), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n313), .A2(G159), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n382), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n261), .B2(new_n228), .ZN(new_n396));
  INV_X1    g0196(.A(new_n388), .ZN(new_n397));
  OAI21_X1  g0197(.A(G68), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n391), .A2(G20), .B1(G159), .B2(new_n313), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(KEYINPUT16), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n395), .A2(new_n400), .A3(new_n298), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n306), .A2(KEYINPUT80), .A3(new_n311), .A4(new_n301), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n402), .A2(new_n300), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT80), .B1(new_n324), .B2(new_n301), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n324), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n403), .A2(new_n405), .B1(new_n299), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G87), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n267), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(G223), .A2(G1698), .ZN(new_n411));
  INV_X1    g0211(.A(G226), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(G1698), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n410), .B1(new_n413), .B2(new_n256), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT81), .B1(new_n414), .B2(new_n269), .ZN(new_n415));
  OR2_X1    g0215(.A1(G223), .A2(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(G1698), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(new_n259), .C2(new_n260), .ZN(new_n418));
  INV_X1    g0218(.A(new_n410), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n269), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT81), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n279), .A2(new_n274), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n269), .A2(G232), .A3(new_n271), .ZN(new_n424));
  INV_X1    g0224(.A(G179), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n415), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G169), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n423), .A2(new_n424), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(new_n420), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT82), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n427), .A2(KEYINPUT82), .A3(new_n430), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n408), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT18), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n408), .A2(new_n433), .A3(new_n437), .A4(new_n434), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G190), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n423), .A2(new_n424), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n415), .A2(new_n422), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G200), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n429), .B2(new_n420), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n401), .A2(new_n445), .A3(new_n407), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT17), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n401), .A2(new_n445), .A3(new_n407), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n256), .A2(G232), .A3(new_n257), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n256), .A2(G238), .A3(G1698), .ZN(new_n453));
  INV_X1    g0253(.A(G107), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(new_n256), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n265), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n272), .A2(G244), .B1(new_n274), .B2(new_n279), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n425), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n300), .A2(G77), .A3(new_n301), .ZN(new_n461));
  INV_X1    g0261(.A(new_n299), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n305), .A2(new_n353), .B1(new_n228), .B2(new_n350), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT15), .B(G87), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n463), .B1(new_n308), .B2(new_n465), .ZN(new_n466));
  OAI221_X1 g0266(.A(new_n461), .B1(G77), .B2(new_n462), .C1(new_n466), .C2(new_n321), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n458), .A2(new_n428), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n460), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n458), .A2(G200), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n467), .B1(new_n459), .B2(G190), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n381), .A2(new_n439), .A3(new_n451), .A4(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n425), .B1(new_n289), .B2(new_n290), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n304), .B1(new_n320), .B2(new_n321), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n283), .A2(new_n428), .A3(new_n284), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n338), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n228), .C1(G33), .C2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT86), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G20), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n298), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n483), .B1(new_n298), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n482), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(KEYINPUT20), .B(new_n482), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n270), .A2(G33), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n300), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G116), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n462), .A2(new_n484), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n256), .A2(G264), .A3(G1698), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n256), .A2(G257), .A3(new_n257), .ZN(new_n500));
  INV_X1    g0300(.A(G303), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n499), .B(new_n500), .C1(new_n501), .C2(new_n256), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n265), .ZN(new_n503));
  AND2_X1   g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  NOR2_X1   g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n270), .B(G45), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(G270), .A3(new_n269), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT5), .B(G41), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n508), .A2(new_n270), .A3(G45), .A4(G274), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n507), .A2(KEYINPUT85), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT85), .B1(new_n507), .B2(new_n509), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n503), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G169), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n498), .A2(KEYINPUT21), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT21), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n490), .A2(new_n491), .B1(new_n495), .B2(new_n496), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n517), .B2(new_n513), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n503), .B(G179), .C1(new_n510), .C2(new_n511), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n498), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n515), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  OR2_X1    g0323(.A1(new_n512), .A2(new_n440), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n512), .A2(G200), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n517), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n524), .A2(new_n517), .A3(KEYINPUT87), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(G244), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n531));
  OAI211_X1 g0331(.A(G238), .B(new_n257), .C1(new_n259), .C2(new_n260), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(new_n532), .C1(new_n267), .C2(new_n484), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n265), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n274), .A2(G45), .ZN(new_n535));
  OAI21_X1  g0335(.A(G250), .B1(new_n275), .B2(G1), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(new_n265), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n534), .A2(new_n425), .A3(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n321), .A2(new_n462), .A3(new_n493), .A4(new_n465), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT19), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n228), .B1(new_n340), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n409), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n228), .B(G68), .C1(new_n259), .C2(new_n260), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n541), .B1(new_n307), .B2(new_n481), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n298), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n464), .A2(new_n299), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n540), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n537), .B1(new_n533), .B2(new_n265), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n539), .B(new_n551), .C1(G169), .C2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n552), .A2(new_n443), .ZN(new_n555));
  AOI211_X1 g0355(.A(new_n440), .B(new_n537), .C1(new_n533), .C2(new_n265), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n321), .A2(G87), .A3(new_n462), .A4(new_n493), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n557), .A2(new_n549), .A3(new_n550), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT84), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n534), .A2(new_n538), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G200), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n552), .A2(G190), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n557), .A2(new_n549), .A3(new_n550), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT84), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(new_n553), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n256), .A2(G257), .A3(G1698), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n256), .A2(G250), .A3(new_n257), .ZN(new_n569));
  INV_X1    g0369(.A(G294), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n568), .B(new_n569), .C1(new_n267), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n506), .A2(new_n269), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n571), .A2(new_n265), .B1(new_n573), .B2(G264), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n509), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n428), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n425), .A3(new_n509), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n228), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n578));
  AND2_X1   g0378(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n579));
  NOR2_X1   g0379(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n256), .A2(new_n228), .A3(G87), .A4(new_n579), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT23), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n228), .B2(G107), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n454), .A2(KEYINPUT23), .A3(G20), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n267), .A2(new_n484), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n585), .A2(new_n586), .B1(new_n587), .B2(new_n228), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n582), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT24), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT24), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n582), .A2(new_n583), .A3(new_n588), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n321), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n299), .A2(new_n454), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT25), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n594), .B(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n494), .B2(new_n454), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n576), .B(new_n577), .C1(new_n593), .C2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n560), .A2(new_n567), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n454), .A2(KEYINPUT6), .A3(G97), .ZN(new_n600));
  AND2_X1   g0400(.A1(G97), .A2(G107), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n543), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n600), .B1(new_n602), .B2(KEYINPUT6), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(G20), .B1(G77), .B2(new_n313), .ZN(new_n604));
  OAI21_X1  g0404(.A(G107), .B1(new_n396), .B2(new_n397), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n321), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n300), .A2(G97), .A3(new_n493), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n462), .A2(G97), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(G257), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n509), .B1(new_n572), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(G244), .B(new_n257), .C1(new_n259), .C2(new_n260), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT4), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n257), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n480), .A4(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n612), .B1(new_n265), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G190), .ZN(new_n620));
  OAI21_X1  g0420(.A(G200), .B1(new_n619), .B2(KEYINPUT83), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n618), .A2(new_n265), .ZN(new_n622));
  INV_X1    g0422(.A(new_n612), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n622), .A2(new_n623), .A3(KEYINPUT83), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n610), .B(new_n620), .C1(new_n621), .C2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n593), .A2(new_n597), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n575), .A2(G200), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n574), .A2(G190), .A3(new_n509), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n609), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n604), .A2(new_n605), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n607), .B(new_n630), .C1(new_n631), .C2(new_n321), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n619), .A2(new_n425), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n622), .A2(new_n623), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n428), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n625), .A2(new_n629), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n599), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n479), .A2(new_n523), .A3(new_n530), .A4(new_n638), .ZN(new_n639));
  XOR2_X1   g0439(.A(new_n639), .B(KEYINPUT89), .Z(G372));
  NAND2_X1  g0440(.A1(new_n636), .A2(KEYINPUT92), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT91), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n534), .A2(KEYINPUT90), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n533), .A2(new_n644), .A3(new_n265), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n537), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n646), .B2(G169), .ZN(new_n647));
  INV_X1    g0447(.A(new_n645), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n644), .B1(new_n533), .B2(new_n265), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n538), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(KEYINPUT91), .A3(new_n428), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n539), .A2(new_n551), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n647), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n563), .B(new_n564), .C1(new_n646), .C2(new_n443), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT92), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n632), .A2(new_n635), .A3(new_n656), .A4(new_n633), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n641), .A2(new_n654), .A3(new_n655), .A4(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n565), .A2(new_n566), .A3(new_n553), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n566), .B1(new_n565), .B2(new_n553), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n661), .A2(new_n662), .A3(new_n636), .ZN(new_n663));
  XNOR2_X1  g0463(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n654), .ZN(new_n667));
  AND4_X1   g0467(.A1(new_n625), .A2(new_n629), .A3(new_n636), .A4(new_n655), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n515), .A2(new_n518), .A3(new_n521), .A4(new_n598), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n479), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n337), .A2(new_n335), .ZN(new_n673));
  INV_X1    g0473(.A(new_n331), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n451), .A2(new_n371), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n470), .B1(new_n380), .B2(new_n366), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n439), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n478), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n672), .A2(new_n679), .ZN(G369));
  NAND3_X1  g0480(.A1(new_n270), .A2(new_n228), .A3(G13), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT94), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g0485(.A(KEYINPUT95), .B(G343), .Z(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n523), .B(new_n530), .C1(new_n517), .C2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n522), .A2(new_n498), .A3(new_n687), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n598), .A2(new_n687), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n629), .B1(new_n626), .B2(new_n688), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n598), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n522), .A2(new_n688), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT96), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n695), .ZN(new_n700));
  INV_X1    g0500(.A(new_n693), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n697), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n235), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n544), .A2(G116), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n225), .B2(new_n706), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  AOI211_X1 g0510(.A(KEYINPUT29), .B(new_n687), .C1(new_n666), .C2(new_n670), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n658), .A2(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n670), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n712), .B1(new_n714), .B2(new_n688), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n638), .A2(new_n523), .A3(new_n530), .A4(new_n688), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n574), .A2(new_n552), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n520), .A2(new_n718), .A3(KEYINPUT30), .A4(new_n619), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n619), .A2(new_n574), .A3(new_n552), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n519), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n619), .A2(G179), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n650), .A3(new_n512), .A4(new_n575), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n719), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n725), .B2(new_n687), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n716), .B1(new_n717), .B2(new_n728), .ZN(new_n729));
  OR3_X1    g0529(.A1(new_n711), .A2(new_n715), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n710), .B1(new_n731), .B2(G1), .ZN(G364));
  NOR2_X1   g0532(.A1(new_n233), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n270), .B1(new_n733), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n705), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n227), .B1(G20), .B2(new_n428), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n228), .A2(new_n425), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G190), .ZN(new_n742));
  INV_X1    g0542(.A(G317), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT33), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n743), .A2(KEYINPUT33), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n440), .A2(G179), .A3(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n228), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n228), .A2(G179), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n746), .B1(new_n570), .B2(new_n748), .C1(new_n501), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G190), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n256), .B1(new_n754), .B2(G329), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n740), .A2(G190), .A3(new_n443), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G322), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n740), .A2(new_n752), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n755), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n741), .A2(new_n440), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G326), .ZN(new_n763));
  INV_X1    g0563(.A(G283), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n749), .A2(new_n440), .A3(G200), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n751), .A2(new_n761), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT100), .ZN(new_n768));
  INV_X1    g0568(.A(new_n760), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n757), .A2(G58), .B1(new_n769), .B2(G77), .ZN(new_n770));
  INV_X1    g0570(.A(new_n762), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n207), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT98), .ZN(new_n773));
  INV_X1    g0573(.A(new_n748), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G97), .A2(new_n774), .B1(new_n742), .B2(G68), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT99), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n753), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n750), .A2(new_n409), .ZN(new_n780));
  INV_X1    g0580(.A(new_n765), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n261), .B(new_n780), .C1(G107), .C2(new_n781), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n773), .A2(new_n776), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n739), .B1(new_n768), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G13), .A2(G33), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n738), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n235), .A2(new_n256), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT97), .Z(new_n790));
  AOI22_X1  g0590(.A1(new_n790), .A2(G355), .B1(new_n484), .B2(new_n704), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n704), .A2(new_n256), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n276), .A2(new_n278), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n792), .B1(new_n254), .B2(new_n275), .C1(new_n225), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n737), .B(new_n784), .C1(new_n788), .C2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n787), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n691), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT101), .ZN(new_n800));
  INV_X1    g0600(.A(new_n692), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n736), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(G330), .B2(new_n691), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n800), .A2(new_n803), .ZN(G396));
  NAND2_X1  g0604(.A1(new_n473), .A2(new_n688), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n671), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n671), .A2(new_n688), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n469), .A2(new_n687), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n472), .A2(new_n471), .B1(new_n467), .B2(new_n687), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n470), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n807), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n729), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n736), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n738), .A2(new_n785), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n737), .B1(new_n350), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n256), .B1(new_n754), .B2(G311), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n821), .B1(new_n484), .B2(new_n760), .C1(new_n570), .C2(new_n756), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n762), .A2(G303), .B1(new_n781), .B2(G87), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n454), .B2(new_n750), .ZN(new_n824));
  INV_X1    g0624(.A(new_n742), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n825), .A2(new_n764), .B1(new_n481), .B2(new_n748), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n822), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n256), .B1(new_n753), .B2(new_n828), .C1(new_n207), .C2(new_n750), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n748), .A2(new_n202), .B1(new_n765), .B2(new_n203), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n757), .A2(G143), .B1(new_n769), .B2(G159), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G137), .A2(new_n762), .B1(new_n742), .B2(G150), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT102), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(KEYINPUT102), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n829), .B(new_n830), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n827), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n820), .B1(new_n739), .B2(new_n840), .C1(new_n814), .C2(new_n786), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n818), .A2(new_n841), .ZN(G384));
  NOR2_X1   g0642(.A1(new_n733), .A2(new_n270), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n805), .B1(new_n666), .B2(new_n670), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n844), .A2(new_n810), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n687), .A2(new_n366), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n381), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n366), .B(new_n687), .C1(new_n380), .C2(new_n372), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT103), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT103), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n849), .B(new_n852), .C1(new_n844), .C2(new_n810), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n436), .A2(new_n438), .A3(new_n450), .A4(new_n447), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n402), .A2(new_n300), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n855), .A2(new_n404), .B1(new_n462), .B2(new_n324), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT104), .B1(new_n389), .B2(new_n394), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT104), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n398), .A2(new_n858), .A3(new_n399), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n857), .A2(new_n859), .A3(new_n382), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n389), .A2(new_n394), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n321), .B1(new_n861), .B2(KEYINPUT16), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n856), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(new_n685), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n854), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT82), .B1(new_n427), .B2(new_n430), .ZN(new_n866));
  INV_X1    g0666(.A(new_n434), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n863), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n448), .B1(new_n863), .B2(new_n685), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n685), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n408), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n435), .A2(new_n872), .A3(new_n873), .A4(new_n448), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n865), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n865), .A2(new_n875), .A3(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n851), .A2(new_n853), .A3(new_n880), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n439), .A2(new_n871), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n380), .A2(new_n366), .A3(new_n688), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n878), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n867), .A2(new_n866), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n446), .B1(new_n886), .B2(new_n408), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n887), .A2(KEYINPUT105), .A3(new_n873), .A4(new_n872), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT105), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n874), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n435), .A2(new_n448), .A3(new_n872), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n888), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n854), .A2(new_n408), .A3(new_n871), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n879), .A2(KEYINPUT106), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT106), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n865), .A2(new_n875), .A3(new_n897), .A4(KEYINPUT38), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n895), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n884), .B(new_n885), .C1(new_n899), .C2(KEYINPUT39), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n881), .A2(new_n882), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n479), .B1(new_n711), .B2(new_n715), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n902), .A2(new_n679), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n901), .B(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT107), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n717), .A2(new_n728), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n813), .B1(new_n847), .B2(new_n848), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT40), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n905), .B1(new_n899), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n893), .A2(new_n894), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n877), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n854), .A2(new_n864), .B1(new_n870), .B2(new_n874), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n897), .B1(new_n912), .B2(KEYINPUT38), .ZN(new_n913));
  AND4_X1   g0713(.A1(new_n897), .A2(new_n865), .A3(new_n875), .A4(KEYINPUT38), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n906), .A2(KEYINPUT40), .A3(new_n907), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(KEYINPUT107), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n880), .A2(new_n906), .A3(new_n907), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n909), .A2(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n479), .A2(new_n906), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n716), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n843), .B1(new_n904), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n904), .B2(new_n923), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n603), .A2(KEYINPUT35), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n603), .A2(KEYINPUT35), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n926), .A2(G116), .A3(new_n229), .A4(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT36), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n226), .A2(G77), .A3(new_n390), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(G50), .B2(new_n203), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(G1), .A3(new_n233), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n925), .A2(new_n929), .A3(new_n932), .ZN(G367));
  OAI211_X1 g0733(.A(new_n625), .B(new_n636), .C1(new_n610), .C2(new_n688), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n636), .A2(new_n688), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n699), .A2(new_n695), .A3(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n937), .A2(KEYINPUT42), .ZN(new_n938));
  INV_X1    g0738(.A(new_n598), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n625), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n687), .B1(new_n940), .B2(new_n636), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n937), .B2(KEYINPUT42), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n687), .A2(new_n558), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n654), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n654), .A2(new_n655), .A3(new_n944), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n943), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n938), .A2(new_n942), .A3(new_n949), .A4(new_n948), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n697), .ZN(new_n955));
  INV_X1    g0755(.A(new_n936), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n954), .B(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n705), .B(KEYINPUT41), .Z(new_n959));
  AOI21_X1  g0759(.A(new_n936), .B1(new_n700), .B2(new_n701), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT44), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n960), .B(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n702), .B2(new_n956), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n700), .A2(new_n701), .A3(new_n936), .A4(new_n963), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n697), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT96), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n698), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n696), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n700), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(new_n801), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n731), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n965), .A2(new_n966), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n702), .A2(new_n956), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n961), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n702), .A2(KEYINPUT44), .A3(new_n956), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n976), .A2(new_n980), .A3(new_n955), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n968), .A2(new_n975), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n959), .B1(new_n982), .B2(new_n731), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n958), .B1(new_n983), .B2(new_n735), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n792), .A2(new_n246), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n788), .B1(new_n235), .B2(new_n464), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n825), .A2(new_n570), .B1(new_n765), .B2(new_n481), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n771), .A2(new_n759), .B1(new_n454), .B2(new_n748), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n261), .B1(new_n760), .B2(new_n764), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n756), .A2(new_n501), .B1(new_n753), .B2(new_n743), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n750), .A2(new_n484), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n990), .B(new_n991), .C1(KEYINPUT46), .C2(new_n992), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n989), .B(new_n993), .C1(KEYINPUT46), .C2(new_n992), .ZN(new_n994));
  INV_X1    g0794(.A(G150), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n748), .A2(new_n203), .B1(new_n756), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT109), .ZN(new_n997));
  AOI22_X1  g0797(.A1(G143), .A2(new_n762), .B1(new_n742), .B2(G159), .ZN(new_n998));
  INV_X1    g0798(.A(G137), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n256), .B1(new_n753), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G50), .B2(new_n769), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n765), .A2(new_n350), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n750), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1002), .B1(G58), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n998), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n994), .B1(new_n997), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT47), .Z(new_n1007));
  OAI221_X1 g0807(.A(new_n736), .B1(new_n985), .B2(new_n986), .C1(new_n1007), .C2(new_n739), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT110), .Z(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n798), .B2(new_n947), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n984), .A2(new_n1010), .ZN(G387));
  NAND2_X1  g0811(.A1(new_n973), .A2(new_n735), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n756), .A2(new_n207), .B1(new_n760), .B2(new_n203), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n261), .B(new_n1013), .C1(G150), .C2(new_n754), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n762), .A2(G159), .B1(new_n781), .B2(G97), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n748), .A2(new_n464), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G77), .B2(new_n1003), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n742), .A2(new_n324), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n756), .A2(new_n743), .B1(new_n760), .B2(new_n501), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT111), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(KEYINPUT111), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G311), .A2(new_n742), .B1(new_n762), .B2(G322), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n748), .A2(new_n764), .B1(new_n750), .B2(new_n570), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1026), .A2(KEYINPUT49), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n256), .B1(new_n754), .B2(G326), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(new_n484), .C2(new_n765), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT49), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1019), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT112), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n739), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n1034), .B2(new_n1033), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n696), .A2(new_n787), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n790), .B1(G116), .B2(new_n544), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n243), .A2(new_n793), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n305), .A2(G50), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT50), .Z(new_n1041));
  OAI211_X1 g0841(.A(new_n707), .B(new_n275), .C1(new_n203), .C2(new_n350), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n792), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1038), .B1(G107), .B2(new_n235), .C1(new_n1039), .C2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n737), .B1(new_n1044), .B2(new_n788), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1036), .A2(new_n1037), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n974), .A2(new_n705), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n973), .A2(new_n731), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1012), .B(new_n1046), .C1(new_n1047), .C2(new_n1048), .ZN(G393));
  NAND3_X1  g0849(.A1(new_n968), .A2(new_n981), .A3(new_n735), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n788), .B1(new_n481), .B2(new_n235), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n251), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1051), .B1(new_n1052), .B2(new_n792), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1053), .A2(new_n737), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G150), .A2(new_n762), .B1(new_n757), .B2(G159), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT113), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT51), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n261), .B1(new_n754), .B2(G143), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n203), .B2(new_n750), .C1(new_n409), .C2(new_n765), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT114), .Z(new_n1060));
  NOR2_X1   g0860(.A1(new_n748), .A2(new_n350), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n305), .B2(new_n760), .C1(new_n207), .C2(new_n825), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n1057), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n771), .A2(new_n743), .B1(new_n759), .B2(new_n756), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT52), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n825), .A2(new_n501), .B1(new_n765), .B2(new_n454), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n256), .B1(new_n754), .B2(G322), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n570), .B2(new_n760), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n748), .A2(new_n484), .B1(new_n750), .B2(new_n764), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1064), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1054), .B1(new_n936), .B2(new_n798), .C1(new_n1072), .C2(new_n739), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n982), .A2(new_n705), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n975), .B1(new_n968), .B2(new_n981), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1050), .B(new_n1073), .C1(new_n1074), .C2(new_n1075), .ZN(G390));
  INV_X1    g0876(.A(new_n819), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1062), .B1(new_n771), .B2(new_n764), .C1(new_n454), .C2(new_n825), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n757), .A2(G116), .B1(new_n754), .B2(G294), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1079), .B(new_n261), .C1(new_n481), .C2(new_n760), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n765), .A2(new_n203), .ZN(new_n1081));
  NOR4_X1   g0881(.A1(new_n1078), .A2(new_n1080), .A3(new_n780), .A4(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(KEYINPUT54), .B(G143), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n748), .A2(new_n777), .B1(new_n760), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G137), .B2(new_n742), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT117), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n256), .B1(new_n765), .B2(new_n207), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT118), .Z(new_n1088));
  AOI22_X1  g0888(.A1(new_n757), .A2(G132), .B1(new_n754), .B2(G125), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1090));
  OR3_X1    g0890(.A1(new_n1090), .A2(new_n750), .A3(new_n995), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n750), .B2(new_n995), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n762), .A2(G128), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1088), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1082), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n736), .B1(new_n324), .B2(new_n1077), .C1(new_n1096), .C2(new_n739), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n878), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT39), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n915), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1097), .B1(new_n1101), .B2(new_n785), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n847), .A2(KEYINPUT115), .A3(new_n848), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT115), .B1(new_n847), .B2(new_n848), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n687), .B1(new_n713), .B2(new_n670), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n812), .A2(new_n470), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n810), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n915), .B(new_n883), .C1(new_n1107), .C2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n807), .A2(new_n811), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n884), .B1(new_n1113), .B2(new_n849), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1112), .B1(new_n1100), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n729), .A2(new_n849), .A3(new_n814), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1112), .B(new_n1116), .C1(new_n1100), .C2(new_n1114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1103), .B1(new_n1120), .B2(new_n734), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n479), .A2(KEYINPUT116), .A3(new_n729), .ZN(new_n1122));
  AOI21_X1  g0922(.A(KEYINPUT116), .B1(new_n479), .B2(new_n729), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n902), .B(new_n679), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n849), .B1(new_n729), .B2(new_n814), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1113), .B1(new_n1117), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n729), .A2(new_n814), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1111), .B(new_n1116), .C1(new_n1128), .C2(new_n1106), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1124), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n706), .B1(new_n1120), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1118), .A2(new_n1130), .A3(new_n1119), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1121), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(G378));
  NAND3_X1  g0935(.A1(new_n881), .A2(new_n882), .A3(new_n900), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n909), .A2(new_n917), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n716), .B1(new_n919), .B2(new_n918), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n478), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n476), .A2(new_n871), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n675), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n675), .B2(new_n1141), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1145), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n1143), .A3(new_n1139), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1137), .A2(new_n1138), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1149), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1136), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n899), .A2(new_n905), .A3(new_n908), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT107), .B1(new_n915), .B2(new_n916), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1138), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1149), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1137), .A2(new_n1138), .A3(new_n1149), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n901), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n734), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1156), .A2(new_n785), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n736), .B1(G50), .B2(new_n1077), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n261), .B2(new_n268), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n771), .A2(new_n484), .B1(new_n765), .B2(new_n202), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G97), .B2(new_n742), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G41), .B(new_n256), .C1(new_n754), .C2(G283), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n757), .A2(G107), .B1(new_n769), .B2(new_n465), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n774), .A2(G68), .B1(new_n1003), .B2(G77), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT58), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1164), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n762), .A2(G125), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n825), .B2(new_n828), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n757), .A2(G128), .B1(new_n769), .B2(G137), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n750), .B2(new_n1083), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1174), .B(new_n1176), .C1(G150), .C2(new_n774), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT120), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G33), .B(G41), .C1(new_n754), .C2(G124), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(new_n777), .C2(new_n765), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1178), .A2(KEYINPUT120), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1172), .B1(new_n1171), .B2(new_n1170), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1162), .B1(new_n1183), .B2(new_n738), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1161), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1160), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1152), .A2(new_n1159), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1124), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1133), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT57), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n705), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1159), .A2(new_n1152), .B1(new_n1133), .B2(new_n1189), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT57), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1187), .B1(new_n1193), .B2(new_n1195), .ZN(G375));
  OAI22_X1  g0996(.A1(new_n825), .A2(new_n1083), .B1(new_n999), .B2(new_n756), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n202), .A2(new_n765), .B1(new_n750), .B2(new_n777), .ZN(new_n1198));
  INV_X1    g0998(.A(G128), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n256), .B1(new_n753), .B2(new_n1199), .C1(new_n995), .C2(new_n760), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(G50), .C2(new_n774), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT121), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1197), .B(new_n1202), .C1(G132), .C2(new_n762), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G116), .A2(new_n742), .B1(new_n762), .B2(G294), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n481), .B2(new_n750), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n256), .B1(new_n754), .B2(G303), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n454), .B2(new_n760), .C1(new_n764), .C2(new_n756), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1205), .A2(new_n1207), .A3(new_n1002), .A4(new_n1016), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n738), .B1(new_n1203), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n737), .B1(new_n203), .B2(new_n819), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(new_n1106), .C2(new_n786), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1213), .B2(new_n734), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n959), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1131), .A2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1189), .A2(new_n1212), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1215), .B1(new_n1217), .B2(new_n1218), .ZN(G381));
  NOR3_X1   g1019(.A1(G378), .A2(G381), .A3(G390), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT122), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n1223), .A2(G387), .A3(G375), .ZN(G407));
  NAND2_X1  g1024(.A1(new_n686), .A2(G213), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1134), .A2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(G375), .C2(new_n1227), .ZN(G409));
  INV_X1    g1028(.A(G390), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(G387), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT125), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n984), .A2(G390), .A3(new_n1010), .ZN(new_n1232));
  XOR2_X1   g1032(.A(G393), .B(G396), .Z(new_n1233));
  NAND4_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(KEYINPUT125), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1236), .A2(new_n1233), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1150), .A2(new_n1151), .A3(new_n1136), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n901), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n735), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT123), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1243), .A3(new_n1185), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT123), .B1(new_n1160), .B2(new_n1186), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1194), .A2(new_n1216), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1134), .ZN(new_n1248));
  OAI211_X1 g1048(.A(G378), .B(new_n1187), .C1(new_n1193), .C2(new_n1195), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT62), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT60), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1252), .B1(new_n1218), .B2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(KEYINPUT124), .B(KEYINPUT60), .C1(new_n1189), .C2(new_n1212), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1130), .A2(new_n706), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(G384), .A3(new_n1215), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G384), .B1(new_n1258), .B2(new_n1215), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1250), .A2(new_n1251), .A3(new_n1225), .A4(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1226), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1265));
  OAI211_X1 g1065(.A(G2897), .B(new_n1226), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1261), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1226), .A2(G2897), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n1259), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1263), .B(new_n1264), .C1(new_n1265), .C2(new_n1270), .ZN(new_n1271));
  XOR2_X1   g1071(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1265), .B2(new_n1262), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1239), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1270), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1265), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT61), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1265), .A2(new_n1262), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT63), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1265), .A2(KEYINPUT63), .A3(new_n1262), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1277), .A2(new_n1280), .A3(new_n1238), .A4(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1274), .A2(new_n1282), .ZN(G405));
  NAND2_X1  g1083(.A1(new_n1262), .A2(KEYINPUT127), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1262), .A2(KEYINPUT127), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G375), .A2(new_n1134), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1287), .B1(new_n1249), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1236), .A2(new_n1233), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n1234), .A3(new_n1284), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1286), .A2(new_n1289), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1289), .B1(new_n1286), .B2(new_n1293), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(G402));
endmodule


