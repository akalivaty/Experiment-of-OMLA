//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224, new_n1226, new_n1227,
    new_n1228, new_n1229;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT64), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n452), .A2(G2106), .B1(KEYINPUT65), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n459), .B1(KEYINPUT65), .B2(new_n458), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G137), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n462), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g050(.A(KEYINPUT67), .B(new_n470), .C1(new_n475), .C2(new_n464), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n478), .B1(new_n467), .B2(new_n468), .ZN(new_n479));
  AND2_X1   g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  OAI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n475), .A2(G2105), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(G136), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT3), .B(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n489), .B1(new_n492), .B2(G124), .ZN(new_n493));
  INV_X1    g068(.A(G124), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n491), .A2(KEYINPUT68), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n488), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n463), .A2(KEYINPUT69), .A3(G138), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n475), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n490), .A2(G126), .A3(G2105), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n463), .A2(KEYINPUT69), .A3(G138), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n490), .A2(KEYINPUT4), .A3(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n500), .A2(new_n501), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT70), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT70), .A2(G651), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT6), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n510), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n510), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n511), .A2(new_n512), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n516), .A2(G88), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n513), .B2(new_n515), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n522), .A2(new_n525), .ZN(G166));
  INV_X1    g101(.A(KEYINPUT5), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(new_n523), .ZN(new_n528));
  NAND2_X1  g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n516), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n524), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(new_n516), .A2(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n524), .A2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n510), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(new_n521), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(G171));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n510), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n524), .A2(G43), .B1(new_n549), .B2(new_n521), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n516), .A2(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT6), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT70), .ZN(new_n561));
  INV_X1    g136(.A(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(KEYINPUT70), .A2(G651), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(G543), .B1(new_n565), .B2(new_n514), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI211_X1 g142(.A(KEYINPUT72), .B(new_n559), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n510), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n516), .A2(G91), .B1(new_n571), .B2(G651), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT72), .B1(new_n566), .B2(new_n567), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n524), .A2(new_n575), .A3(G53), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(KEYINPUT9), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G299));
  NAND3_X1  g153(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT73), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(G301));
  NAND2_X1  g156(.A1(new_n522), .A2(new_n525), .ZN(G303));
  NAND2_X1  g157(.A1(new_n524), .A2(G49), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n516), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  OAI211_X1 g161(.A(G48), .B(G543), .C1(new_n565), .C2(new_n514), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n530), .B1(new_n565), .B2(new_n514), .ZN(new_n588));
  INV_X1    g163(.A(G86), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(G61), .B1(new_n508), .B2(new_n509), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(KEYINPUT74), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n595), .B(G61), .C1(new_n508), .C2(new_n509), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n520), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n510), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n521), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT75), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(G47), .A2(new_n524), .B1(new_n516), .B2(G85), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(G301), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n510), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n524), .A2(G54), .B1(new_n612), .B2(G651), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n516), .A2(KEYINPUT10), .A3(G92), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(KEYINPUT10), .B1(new_n516), .B2(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT76), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  INV_X1    g195(.A(G92), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n588), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n614), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n623), .A2(KEYINPUT76), .A3(new_n613), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n609), .B1(new_n608), .B2(new_n625), .ZN(G284));
  AOI21_X1  g201(.A(new_n609), .B1(new_n608), .B2(new_n625), .ZN(G321));
  NAND2_X1  g202(.A1(G299), .A2(new_n608), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n608), .B2(G168), .ZN(G280));
  XNOR2_X1  g204(.A(G280), .B(KEYINPUT77), .ZN(G297));
  XOR2_X1   g205(.A(KEYINPUT78), .B(G559), .Z(new_n631));
  OAI21_X1  g206(.A(new_n625), .B1(G860), .B2(new_n631), .ZN(G148));
  NAND2_X1  g207(.A1(new_n552), .A2(new_n608), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n625), .A2(new_n631), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n633), .B1(new_n635), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g212(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n638));
  NOR3_X1   g213(.A1(new_n465), .A2(new_n466), .A3(G2105), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n641), .A2(G2100), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT80), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n487), .A2(G135), .ZN(new_n644));
  OR2_X1    g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n645), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n646));
  INV_X1    g221(.A(G123), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n646), .C1(new_n647), .C2(new_n491), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2096), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(G2100), .B2(new_n641), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n643), .A2(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2443), .B(G2446), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT81), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(G14), .B1(new_n662), .B2(new_n664), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2100), .ZN(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G2096), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n685), .A2(new_n688), .A3(new_n692), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT83), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT84), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n699), .B(new_n702), .ZN(G229));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G6), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n598), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT86), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT32), .B(G1981), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n704), .A2(G23), .ZN(new_n712));
  INV_X1    g287(.A(G288), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n704), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT33), .B(G1976), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n704), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n704), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT87), .B(G1971), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  AND4_X1   g295(.A1(new_n710), .A2(new_n711), .A3(new_n716), .A4(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT34), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  MUX2_X1   g299(.A(G24), .B(G290), .S(G16), .Z(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT85), .B(G1986), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n492), .A2(G119), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n487), .A2(G131), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n463), .A2(G107), .ZN(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  MUX2_X1   g307(.A(G25), .B(new_n732), .S(G29), .Z(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n727), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n723), .A2(new_n724), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT88), .B(KEYINPUT36), .Z(new_n739));
  AND2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(G168), .A2(G16), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G16), .B2(G21), .ZN(new_n744));
  INV_X1    g319(.A(G1966), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G1961), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n579), .A2(G16), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n704), .A2(G5), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI22_X1  g325(.A1(new_n744), .A2(new_n745), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G35), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G162), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT29), .ZN(new_n754));
  INV_X1    g329(.A(G2090), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n746), .B(new_n751), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G32), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n487), .A2(G141), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT94), .ZN(new_n762));
  AND3_X1   g337(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT26), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n763), .B(new_n765), .C1(new_n492), .C2(G129), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n760), .B1(new_n768), .B2(new_n759), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT27), .B(G1996), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n750), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(G1961), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  INV_X1    g349(.A(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n774), .B2(new_n775), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G160), .B2(new_n759), .ZN(new_n778));
  INV_X1    g353(.A(G2084), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(G164), .A2(G29), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G27), .B2(G29), .ZN(new_n782));
  INV_X1    g357(.A(G2078), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT30), .B(G28), .ZN(new_n785));
  OR2_X1    g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  NAND2_X1  g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n785), .A2(new_n759), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n648), .B2(new_n759), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n780), .B(new_n790), .C1(new_n783), .C2(new_n782), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n773), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n487), .A2(G139), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT91), .ZN(new_n794));
  NAND2_X1  g369(.A1(G115), .A2(G2104), .ZN(new_n795));
  INV_X1    g370(.A(G127), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n475), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT25), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n797), .A2(G2105), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n794), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT92), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n794), .A2(KEYINPUT92), .A3(new_n802), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(G29), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G33), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(G29), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT93), .B(G2072), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n758), .A2(new_n792), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n704), .A2(G4), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n625), .B2(new_n704), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(G1348), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(G1348), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n704), .A2(G19), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n553), .B2(new_n704), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(G1341), .Z(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n759), .A2(G26), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n492), .A2(G128), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n487), .A2(G140), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n463), .A2(G116), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n825), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n824), .B1(new_n829), .B2(G29), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G2067), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n817), .A2(new_n818), .A3(new_n821), .A4(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(KEYINPUT90), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(KEYINPUT90), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n704), .A2(G20), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT23), .Z(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G299), .B2(G16), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G1956), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n814), .A2(new_n833), .A3(new_n834), .A4(new_n838), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n740), .A2(new_n742), .A3(new_n839), .ZN(G311));
  OR3_X1    g415(.A1(new_n740), .A2(new_n742), .A3(new_n839), .ZN(G150));
  NAND2_X1  g416(.A1(new_n625), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT95), .B(G93), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n516), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n524), .A2(G55), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n530), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n845), .B(new_n846), .C1(new_n520), .C2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n552), .B(new_n848), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n843), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n852));
  AOI21_X1  g427(.A(G860), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n848), .A2(G860), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT96), .B(KEYINPUT37), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(G145));
  AOI21_X1  g433(.A(new_n768), .B1(new_n805), .B2(new_n807), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n805), .A2(new_n768), .A3(new_n807), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n492), .A2(G130), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n487), .A2(G142), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n463), .A2(G118), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n862), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n732), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n860), .A2(new_n861), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n861), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n867), .B1(new_n870), .B2(new_n859), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n829), .B(new_n506), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n640), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(G162), .B(new_n482), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(new_n648), .Z(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n869), .A2(new_n871), .A3(new_n874), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n876), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n876), .A2(new_n880), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT97), .B1(new_n884), .B2(new_n878), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT97), .ZN(new_n886));
  AOI211_X1 g461(.A(new_n886), .B(new_n879), .C1(new_n876), .C2(new_n880), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n883), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(G395));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n605), .A2(new_n713), .A3(new_n606), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n713), .B1(new_n605), .B2(new_n606), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(G290), .A2(G288), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(KEYINPUT100), .A3(new_n892), .ZN(new_n897));
  XNOR2_X1  g472(.A(G166), .B(new_n598), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT100), .B1(new_n896), .B2(new_n892), .ZN(new_n900));
  INV_X1    g475(.A(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT102), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n906));
  AOI211_X1 g481(.A(new_n906), .B(KEYINPUT42), .C1(new_n899), .C2(new_n902), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n635), .A2(new_n850), .ZN(new_n909));
  NAND2_X1  g484(.A1(G299), .A2(new_n617), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n573), .A2(new_n577), .A3(new_n623), .A4(new_n613), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n634), .A2(new_n849), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT99), .B1(new_n912), .B2(KEYINPUT41), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(KEYINPUT41), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n910), .A2(new_n917), .A3(new_n911), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n915), .B1(new_n919), .B2(KEYINPUT99), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n909), .A2(new_n913), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n914), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n903), .A2(KEYINPUT101), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n899), .A2(new_n924), .A3(new_n902), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(KEYINPUT42), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n908), .A2(new_n922), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n922), .B1(new_n908), .B2(new_n926), .ZN(new_n929));
  OAI21_X1  g504(.A(G868), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n848), .A2(new_n608), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(G295));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n933), .A3(new_n931), .ZN(new_n934));
  INV_X1    g509(.A(new_n907), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n903), .A2(new_n904), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n906), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n926), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  MUX2_X1   g513(.A(new_n912), .B(new_n920), .S(new_n921), .Z(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n608), .B1(new_n940), .B2(new_n927), .ZN(new_n941));
  INV_X1    g516(.A(new_n931), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT103), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n934), .A2(new_n943), .ZN(G331));
  INV_X1    g519(.A(new_n925), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n924), .B1(new_n899), .B2(new_n902), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(G286), .A2(new_n579), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n579), .B(KEYINPUT73), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n949), .B2(G168), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n950), .A2(new_n849), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(new_n912), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(G168), .ZN(new_n953));
  INV_X1    g528(.A(new_n948), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n849), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n950), .A2(KEYINPUT105), .A3(new_n849), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n951), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n947), .B(new_n956), .C1(new_n920), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n923), .A2(new_n925), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n920), .A2(new_n960), .ZN(new_n963));
  INV_X1    g538(.A(new_n956), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n961), .A2(new_n965), .A3(new_n966), .A4(new_n882), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n958), .A2(new_n959), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n952), .ZN(new_n969));
  INV_X1    g544(.A(new_n955), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n919), .B1(new_n970), .B2(new_n951), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G37), .B1(new_n972), .B2(new_n962), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n961), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(KEYINPUT44), .B(new_n967), .C1(new_n974), .C2(new_n966), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n961), .A2(new_n965), .A3(new_n882), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n963), .A2(new_n964), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT43), .B1(new_n977), .B2(new_n947), .ZN(new_n978));
  AOI22_X1  g553(.A1(KEYINPUT43), .A2(new_n976), .B1(new_n978), .B2(new_n973), .ZN(new_n979));
  XOR2_X1   g554(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n980));
  OAI21_X1  g555(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(G397));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n506), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n472), .A2(new_n481), .A3(G40), .A4(new_n476), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  OR3_X1    g563(.A1(new_n988), .A2(G1986), .A3(G290), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(G290), .A3(G1986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT106), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n987), .A2(G1996), .A3(new_n767), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT107), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n767), .A2(G1996), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n829), .B(G2067), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n987), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n732), .B(new_n734), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n999), .A2(KEYINPUT108), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(KEYINPUT108), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n987), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n992), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1971), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n984), .A2(G1384), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n506), .A2(new_n1006), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n481), .A2(G40), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n477), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT45), .B1(new_n506), .B2(new_n982), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1005), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT109), .ZN(new_n1012));
  INV_X1    g587(.A(new_n986), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n506), .A2(new_n982), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT50), .B1(new_n506), .B2(new_n982), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n755), .B(new_n1013), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n506), .A2(new_n982), .A3(new_n1014), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n475), .A2(new_n498), .A3(new_n499), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT4), .B1(new_n490), .B2(new_n502), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n501), .A2(new_n505), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1384), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1020), .B1(new_n1025), .B2(KEYINPUT50), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1026), .A2(KEYINPUT111), .A3(new_n755), .A4(new_n1013), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(new_n1005), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1012), .A2(new_n1019), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G303), .A2(G8), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT55), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1030), .A2(G8), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(G8), .B1(new_n983), .B2(new_n986), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n713), .A2(G1976), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G288), .A2(new_n1038), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT52), .B1(new_n1035), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(G1981), .B1(new_n590), .B2(new_n597), .ZN(new_n1045));
  INV_X1    g620(.A(G61), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n528), .B2(new_n529), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n591), .B1(new_n1047), .B2(new_n595), .ZN(new_n1048));
  INV_X1    g623(.A(new_n596), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n521), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n516), .A2(G86), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n587), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1045), .A2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1045), .A2(new_n1053), .A3(KEYINPUT49), .ZN(new_n1057));
  AND4_X1   g632(.A1(KEYINPUT113), .A2(new_n1056), .A3(new_n1057), .A4(new_n1036), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1035), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT113), .B1(new_n1059), .B2(new_n1057), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1044), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1034), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n985), .A2(new_n783), .A3(new_n1013), .A4(new_n1007), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n747), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n986), .B1(new_n506), .B2(new_n1006), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(KEYINPUT53), .A3(new_n783), .A4(new_n985), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT123), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1065), .A2(new_n1067), .A3(G301), .A4(new_n1069), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1073), .A2(KEYINPUT54), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1075), .A3(G171), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1014), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1078), .B(new_n1013), .C1(new_n1025), .C2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n506), .B2(new_n982), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT115), .B1(new_n1081), .B2(new_n986), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n983), .A2(KEYINPUT50), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1011), .B1(new_n1085), .B2(G2090), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G8), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1032), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1070), .A2(new_n949), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1073), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1062), .A2(new_n1077), .A3(new_n1088), .A4(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n745), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n779), .B(new_n1013), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1094), .A2(new_n1095), .A3(G168), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  AND2_X1   g672(.A1(KEYINPUT121), .A2(G8), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(G8), .A3(G286), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1097), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT122), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT51), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1101), .A4(new_n1099), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT124), .B1(new_n1093), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1077), .A2(new_n1092), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1059), .A2(new_n1057), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT113), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1059), .A2(KEYINPUT113), .A3(new_n1057), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1043), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1030), .A2(G8), .A3(new_n1033), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1118), .A2(new_n1088), .A3(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1112), .A2(new_n1113), .A3(new_n1109), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1956), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1085), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n573), .A2(new_n1124), .A3(new_n577), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1124), .B1(new_n573), .B2(new_n577), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT56), .B(G2072), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1068), .A2(new_n985), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1123), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n1131));
  INV_X1    g706(.A(new_n625), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n983), .A2(new_n986), .A3(G2067), .ZN(new_n1133));
  INV_X1    g708(.A(G1348), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n1066), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1131), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(G1348), .B1(new_n1026), .B2(new_n1013), .ZN(new_n1137));
  OAI211_X1 g712(.A(KEYINPUT117), .B(new_n625), .C1(new_n1137), .C2(new_n1133), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1127), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1130), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT118), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1143), .B(new_n1130), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT61), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n986), .B1(new_n983), .B2(new_n1014), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1083), .B1(new_n1147), .B2(new_n1078), .ZN(new_n1148));
  AOI21_X1  g723(.A(G1956), .B1(new_n1148), .B2(new_n1082), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1129), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1149), .A2(new_n1150), .B1(new_n1126), .B2(new_n1125), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1151), .A2(new_n1130), .A3(KEYINPUT120), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n619), .A2(new_n1154), .A3(new_n624), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1135), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n625), .A2(KEYINPUT60), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1151), .A2(new_n1130), .A3(KEYINPUT61), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1009), .A2(G1996), .A3(new_n1010), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n983), .A2(new_n986), .ZN(new_n1163));
  XOR2_X1   g738(.A(KEYINPUT58), .B(G1341), .Z(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1161), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(G1996), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1068), .A2(new_n1168), .A3(new_n985), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1169), .B(KEYINPUT119), .C1(new_n1163), .C2(new_n1165), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1160), .B1(new_n1171), .B2(new_n553), .ZN(new_n1172));
  AOI211_X1 g747(.A(KEYINPUT59), .B(new_n552), .C1(new_n1167), .C2(new_n1170), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1158), .B(new_n1159), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1142), .B(new_n1144), .C1(new_n1153), .C2(new_n1174), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1111), .A2(new_n1121), .A3(new_n1175), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1038), .B(new_n713), .C1(new_n1058), .C2(new_n1060), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1035), .B1(new_n1177), .B2(new_n1053), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1061), .A2(new_n1119), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT114), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n713), .A2(new_n1038), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1181), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1053), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1036), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT114), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1118), .A2(new_n1034), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1180), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1100), .A2(G8), .A3(G168), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT116), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1191), .A2(new_n1088), .A3(new_n1119), .A4(new_n1118), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1030), .A2(G8), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1032), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1062), .A2(KEYINPUT63), .A3(new_n1191), .A4(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1089), .ZN(new_n1199));
  AND4_X1   g774(.A1(new_n1088), .A2(new_n1118), .A3(new_n1119), .A4(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1104), .A2(new_n1201), .A3(new_n1108), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1201), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1203));
  OAI211_X1 g778(.A(new_n1200), .B(new_n1202), .C1(new_n1203), .C2(KEYINPUT125), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1203), .A2(KEYINPUT125), .ZN(new_n1205));
  OAI211_X1 g780(.A(new_n1188), .B(new_n1198), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1004), .B1(new_n1176), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g782(.A(KEYINPUT46), .B1(new_n987), .B2(new_n1168), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1208), .B(KEYINPUT126), .Z(new_n1209));
  NAND3_X1  g784(.A1(new_n987), .A2(KEYINPUT46), .A3(new_n1168), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT127), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n987), .B1(new_n996), .B2(new_n767), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1209), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  XOR2_X1   g788(.A(new_n1213), .B(KEYINPUT47), .Z(new_n1214));
  NOR2_X1   g789(.A1(new_n829), .A2(G2067), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n732), .A2(new_n735), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1215), .B1(new_n998), .B2(new_n1216), .ZN(new_n1217));
  XOR2_X1   g792(.A(new_n989), .B(KEYINPUT48), .Z(new_n1218));
  OAI22_X1  g793(.A1(new_n1217), .A2(new_n988), .B1(new_n1003), .B2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g794(.A1(new_n1214), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1207), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g796(.A1(G229), .A2(new_n460), .A3(G227), .ZN(new_n1223));
  NAND3_X1  g797(.A1(new_n888), .A2(new_n670), .A3(new_n1223), .ZN(new_n1224));
  NOR2_X1   g798(.A1(new_n1224), .A2(new_n979), .ZN(G308));
  INV_X1    g799(.A(new_n1223), .ZN(new_n1226));
  AOI21_X1  g800(.A(new_n1226), .B1(new_n667), .B2(new_n669), .ZN(new_n1227));
  AND2_X1   g801(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n1228));
  AND2_X1   g802(.A1(new_n978), .A2(new_n973), .ZN(new_n1229));
  OAI211_X1 g803(.A(new_n888), .B(new_n1227), .C1(new_n1228), .C2(new_n1229), .ZN(G225));
endmodule


