//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  OAI21_X1  g0004(.A(G50), .B1(G58), .B2(G68), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n210), .B(new_n214), .C1(new_n223), .C2(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G250), .B(G257), .Z(new_n226));
  XNOR2_X1  g0026(.A(G264), .B(G270), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT65), .Z(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n229), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(G1698), .ZN(new_n249));
  AND2_X1   g0049(.A1(new_n249), .A2(G222), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT3), .B(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  INV_X1    g0053(.A(G77), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n251), .ZN(new_n255));
  OR3_X1    g0055(.A1(new_n250), .A2(new_n255), .A3(KEYINPUT68), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT68), .B1(new_n250), .B2(new_n255), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n256), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n264), .A2(new_n258), .A3(G274), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT67), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT67), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n258), .A2(new_n270), .A3(new_n267), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n265), .B1(new_n272), .B2(G226), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n261), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G179), .ZN(new_n275));
  AOI21_X1  g0075(.A(G169), .B1(new_n261), .B2(new_n273), .ZN(new_n276));
  INV_X1    g0076(.A(G50), .ZN(new_n277));
  INV_X1    g0077(.A(G58), .ZN(new_n278));
  INV_X1    g0078(.A(G68), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n280), .A2(G20), .B1(G150), .B2(new_n281), .ZN(new_n282));
  OR2_X1    g0082(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT69), .A2(KEYINPUT8), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n278), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT70), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT8), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT70), .B1(new_n288), .B2(G58), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n287), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n208), .A2(G33), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n282), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n207), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n293), .A2(new_n207), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G1), .B2(new_n208), .ZN(new_n298));
  MUX2_X1   g0098(.A(new_n296), .B(new_n298), .S(G50), .Z(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n275), .A2(new_n276), .A3(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n249), .A2(G232), .B1(G107), .B2(new_n248), .ZN(new_n303));
  INV_X1    g0103(.A(G238), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n252), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n259), .ZN(new_n306));
  INV_X1    g0106(.A(G274), .ZN(new_n307));
  AND2_X1   g0107(.A1(G1), .A2(G13), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n257), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n264), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n272), .A2(G244), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n306), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT72), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT8), .B(G58), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(new_n281), .B1(G20), .B2(G77), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT15), .B(G87), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n291), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n296), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n266), .A2(KEYINPUT71), .A3(G13), .A4(G20), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n318), .A2(new_n294), .B1(new_n254), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n294), .B1(new_n320), .B2(new_n321), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n325), .B(G77), .C1(G1), .C2(new_n208), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n312), .A2(G190), .B1(new_n313), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n324), .A2(new_n326), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n306), .A2(new_n310), .A3(new_n311), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n329), .A2(KEYINPUT72), .B1(new_n330), .B2(G200), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n312), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n327), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n300), .B(KEYINPUT9), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n274), .A2(G200), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n261), .A2(G190), .A3(new_n273), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT10), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT10), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n339), .A2(new_n344), .A3(new_n340), .A4(new_n341), .ZN(new_n345));
  AOI211_X1 g0145(.A(new_n302), .B(new_n338), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(G58), .B(G68), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G20), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n281), .A2(G159), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n248), .A2(new_n208), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT75), .B1(new_n246), .B2(G33), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT75), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(new_n244), .A3(KEYINPUT3), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n356), .A3(new_n247), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n353), .A2(G20), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n352), .A2(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n351), .B1(new_n359), .B2(new_n279), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n297), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT7), .B1(new_n248), .B2(new_n208), .ZN(new_n363));
  AOI211_X1 g0163(.A(new_n353), .B(G20), .C1(new_n245), .C2(new_n247), .ZN(new_n364));
  OAI21_X1  g0164(.A(G68), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(KEYINPUT16), .A3(new_n351), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(KEYINPUT74), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT74), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n353), .B1(new_n251), .B2(G20), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n248), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n350), .B1(new_n371), .B2(G68), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n368), .B1(new_n372), .B2(KEYINPUT16), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n362), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n290), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n298), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n290), .A2(new_n296), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G1698), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n253), .A2(new_n380), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n380), .A2(G226), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n251), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G87), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n258), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n310), .B1(new_n231), .B2(new_n268), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n387), .A2(new_n335), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(G179), .B2(new_n387), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n379), .A2(KEYINPUT18), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT76), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n389), .B1(new_n374), .B2(new_n378), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(KEYINPUT76), .A3(KEYINPUT18), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT18), .ZN(new_n396));
  INV_X1    g0196(.A(new_n378), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n366), .A2(KEYINPUT74), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n372), .A2(new_n368), .A3(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n400), .B2(new_n362), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n396), .B1(new_n401), .B2(new_n389), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n393), .A2(new_n395), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G190), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n387), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(G200), .B2(new_n387), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n374), .A2(new_n378), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT17), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(KEYINPUT77), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n279), .A2(G20), .ZN(new_n410));
  INV_X1    g0210(.A(new_n281), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n410), .B1(new_n291), .B2(new_n254), .C1(new_n411), .C2(new_n277), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n294), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT11), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n325), .B(G68), .C1(G1), .C2(new_n208), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G13), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(G1), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n419), .A2(new_n410), .A3(KEYINPUT12), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n323), .A2(new_n279), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(KEYINPUT12), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT73), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  NOR2_X1   g0225(.A1(G226), .A2(G1698), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n231), .B2(G1698), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n427), .A2(new_n251), .B1(G33), .B2(G97), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n310), .B1(new_n428), .B2(new_n258), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n304), .B1(new_n269), .B2(new_n271), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT13), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n231), .A2(G1698), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G226), .B2(G1698), .ZN(new_n434));
  INV_X1    g0234(.A(G97), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n434), .A2(new_n248), .B1(new_n244), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n265), .B1(new_n436), .B2(new_n259), .ZN(new_n437));
  INV_X1    g0237(.A(new_n271), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n270), .B1(new_n258), .B2(new_n267), .ZN(new_n439));
  OAI21_X1  g0239(.A(G238), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n432), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n425), .B(G169), .C1(new_n431), .C2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT13), .B1(new_n429), .B2(new_n430), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n437), .A2(new_n440), .A3(new_n432), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(G179), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n444), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n425), .B1(new_n447), .B2(G169), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n424), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(G169), .B1(new_n431), .B2(new_n441), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT14), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(KEYINPUT73), .A3(new_n445), .A4(new_n442), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n423), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n447), .A2(G200), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n443), .A2(G190), .A3(new_n444), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n423), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n346), .A2(new_n409), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n403), .A2(new_n408), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT77), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n208), .C1(G33), .C2(new_n435), .ZN(new_n465));
  INV_X1    g0265(.A(G116), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G20), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n294), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n465), .A2(KEYINPUT20), .A3(new_n294), .A4(new_n467), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n466), .B1(new_n266), .B2(G33), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n470), .A2(new_n471), .B1(new_n325), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT83), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n322), .B2(G116), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n320), .A2(KEYINPUT83), .A3(new_n466), .A4(new_n321), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT84), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n473), .A2(new_n477), .A3(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT78), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(G41), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n262), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n263), .A2(G1), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n488), .A2(new_n258), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G270), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n309), .A2(new_n486), .A3(new_n485), .A4(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n245), .A2(new_n247), .A3(G257), .A4(new_n380), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT81), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT81), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n251), .A2(new_n496), .A3(G257), .A4(new_n380), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n248), .A2(G303), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n251), .A2(G264), .A3(G1698), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT82), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n500), .A2(new_n501), .A3(new_n259), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n500), .B2(new_n259), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n493), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n482), .A2(G169), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT21), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(G200), .ZN(new_n508));
  INV_X1    g0308(.A(new_n481), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT84), .B1(new_n473), .B2(new_n477), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n493), .B(G190), .C1(new_n502), .C2(new_n503), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n500), .A2(new_n259), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n500), .A2(new_n501), .A3(new_n259), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n492), .A2(new_n333), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n482), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n482), .A2(KEYINPUT21), .A3(G169), .A4(new_n504), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n507), .A2(new_n513), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G107), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n357), .A2(new_n358), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(new_n369), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n522), .A2(KEYINPUT6), .A3(G97), .ZN(new_n525));
  XNOR2_X1  g0325(.A(G97), .B(G107), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n528), .A2(new_n208), .B1(new_n254), .B2(new_n411), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n294), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n418), .A2(G20), .A3(new_n435), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n266), .A2(G33), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n297), .A2(new_n296), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n533), .B2(new_n435), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n488), .A2(G257), .A3(new_n258), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n491), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n245), .A2(new_n247), .A3(G244), .A4(new_n380), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n251), .A2(KEYINPUT4), .A3(G244), .A4(new_n380), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n251), .A2(G250), .A3(G1698), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n464), .A4(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n537), .B1(new_n543), .B2(new_n259), .ZN(new_n544));
  INV_X1    g0344(.A(G200), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n530), .B(new_n535), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(G190), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT79), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n544), .A2(KEYINPUT79), .A3(G190), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n544), .A2(new_n333), .ZN(new_n552));
  AND2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n527), .B1(new_n553), .B2(new_n202), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n522), .A2(KEYINPUT6), .A3(G97), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(G20), .B1(G77), .B2(new_n281), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n359), .B2(new_n522), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n534), .B1(new_n558), .B2(new_n294), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n543), .A2(new_n259), .ZN(new_n560));
  INV_X1    g0360(.A(new_n537), .ZN(new_n561));
  AOI21_X1  g0361(.A(G169), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n552), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(G87), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n533), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n245), .A2(new_n247), .A3(new_n208), .A4(G68), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n291), .B2(new_n435), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n208), .A2(new_n570), .B1(new_n202), .B2(new_n564), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n294), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n323), .A2(new_n317), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n565), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n245), .A2(new_n247), .A3(G244), .A4(G1698), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n245), .A2(new_n247), .A3(G238), .A4(new_n380), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G116), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n259), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n258), .A2(G274), .A3(new_n487), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n266), .A2(G45), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n258), .A2(G250), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G200), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n259), .B2(new_n579), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G190), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n575), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n586), .A2(new_n335), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n317), .B(KEYINPUT80), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n572), .B(new_n573), .C1(new_n533), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n333), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n551), .A2(new_n563), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n488), .A2(G264), .A3(new_n258), .ZN(new_n598));
  MUX2_X1   g0398(.A(G250), .B(G257), .S(G1698), .Z(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(new_n251), .B1(G33), .B2(G294), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n491), .B(new_n598), .C1(new_n600), .C2(new_n258), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G169), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT87), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n598), .A2(KEYINPUT88), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT88), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n488), .A2(new_n606), .A3(G264), .A4(new_n258), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n599), .A2(new_n251), .ZN(new_n609));
  NAND2_X1  g0409(.A1(G33), .A2(G294), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n258), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n608), .A2(new_n612), .A3(G179), .A4(new_n491), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n601), .A2(KEYINPUT87), .A3(G169), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n604), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n245), .A2(new_n247), .A3(new_n208), .A4(G87), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT22), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT22), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n251), .A2(new_n618), .A3(new_n208), .A4(G87), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n578), .A2(G20), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n522), .A2(KEYINPUT23), .A3(G20), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT23), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n208), .B2(G107), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n621), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g0426(.A(KEYINPUT85), .B(KEYINPUT24), .Z(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n620), .A2(new_n625), .A3(new_n627), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n294), .A3(new_n630), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n419), .A2(new_n208), .A3(G107), .ZN(new_n632));
  NAND2_X1  g0432(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n633));
  OR2_X1    g0433(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  OAI221_X1 g0435(.A(new_n635), .B1(new_n633), .B2(new_n632), .C1(new_n533), .C2(new_n522), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n615), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n611), .B1(new_n605), .B2(new_n607), .ZN(new_n640));
  AOI21_X1  g0440(.A(G200), .B1(new_n640), .B2(new_n491), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n601), .A2(G190), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n631), .B(new_n637), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT89), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n639), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n639), .B2(new_n643), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n597), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n463), .A2(new_n521), .A3(new_n647), .ZN(G372));
  NAND2_X1  g0448(.A1(new_n343), .A2(new_n345), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n407), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n449), .A2(new_n452), .ZN(new_n652));
  INV_X1    g0452(.A(new_n423), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n337), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n456), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n402), .A2(new_n391), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n649), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n302), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT90), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n574), .B(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n587), .A2(new_n589), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n595), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n640), .A2(new_n491), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n642), .B1(new_n667), .B2(new_n545), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(new_n638), .ZN(new_n669));
  NOR4_X1   g0469(.A1(new_n666), .A2(new_n669), .A3(new_n551), .A4(new_n563), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n507), .A2(new_n519), .A3(new_n520), .ZN(new_n671));
  INV_X1    g0471(.A(new_n639), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n596), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n563), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT26), .ZN(new_n676));
  INV_X1    g0476(.A(new_n595), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n664), .B2(new_n663), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT26), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(new_n563), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n676), .A2(new_n680), .A3(new_n595), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n673), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n661), .B1(new_n463), .B2(new_n684), .ZN(G369));
  OR3_X1    g0485(.A1(new_n419), .A2(KEYINPUT27), .A3(G20), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT27), .B1(new_n419), .B2(G20), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G213), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G343), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n511), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n671), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n521), .B2(new_n692), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  INV_X1    g0495(.A(new_n646), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n639), .A2(new_n643), .A3(new_n644), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n638), .A2(new_n690), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n639), .B2(new_n691), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n695), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n671), .A2(new_n691), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n698), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n672), .A2(new_n691), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n212), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n205), .B2(new_n712), .ZN(new_n715));
  XOR2_X1   g0515(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n716));
  XNOR2_X1  g0516(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT93), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n608), .A2(new_n612), .A3(new_n588), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n517), .A2(new_n518), .A3(new_n544), .A4(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n721), .B(new_n537), .C1(new_n259), .C2(new_n543), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n517), .A2(new_n723), .A3(new_n518), .A4(new_n719), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n544), .A2(G179), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n580), .A2(KEYINPUT92), .A3(new_n585), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT92), .B1(new_n580), .B2(new_n585), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n504), .A2(new_n667), .A3(new_n725), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n722), .A2(new_n724), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT31), .B1(new_n730), .B2(new_n690), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n718), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AND4_X1   g0533(.A1(new_n507), .A2(new_n513), .A3(new_n519), .A4(new_n520), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n698), .A2(new_n734), .A3(new_n597), .A4(new_n691), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n720), .A2(new_n721), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n729), .A2(new_n724), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n690), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(KEYINPUT93), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n733), .A2(new_n735), .A3(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n595), .B1(new_n675), .B2(KEYINPUT26), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n679), .B1(new_n678), .B2(new_n563), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n690), .B1(new_n673), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT29), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(KEYINPUT29), .B(new_n690), .C1(new_n673), .C2(new_n682), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n744), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n717), .B1(new_n752), .B2(G1), .ZN(G364));
  NOR2_X1   g0553(.A1(new_n417), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n266), .B1(new_n754), .B2(G45), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n711), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n695), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G330), .B2(new_n694), .ZN(new_n759));
  INV_X1    g0559(.A(new_n757), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n208), .A2(G179), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n761), .A2(new_n404), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(G283), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G329), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n762), .A2(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT97), .Z(new_n768));
  NOR3_X1   g0568(.A1(new_n404), .A2(G179), .A3(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n208), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n208), .A2(new_n333), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n404), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G294), .A2(new_n771), .B1(new_n774), .B2(G326), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n772), .A2(new_n764), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n248), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n772), .A2(G190), .A3(new_n545), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n778), .B1(G322), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n773), .A2(G190), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT33), .B(G317), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n761), .A2(G190), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n782), .A2(new_n783), .B1(new_n785), .B2(G303), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n775), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n251), .B1(new_n776), .B2(new_n254), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G58), .B2(new_n780), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n771), .A2(G97), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n785), .A2(G87), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT32), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n765), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n762), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n792), .A2(new_n794), .B1(new_n795), .B2(G107), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n789), .A2(new_n790), .A3(new_n791), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n782), .A2(G68), .ZN(new_n798));
  INV_X1    g0598(.A(new_n774), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n798), .B1(new_n792), .B2(new_n794), .C1(new_n799), .C2(new_n277), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n768), .A2(new_n787), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n207), .B1(G20), .B2(new_n335), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n760), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n239), .A2(G45), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n710), .A2(new_n251), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n804), .B(new_n805), .C1(G45), .C2(new_n205), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n251), .A2(new_n212), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT94), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n808), .A2(G355), .B1(new_n466), .B2(new_n710), .ZN(new_n809));
  AOI21_X1  g0609(.A(KEYINPUT95), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n806), .A2(KEYINPUT95), .A3(new_n809), .ZN(new_n811));
  NOR2_X1   g0611(.A1(G13), .A2(G33), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(G20), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT96), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n802), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n803), .B1(new_n810), .B2(new_n818), .C1(new_n694), .C2(new_n815), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n759), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  AOI21_X1  g0621(.A(new_n690), .B1(new_n673), .B2(new_n682), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n337), .A2(new_n690), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n327), .A2(new_n690), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n332), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n823), .B1(new_n825), .B2(new_n337), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n822), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n743), .A2(G330), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n757), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  INV_X1    g0630(.A(new_n776), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n780), .A2(G143), .B1(new_n831), .B2(G159), .ZN(new_n832));
  INV_X1    g0632(.A(G137), .ZN(new_n833));
  INV_X1    g0633(.A(G150), .ZN(new_n834));
  INV_X1    g0634(.A(new_n782), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n832), .B1(new_n799), .B2(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n795), .A2(G68), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n840), .B(new_n251), .C1(new_n841), .C2(new_n765), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n770), .A2(new_n278), .B1(new_n784), .B2(new_n277), .ZN(new_n843));
  NOR4_X1   g0643(.A1(new_n838), .A2(new_n839), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n774), .A2(G303), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n835), .B2(new_n763), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n776), .A2(new_n466), .B1(new_n765), .B2(new_n777), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n251), .B(new_n847), .C1(G294), .C2(new_n780), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n762), .A2(new_n564), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n848), .A2(new_n790), .A3(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n846), .B(new_n851), .C1(G107), .C2(new_n785), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n802), .B1(new_n844), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n802), .A2(new_n812), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n760), .B1(new_n254), .B2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(new_n826), .C2(new_n813), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n830), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(G384));
  OR2_X1    g0658(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n859), .A2(new_n860), .A3(G116), .A4(new_n209), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT36), .Z(new_n862));
  OAI211_X1 g0662(.A(new_n206), .B(G77), .C1(new_n278), .C2(new_n279), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n277), .A2(G68), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n266), .B(G13), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n823), .B1(new_n822), .B2(new_n826), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n449), .A2(new_n452), .A3(new_n456), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT98), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n423), .A2(new_n691), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n871), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n654), .A2(new_n456), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n870), .B1(new_n869), .B2(new_n871), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT99), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n877), .B(new_n294), .C1(new_n372), .C2(KEYINPUT16), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT16), .B1(new_n365), .B2(new_n351), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT99), .B1(new_n879), .B2(new_n297), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n400), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n389), .B1(new_n881), .B2(new_n378), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n374), .A2(new_n378), .A3(new_n406), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT100), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT100), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n294), .B1(new_n372), .B2(KEYINPUT16), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n399), .A2(new_n398), .B1(new_n886), .B2(KEYINPUT99), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n397), .B1(new_n887), .B2(new_n878), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n885), .B(new_n407), .C1(new_n888), .C2(new_n389), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n881), .A2(new_n378), .ZN(new_n890));
  INV_X1    g0690(.A(new_n688), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n884), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT37), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n883), .A2(new_n394), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n379), .A2(new_n891), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n892), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n460), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n379), .A2(new_n390), .ZN(new_n903));
  AND4_X1   g0703(.A1(new_n896), .A2(new_n903), .A3(new_n897), .A4(new_n407), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n893), .B2(KEYINPUT37), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n892), .B1(new_n403), .B2(new_n408), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n868), .B(new_n876), .C1(new_n902), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n658), .A2(new_n688), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n654), .A2(new_n690), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT39), .B1(new_n902), .B2(new_n908), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT101), .B1(new_n915), .B2(new_n904), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n903), .A2(new_n407), .ZN(new_n917));
  INV_X1    g0717(.A(new_n897), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT37), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT101), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n898), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n918), .B1(new_n658), .B2(new_n651), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n916), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n907), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n925));
  XOR2_X1   g0725(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n913), .B1(new_n914), .B2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n911), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n459), .B(new_n462), .C1(new_n750), .C2(new_n751), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n661), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT103), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n929), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n825), .A2(new_n337), .ZN(new_n934));
  INV_X1    g0734(.A(new_n823), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n731), .A2(new_n732), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n937), .B2(new_n735), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n938), .A2(new_n876), .A3(KEYINPUT104), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT104), .B1(new_n938), .B2(new_n876), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT40), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n924), .B2(new_n925), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n647), .A2(new_n521), .A3(new_n690), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n740), .A2(new_n741), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n826), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n869), .A2(new_n871), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT98), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n453), .A2(new_n457), .A3(new_n871), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n902), .B2(new_n908), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n941), .A2(new_n943), .B1(new_n953), .B2(new_n942), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n463), .B1(new_n735), .B2(new_n937), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(G330), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n955), .B2(new_n957), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n933), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n933), .A2(new_n959), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT105), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n960), .B1(new_n266), .B2(new_n754), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n961), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(KEYINPUT105), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n866), .B1(new_n963), .B2(new_n965), .ZN(G367));
  NOR2_X1   g0766(.A1(new_n551), .A2(new_n563), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n559), .B2(new_n691), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n563), .A2(new_n690), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n705), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT42), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n968), .A2(new_n639), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n691), .B1(new_n974), .B2(new_n563), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n663), .A2(new_n691), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT106), .B1(new_n978), .B2(new_n678), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n978), .A2(KEYINPUT106), .A3(new_n678), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n979), .B(new_n980), .C1(new_n677), .C2(new_n977), .ZN(new_n981));
  XNOR2_X1  g0781(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT43), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n976), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT108), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT108), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n976), .A2(new_n988), .A3(new_n983), .A4(new_n985), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n987), .B(new_n989), .C1(new_n976), .C2(new_n983), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n702), .A2(new_n971), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n990), .B(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n711), .B(KEYINPUT41), .Z(new_n995));
  INV_X1    g0795(.A(KEYINPUT44), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT109), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n707), .A2(new_n997), .A3(new_n971), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n997), .B1(new_n707), .B2(new_n971), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n996), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1000), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1002), .A2(KEYINPUT44), .A3(new_n998), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n708), .A2(KEYINPUT45), .A3(new_n970), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT45), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n707), .B2(new_n971), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1001), .A2(new_n1003), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n702), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT110), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT110), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1008), .A2(new_n1012), .A3(new_n1009), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n705), .B1(new_n701), .B2(new_n704), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(new_n695), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n752), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1001), .A2(new_n1003), .A3(new_n702), .A4(new_n1007), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1011), .A2(new_n1013), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n995), .B1(new_n1019), .B2(new_n752), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n994), .B1(new_n1020), .B2(new_n756), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n817), .B1(new_n212), .B2(new_n317), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n228), .A2(new_n710), .A3(new_n251), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n757), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n762), .A2(new_n254), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n770), .A2(new_n279), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(G58), .C2(new_n785), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n248), .B1(new_n780), .B2(G150), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n765), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G50), .A2(new_n831), .B1(new_n1029), .B2(G137), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G143), .A2(new_n774), .B1(new_n782), .B2(G159), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n780), .A2(G303), .B1(new_n831), .B2(G283), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT46), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n784), .B2(new_n466), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n785), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(KEYINPUT111), .B(G317), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n251), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n762), .A2(new_n435), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G294), .B2(new_n782), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n522), .B2(new_n770), .C1(new_n777), .C2(new_n799), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1032), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT47), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1024), .B1(new_n1044), .B2(new_n802), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT112), .Z(new_n1046));
  NAND2_X1  g0846(.A1(new_n981), .A2(new_n816), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1021), .A2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT113), .Z(G387));
  OR2_X1    g0851(.A1(new_n234), .A2(new_n263), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n713), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n1052), .A2(new_n805), .B1(new_n1053), .B2(new_n808), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n713), .B(new_n263), .C1(new_n279), .C2(new_n254), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT50), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n315), .B2(new_n277), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n314), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n1054), .A2(new_n1059), .B1(G107), .B2(new_n212), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n817), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n757), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n701), .A2(new_n815), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n779), .A2(new_n277), .B1(new_n776), .B2(new_n279), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n248), .B(new_n1064), .C1(G150), .C2(new_n1029), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n375), .A2(new_n782), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n784), .A2(new_n254), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1040), .B(new_n1067), .C1(G159), .C2(new_n774), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n592), .A2(new_n770), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n251), .B1(new_n1029), .B2(G326), .ZN(new_n1071));
  INV_X1    g0871(.A(G294), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n770), .A2(new_n763), .B1(new_n784), .B2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n780), .A2(new_n1037), .B1(new_n831), .B2(G303), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n774), .A2(G322), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n777), .C2(new_n835), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT49), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1071), .B1(new_n466), .B2(new_n762), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1070), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1062), .B(new_n1063), .C1(new_n802), .C2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1015), .B2(new_n756), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1016), .A2(new_n711), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1015), .A2(new_n752), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(G393));
  AND2_X1   g0888(.A1(new_n1010), .A2(new_n1018), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1019), .B(new_n711), .C1(new_n1017), .C2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n971), .A2(new_n816), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n817), .B1(new_n435), .B2(new_n212), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n242), .A2(new_n805), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n757), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n782), .A2(G50), .B1(new_n831), .B2(new_n315), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1095), .A2(KEYINPUT114), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(KEYINPUT114), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n248), .B(new_n849), .C1(G143), .C2(new_n1029), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n771), .A2(G77), .B1(new_n785), .B2(G68), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G150), .A2(new_n774), .B1(new_n780), .B2(G159), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT51), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G317), .A2(new_n774), .B1(new_n780), .B2(G311), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT52), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n771), .A2(G116), .B1(new_n785), .B2(G283), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n782), .A2(G303), .B1(new_n795), .B2(G107), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n831), .A2(G294), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n251), .B1(new_n1029), .B2(G322), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1100), .A2(new_n1102), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1094), .B1(new_n1110), .B2(new_n802), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1089), .A2(new_n756), .B1(new_n1091), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1090), .A2(new_n1112), .ZN(G390));
  NAND3_X1  g0913(.A1(new_n914), .A2(new_n812), .A3(new_n927), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n802), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n791), .A2(new_n248), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT117), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n776), .A2(new_n435), .B1(new_n765), .B2(new_n1072), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G116), .B2(new_n780), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G107), .A2(new_n782), .B1(new_n774), .B2(G283), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n771), .A2(G77), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n840), .A4(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n774), .A2(G128), .B1(new_n795), .B2(G50), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n833), .B2(new_n835), .C1(new_n793), .C2(new_n770), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n780), .A2(G132), .B1(new_n1029), .B2(G125), .ZN(new_n1125));
  OR3_X1    g0925(.A1(new_n784), .A2(KEYINPUT53), .A3(new_n834), .ZN(new_n1126));
  OAI21_X1  g0926(.A(KEYINPUT53), .B1(new_n784), .B2(new_n834), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n248), .B1(new_n831), .B2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1117), .A2(new_n1122), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT118), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1115), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1133), .B2(new_n1132), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n760), .B1(new_n290), .B2(new_n854), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1114), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n913), .B1(new_n867), .B2(new_n951), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n914), .A2(new_n1138), .A3(new_n927), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n924), .A2(new_n925), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n823), .B1(new_n748), .B2(new_n934), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n913), .C1(new_n951), .C2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n938), .A2(new_n876), .A3(G330), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT115), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n744), .A2(new_n1147), .A3(new_n826), .A4(new_n876), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n743), .A2(new_n876), .A3(G330), .A4(new_n826), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(KEYINPUT115), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1151), .A2(new_n1139), .A3(new_n1142), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n937), .A2(new_n735), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n459), .A2(G330), .A3(new_n462), .A4(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n930), .A2(new_n1155), .A3(new_n661), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(G330), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n951), .B1(new_n946), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n1141), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n951), .B1(new_n828), .B2(new_n936), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n867), .B1(new_n1162), .B2(new_n1144), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1157), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT116), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1151), .A2(new_n1139), .A3(new_n1142), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1144), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1164), .B(new_n1165), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1160), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1150), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1149), .A2(KEYINPUT115), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1162), .A2(new_n1144), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n868), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1156), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(new_n1146), .A3(new_n1152), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1168), .A2(new_n711), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1165), .B1(new_n1153), .B2(new_n1164), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1137), .B1(new_n755), .B2(new_n1153), .C1(new_n1177), .C2(new_n1178), .ZN(G378));
  NAND2_X1  g0979(.A1(new_n649), .A2(new_n660), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n301), .A2(new_n688), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n649), .B(new_n660), .C1(new_n301), .C2(new_n688), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1184), .B(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n954), .B2(G330), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n953), .A2(new_n942), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT104), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n946), .B2(new_n951), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n938), .A2(new_n876), .A3(KEYINPUT104), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1140), .A2(KEYINPUT40), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  AND4_X1   g0993(.A1(G330), .A2(new_n1189), .A3(new_n1193), .A4(new_n1187), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n929), .B1(new_n1188), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1189), .A2(new_n1193), .A3(G330), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1187), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n954), .A2(G330), .A3(new_n1187), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n911), .A2(new_n928), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1195), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1176), .A2(new_n1157), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(KEYINPUT57), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n711), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G128), .A2(new_n780), .B1(new_n785), .B2(new_n1129), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT121), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G150), .A2(new_n771), .B1(new_n782), .B2(G132), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n774), .A2(G125), .B1(new_n831), .B2(G137), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT122), .Z(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n795), .A2(G159), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G33), .B(G41), .C1(new_n1029), .C2(G124), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n251), .A2(G41), .ZN(new_n1220));
  AOI211_X1 g1020(.A(G50), .B(new_n1220), .C1(new_n244), .C2(new_n262), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT119), .Z(new_n1222));
  NOR2_X1   g1022(.A1(new_n762), .A2(new_n278), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n835), .A2(new_n435), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(G116), .C2(new_n774), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1220), .B1(new_n763), .B2(new_n765), .C1(new_n522), .C2(new_n779), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1226), .A2(new_n1026), .A3(new_n1067), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1225), .B(new_n1227), .C1(new_n592), .C2(new_n776), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT58), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1222), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT120), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n1230), .A2(new_n1231), .B1(new_n1229), .B2(new_n1228), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1231), .B2(new_n1230), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1115), .B1(new_n1219), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n854), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n757), .B1(G50), .B2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1234), .B(new_n1236), .C1(new_n1197), .C2(new_n812), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1202), .B2(new_n756), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1207), .A2(new_n1238), .ZN(G375));
  AOI22_X1  g1039(.A1(G150), .A2(new_n831), .B1(new_n1029), .B2(G128), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1240), .B(new_n251), .C1(new_n833), .C2(new_n779), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1223), .B(new_n1241), .C1(new_n782), .C2(new_n1129), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n770), .A2(new_n277), .B1(new_n784), .B2(new_n793), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G132), .B2(new_n774), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n466), .A2(new_n835), .B1(new_n799), .B2(new_n1072), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1025), .B(new_n1245), .C1(G97), .C2(new_n785), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n251), .B1(new_n1029), .B2(G303), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n780), .A2(G283), .B1(new_n831), .B2(G107), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1069), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1242), .A2(new_n1244), .B1(new_n1246), .B2(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n757), .B1(G68), .B2(new_n1235), .C1(new_n1250), .C2(new_n1115), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n951), .B2(new_n812), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1252), .B1(new_n1254), .B2(new_n756), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1157), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n995), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1164), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1255), .B1(new_n1256), .B2(new_n1258), .ZN(G381));
  INV_X1    g1059(.A(G387), .ZN(new_n1260));
  INV_X1    g1060(.A(G375), .ZN(new_n1261));
  OR2_X1    g1061(.A1(G393), .A2(G396), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1262), .A2(G384), .ZN(new_n1263));
  NOR4_X1   g1063(.A1(G378), .A2(G390), .A3(new_n1263), .A4(G381), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1260), .A2(new_n1261), .A3(new_n1264), .ZN(G407));
  OAI21_X1  g1065(.A(new_n1137), .B1(new_n1153), .B2(new_n755), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1168), .A2(new_n711), .A3(new_n1176), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1178), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1261), .A2(new_n689), .A3(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(G407), .A2(G213), .A3(new_n1270), .ZN(G409));
  NAND2_X1  g1071(.A1(G393), .A2(G396), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT113), .B1(new_n1262), .B2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(G390), .A2(new_n1273), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1090), .A2(new_n1112), .B1(new_n1262), .B2(new_n1272), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1021), .B(new_n1049), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1262), .A2(new_n1272), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1090), .B(new_n1112), .C1(new_n1277), .C2(KEYINPUT113), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1262), .A2(new_n1272), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G390), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1020), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n993), .B1(new_n1281), .B2(new_n755), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1278), .B(new_n1280), .C1(new_n1282), .C2(new_n1048), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1276), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G378), .B(new_n1238), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1202), .A2(new_n1257), .A3(new_n1203), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1238), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT123), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1288), .A2(new_n1289), .A3(new_n1269), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1289), .B1(new_n1288), .B2(new_n1269), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1286), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT124), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1164), .A2(KEYINPUT60), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n712), .B1(new_n1295), .B2(new_n1256), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1256), .B2(new_n1295), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1255), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n857), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1297), .A2(G384), .A3(new_n1255), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(KEYINPUT124), .B(new_n1286), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n689), .A2(G213), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1294), .A2(new_n1301), .A3(new_n1302), .A4(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT62), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1292), .A2(new_n1303), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1301), .A2(KEYINPUT62), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1304), .A2(new_n1305), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT61), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n689), .A2(G213), .A3(G2897), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1301), .B(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1309), .B1(new_n1311), .B2(new_n1306), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1285), .B1(new_n1308), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1304), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1294), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1310), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1301), .B(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1292), .A2(new_n1303), .A3(new_n1321), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1276), .A2(new_n1283), .A3(new_n1309), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  AND4_X1   g1125(.A1(new_n1314), .A2(new_n1316), .A3(new_n1320), .A4(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1324), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1314), .B1(new_n1327), .B2(new_n1316), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1313), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(KEYINPUT126), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT126), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1331), .B(new_n1313), .C1(new_n1326), .C2(new_n1328), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1332), .ZN(G405));
  NOR2_X1   g1133(.A1(new_n1261), .A2(G378), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1286), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1301), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  NOR3_X1   g1137(.A1(new_n1334), .A2(new_n1301), .A3(new_n1335), .ZN(new_n1338));
  OAI22_X1  g1138(.A1(new_n1337), .A2(new_n1338), .B1(KEYINPUT127), .B2(new_n1284), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1284), .A2(KEYINPUT127), .ZN(new_n1340));
  XOR2_X1   g1140(.A(new_n1339), .B(new_n1340), .Z(G402));
endmodule


