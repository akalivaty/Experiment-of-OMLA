

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U547 ( .A1(n542), .A2(G651), .ZN(n792) );
  NOR2_X1 U548 ( .A1(n542), .A2(n540), .ZN(n798) );
  AND2_X1 U549 ( .A1(G2105), .A2(G2104), .ZN(n894) );
  NOR2_X1 U550 ( .A1(n649), .A2(n915), .ZN(n600) );
  NOR2_X2 U551 ( .A1(G164), .A2(G1384), .ZN(n704) );
  XNOR2_X2 U552 ( .A(n536), .B(KEYINPUT88), .ZN(G164) );
  INV_X1 U553 ( .A(KEYINPUT104), .ZN(n687) );
  AND2_X1 U554 ( .A1(n933), .A2(n515), .ZN(n690) );
  XNOR2_X1 U555 ( .A(n523), .B(KEYINPUT17), .ZN(n705) );
  INV_X1 U556 ( .A(n598), .ZN(n668) );
  NAND2_X1 U557 ( .A1(n683), .A2(n516), .ZN(n685) );
  BUF_X1 U558 ( .A(n706), .Z(n891) );
  AND2_X1 U559 ( .A1(n700), .A2(n514), .ZN(n701) );
  NAND2_X1 U560 ( .A1(n706), .A2(G101), .ZN(n522) );
  AND2_X1 U561 ( .A1(n526), .A2(n525), .ZN(n513) );
  OR2_X1 U562 ( .A1(n699), .A2(n698), .ZN(n514) );
  OR2_X1 U563 ( .A1(n698), .A2(n689), .ZN(n515) );
  NOR2_X1 U564 ( .A1(n682), .A2(n698), .ZN(n516) );
  INV_X1 U565 ( .A(G2105), .ZN(n521) );
  XOR2_X1 U566 ( .A(n664), .B(n663), .Z(n517) );
  AND2_X1 U567 ( .A1(n939), .A2(n749), .ZN(n518) );
  NOR2_X1 U568 ( .A1(n737), .A2(n518), .ZN(n519) );
  XOR2_X1 U569 ( .A(KEYINPUT98), .B(n628), .Z(n520) );
  INV_X1 U570 ( .A(KEYINPUT26), .ZN(n599) );
  INV_X1 U571 ( .A(KEYINPUT97), .ZN(n621) );
  INV_X1 U572 ( .A(G8), .ZN(n651) );
  NOR2_X1 U573 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U574 ( .A1(G1966), .A2(n698), .ZN(n650) );
  INV_X1 U575 ( .A(KEYINPUT101), .ZN(n663) );
  NOR2_X1 U576 ( .A1(G2084), .A2(n668), .ZN(n652) );
  XNOR2_X1 U577 ( .A(n675), .B(KEYINPUT32), .ZN(n676) );
  INV_X1 U578 ( .A(KEYINPUT94), .ZN(n596) );
  INV_X1 U579 ( .A(KEYINPUT64), .ZN(n684) );
  XNOR2_X1 U580 ( .A(n685), .B(n684), .ZN(n686) );
  INV_X1 U581 ( .A(G2104), .ZN(n524) );
  AND2_X1 U582 ( .A1(n521), .A2(G2104), .ZN(n706) );
  BUF_X1 U583 ( .A(n705), .Z(n890) );
  XOR2_X1 U584 ( .A(KEYINPUT15), .B(n620), .Z(n937) );
  NOR2_X1 U585 ( .A1(n610), .A2(n609), .ZN(n612) );
  XNOR2_X1 U586 ( .A(n522), .B(KEYINPUT23), .ZN(n529) );
  NOR2_X1 U587 ( .A1(n529), .A2(n528), .ZN(G160) );
  NAND2_X1 U588 ( .A1(n521), .A2(n524), .ZN(n523) );
  NAND2_X1 U589 ( .A1(n705), .A2(G137), .ZN(n527) );
  AND2_X1 U590 ( .A1(n524), .A2(G2105), .ZN(n710) );
  NAND2_X1 U591 ( .A1(G125), .A2(n710), .ZN(n526) );
  NAND2_X1 U592 ( .A1(G113), .A2(n894), .ZN(n525) );
  NAND2_X1 U593 ( .A1(n527), .A2(n513), .ZN(n528) );
  NAND2_X1 U594 ( .A1(n705), .A2(G138), .ZN(n535) );
  NAND2_X1 U595 ( .A1(G102), .A2(n706), .ZN(n531) );
  NAND2_X1 U596 ( .A1(G114), .A2(n894), .ZN(n530) );
  AND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n533) );
  NAND2_X1 U598 ( .A1(G126), .A2(n710), .ZN(n532) );
  AND2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  AND2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U601 ( .A1(G543), .A2(G651), .ZN(n801) );
  NAND2_X1 U602 ( .A1(G91), .A2(n801), .ZN(n538) );
  XOR2_X1 U603 ( .A(KEYINPUT0), .B(G543), .Z(n542) );
  INV_X1 U604 ( .A(G651), .ZN(n540) );
  NAND2_X1 U605 ( .A1(G78), .A2(n798), .ZN(n537) );
  NAND2_X1 U606 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U607 ( .A(KEYINPUT66), .B(n539), .Z(n546) );
  NOR2_X1 U608 ( .A1(G543), .A2(n540), .ZN(n541) );
  XOR2_X2 U609 ( .A(KEYINPUT1), .B(n541), .Z(n794) );
  NAND2_X1 U610 ( .A1(G65), .A2(n794), .ZN(n544) );
  NAND2_X1 U611 ( .A1(G53), .A2(n792), .ZN(n543) );
  AND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(G299) );
  NAND2_X1 U614 ( .A1(G52), .A2(n792), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(KEYINPUT65), .ZN(n554) );
  NAND2_X1 U616 ( .A1(G90), .A2(n801), .ZN(n549) );
  NAND2_X1 U617 ( .A1(G77), .A2(n798), .ZN(n548) );
  NAND2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n550), .B(KEYINPUT9), .ZN(n552) );
  NAND2_X1 U620 ( .A1(G64), .A2(n794), .ZN(n551) );
  NAND2_X1 U621 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U622 ( .A1(n554), .A2(n553), .ZN(G171) );
  XNOR2_X1 U623 ( .A(KEYINPUT70), .B(KEYINPUT6), .ZN(n558) );
  NAND2_X1 U624 ( .A1(G63), .A2(n794), .ZN(n556) );
  NAND2_X1 U625 ( .A1(G51), .A2(n792), .ZN(n555) );
  NAND2_X1 U626 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n558), .B(n557), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n801), .A2(G89), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U630 ( .A1(G76), .A2(n798), .ZN(n560) );
  NAND2_X1 U631 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U632 ( .A(KEYINPUT5), .B(n562), .ZN(n563) );
  XNOR2_X1 U633 ( .A(KEYINPUT69), .B(n563), .ZN(n564) );
  NOR2_X1 U634 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U635 ( .A(KEYINPUT7), .B(n566), .Z(G168) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(n801), .A2(G88), .ZN(n567) );
  XNOR2_X1 U638 ( .A(n567), .B(KEYINPUT84), .ZN(n569) );
  NAND2_X1 U639 ( .A1(G75), .A2(n798), .ZN(n568) );
  NAND2_X1 U640 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U641 ( .A1(G62), .A2(n794), .ZN(n571) );
  NAND2_X1 U642 ( .A1(G50), .A2(n792), .ZN(n570) );
  NAND2_X1 U643 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U644 ( .A1(n573), .A2(n572), .ZN(G166) );
  INV_X1 U645 ( .A(G166), .ZN(G303) );
  NAND2_X1 U646 ( .A1(G49), .A2(n792), .ZN(n575) );
  NAND2_X1 U647 ( .A1(G74), .A2(G651), .ZN(n574) );
  NAND2_X1 U648 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U649 ( .A1(n794), .A2(n576), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n542), .A2(G87), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n578), .A2(n577), .ZN(G288) );
  NAND2_X1 U652 ( .A1(G86), .A2(n801), .ZN(n579) );
  XNOR2_X1 U653 ( .A(n579), .B(KEYINPUT82), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G73), .A2(n798), .ZN(n580) );
  XOR2_X1 U655 ( .A(KEYINPUT2), .B(n580), .Z(n581) );
  XNOR2_X1 U656 ( .A(n581), .B(KEYINPUT83), .ZN(n583) );
  NAND2_X1 U657 ( .A1(G48), .A2(n792), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U659 ( .A1(G61), .A2(n794), .ZN(n584) );
  XNOR2_X1 U660 ( .A(KEYINPUT81), .B(n584), .ZN(n585) );
  NOR2_X1 U661 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(G305) );
  NAND2_X1 U663 ( .A1(G85), .A2(n801), .ZN(n590) );
  NAND2_X1 U664 ( .A1(G72), .A2(n798), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G60), .A2(n794), .ZN(n592) );
  NAND2_X1 U667 ( .A1(G47), .A2(n792), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n593) );
  OR2_X1 U669 ( .A1(n594), .A2(n593), .ZN(G290) );
  NAND2_X1 U670 ( .A1(G160), .A2(G40), .ZN(n703) );
  XNOR2_X1 U671 ( .A(n703), .B(n596), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n704), .A2(n597), .ZN(n649) );
  INV_X1 U673 ( .A(n649), .ZN(n598) );
  NAND2_X1 U674 ( .A1(G8), .A2(n652), .ZN(n665) );
  INV_X1 U675 ( .A(G1996), .ZN(n915) );
  XNOR2_X1 U676 ( .A(n600), .B(n599), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n668), .A2(G1341), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n613) );
  XNOR2_X1 U679 ( .A(KEYINPUT67), .B(KEYINPUT13), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n801), .A2(G81), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n603), .B(KEYINPUT12), .ZN(n605) );
  NAND2_X1 U682 ( .A1(G68), .A2(n798), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U684 ( .A(n607), .B(n606), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n794), .A2(G56), .ZN(n608) );
  XOR2_X1 U686 ( .A(KEYINPUT14), .B(n608), .Z(n609) );
  NAND2_X1 U687 ( .A1(n792), .A2(G43), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n936) );
  NOR2_X1 U689 ( .A1(n613), .A2(n936), .ZN(n627) );
  NAND2_X1 U690 ( .A1(G92), .A2(n801), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G79), .A2(n798), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U693 ( .A1(G66), .A2(n794), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G54), .A2(n792), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n627), .A2(n937), .ZN(n622) );
  XNOR2_X1 U698 ( .A(n622), .B(n621), .ZN(n626) );
  INV_X1 U699 ( .A(n668), .ZN(n644) );
  NOR2_X1 U700 ( .A1(n644), .A2(G1348), .ZN(n624) );
  NOR2_X1 U701 ( .A1(G2067), .A2(n668), .ZN(n623) );
  NOR2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n629) );
  NOR2_X1 U704 ( .A1(n627), .A2(n937), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n520), .ZN(n631) );
  INV_X1 U706 ( .A(KEYINPUT99), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n631), .B(n630), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n644), .A2(G2072), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT27), .ZN(n634) );
  INV_X1 U710 ( .A(G1956), .ZN(n967) );
  NOR2_X1 U711 ( .A1(n967), .A2(n644), .ZN(n633) );
  NOR2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n638) );
  INV_X1 U713 ( .A(G299), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n641) );
  NOR2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U717 ( .A(n639), .B(KEYINPUT28), .Z(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n643) );
  XOR2_X1 U719 ( .A(KEYINPUT100), .B(KEYINPUT29), .Z(n642) );
  XNOR2_X1 U720 ( .A(n643), .B(n642), .ZN(n648) );
  OR2_X1 U721 ( .A1(n644), .A2(G1961), .ZN(n646) );
  XNOR2_X1 U722 ( .A(G2078), .B(KEYINPUT25), .ZN(n912) );
  NAND2_X1 U723 ( .A1(n644), .A2(n912), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n646), .A2(n645), .ZN(n656) );
  NAND2_X1 U725 ( .A1(n656), .A2(G171), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n648), .A2(n647), .ZN(n661) );
  NAND2_X1 U727 ( .A1(G8), .A2(n649), .ZN(n698) );
  XOR2_X1 U728 ( .A(KEYINPUT96), .B(n650), .Z(n662) );
  NAND2_X1 U729 ( .A1(n662), .A2(n653), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n654), .B(KEYINPUT30), .ZN(n655) );
  NOR2_X1 U731 ( .A1(G168), .A2(n655), .ZN(n658) );
  NOR2_X1 U732 ( .A1(G171), .A2(n656), .ZN(n657) );
  NOR2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U734 ( .A(KEYINPUT31), .B(n659), .Z(n660) );
  NAND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n666), .A2(n662), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n665), .A2(n517), .ZN(n677) );
  NAND2_X1 U738 ( .A1(G286), .A2(n666), .ZN(n673) );
  NOR2_X1 U739 ( .A1(G1971), .A2(n698), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n667), .B(KEYINPUT102), .ZN(n670) );
  NOR2_X1 U741 ( .A1(n668), .A2(G2090), .ZN(n669) );
  NOR2_X1 U742 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U743 ( .A1(G303), .A2(n671), .ZN(n672) );
  NAND2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U745 ( .A1(n674), .A2(G8), .ZN(n675) );
  NAND2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n679) );
  INV_X1 U747 ( .A(KEYINPUT103), .ZN(n678) );
  XNOR2_X1 U748 ( .A(n679), .B(n678), .ZN(n693) );
  NOR2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n943) );
  NOR2_X1 U750 ( .A1(G1971), .A2(G303), .ZN(n680) );
  NOR2_X1 U751 ( .A1(n943), .A2(n680), .ZN(n681) );
  NAND2_X1 U752 ( .A1(n693), .A2(n681), .ZN(n683) );
  NAND2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n940) );
  INV_X1 U754 ( .A(n940), .ZN(n682) );
  NOR2_X1 U755 ( .A1(n686), .A2(KEYINPUT33), .ZN(n688) );
  XNOR2_X1 U756 ( .A(n688), .B(n687), .ZN(n691) );
  XOR2_X1 U757 ( .A(G1981), .B(G305), .Z(n933) );
  NAND2_X1 U758 ( .A1(n943), .A2(KEYINPUT33), .ZN(n689) );
  NAND2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n702) );
  NOR2_X1 U760 ( .A1(G2090), .A2(G303), .ZN(n692) );
  NAND2_X1 U761 ( .A1(G8), .A2(n692), .ZN(n694) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U763 ( .A1(n695), .A2(n698), .ZN(n700) );
  NOR2_X1 U764 ( .A1(G1981), .A2(G305), .ZN(n696) );
  XNOR2_X1 U765 ( .A(n696), .B(KEYINPUT24), .ZN(n697) );
  XNOR2_X1 U766 ( .A(n697), .B(KEYINPUT95), .ZN(n699) );
  NAND2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n738) );
  NOR2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n749) );
  NAND2_X1 U769 ( .A1(G140), .A2(n890), .ZN(n708) );
  NAND2_X1 U770 ( .A1(G104), .A2(n891), .ZN(n707) );
  NAND2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U772 ( .A(KEYINPUT34), .B(n709), .ZN(n716) );
  NAND2_X1 U773 ( .A1(n710), .A2(G128), .ZN(n711) );
  XOR2_X1 U774 ( .A(KEYINPUT89), .B(n711), .Z(n713) );
  NAND2_X1 U775 ( .A1(n894), .A2(G116), .ZN(n712) );
  NAND2_X1 U776 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U777 ( .A(KEYINPUT35), .B(n714), .Z(n715) );
  NOR2_X1 U778 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U779 ( .A(KEYINPUT36), .B(n717), .Z(n885) );
  XOR2_X1 U780 ( .A(KEYINPUT37), .B(G2067), .Z(n746) );
  AND2_X1 U781 ( .A1(n885), .A2(n746), .ZN(n1009) );
  NAND2_X1 U782 ( .A1(n749), .A2(n1009), .ZN(n744) );
  XOR2_X1 U783 ( .A(KEYINPUT90), .B(G1991), .Z(n911) );
  NAND2_X1 U784 ( .A1(G131), .A2(n890), .ZN(n719) );
  NAND2_X1 U785 ( .A1(G95), .A2(n891), .ZN(n718) );
  NAND2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U787 ( .A1(G119), .A2(n710), .ZN(n721) );
  NAND2_X1 U788 ( .A1(G107), .A2(n894), .ZN(n720) );
  NAND2_X1 U789 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n870) );
  NOR2_X1 U791 ( .A1(n911), .A2(n870), .ZN(n734) );
  XOR2_X1 U792 ( .A(KEYINPUT91), .B(KEYINPUT38), .Z(n725) );
  NAND2_X1 U793 ( .A1(G105), .A2(n891), .ZN(n724) );
  XNOR2_X1 U794 ( .A(n725), .B(n724), .ZN(n732) );
  NAND2_X1 U795 ( .A1(G129), .A2(n710), .ZN(n727) );
  NAND2_X1 U796 ( .A1(G117), .A2(n894), .ZN(n726) );
  NAND2_X1 U797 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U798 ( .A1(n890), .A2(G141), .ZN(n728) );
  XOR2_X1 U799 ( .A(KEYINPUT92), .B(n728), .Z(n729) );
  NOR2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U801 ( .A1(n732), .A2(n731), .ZN(n874) );
  AND2_X1 U802 ( .A1(n874), .A2(G1996), .ZN(n733) );
  NOR2_X1 U803 ( .A1(n734), .A2(n733), .ZN(n1010) );
  XNOR2_X1 U804 ( .A(KEYINPUT93), .B(n749), .ZN(n735) );
  NOR2_X1 U805 ( .A1(n1010), .A2(n735), .ZN(n741) );
  INV_X1 U806 ( .A(n741), .ZN(n736) );
  NAND2_X1 U807 ( .A1(n744), .A2(n736), .ZN(n737) );
  XNOR2_X1 U808 ( .A(G1986), .B(G290), .ZN(n939) );
  NAND2_X1 U809 ( .A1(n738), .A2(n519), .ZN(n752) );
  NOR2_X1 U810 ( .A1(G1996), .A2(n874), .ZN(n998) );
  AND2_X1 U811 ( .A1(n911), .A2(n870), .ZN(n1005) );
  NOR2_X1 U812 ( .A1(G1986), .A2(G290), .ZN(n739) );
  NOR2_X1 U813 ( .A1(n1005), .A2(n739), .ZN(n740) );
  NOR2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U815 ( .A1(n998), .A2(n742), .ZN(n743) );
  XNOR2_X1 U816 ( .A(n743), .B(KEYINPUT39), .ZN(n745) );
  NAND2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n748) );
  NOR2_X1 U818 ( .A1(n885), .A2(n746), .ZN(n747) );
  XNOR2_X1 U819 ( .A(KEYINPUT105), .B(n747), .ZN(n1002) );
  NAND2_X1 U820 ( .A1(n748), .A2(n1002), .ZN(n750) );
  NAND2_X1 U821 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U822 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U823 ( .A(n753), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U824 ( .A(G2443), .B(G2446), .Z(n755) );
  XNOR2_X1 U825 ( .A(G2427), .B(G2451), .ZN(n754) );
  XNOR2_X1 U826 ( .A(n755), .B(n754), .ZN(n761) );
  XOR2_X1 U827 ( .A(G2430), .B(G2454), .Z(n757) );
  XNOR2_X1 U828 ( .A(G1348), .B(G1341), .ZN(n756) );
  XNOR2_X1 U829 ( .A(n757), .B(n756), .ZN(n759) );
  XOR2_X1 U830 ( .A(G2435), .B(G2438), .Z(n758) );
  XNOR2_X1 U831 ( .A(n759), .B(n758), .ZN(n760) );
  XOR2_X1 U832 ( .A(n761), .B(n760), .Z(n762) );
  AND2_X1 U833 ( .A1(G14), .A2(n762), .ZN(G401) );
  AND2_X1 U834 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U835 ( .A(G132), .ZN(G219) );
  INV_X1 U836 ( .A(G82), .ZN(G220) );
  INV_X1 U837 ( .A(G57), .ZN(G237) );
  NAND2_X1 U838 ( .A1(G7), .A2(G661), .ZN(n763) );
  XNOR2_X1 U839 ( .A(n763), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U840 ( .A(G223), .ZN(n828) );
  NAND2_X1 U841 ( .A1(n828), .A2(G567), .ZN(n764) );
  XOR2_X1 U842 ( .A(KEYINPUT11), .B(n764), .Z(G234) );
  INV_X1 U843 ( .A(G860), .ZN(n770) );
  OR2_X1 U844 ( .A1(n936), .A2(n770), .ZN(G153) );
  NAND2_X1 U845 ( .A1(G171), .A2(G868), .ZN(n766) );
  INV_X1 U846 ( .A(G868), .ZN(n811) );
  NAND2_X1 U847 ( .A1(n937), .A2(n811), .ZN(n765) );
  NAND2_X1 U848 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U849 ( .A(KEYINPUT68), .B(n767), .Z(G284) );
  NOR2_X1 U850 ( .A1(G286), .A2(n811), .ZN(n769) );
  NOR2_X1 U851 ( .A1(G868), .A2(G299), .ZN(n768) );
  NOR2_X1 U852 ( .A1(n769), .A2(n768), .ZN(G297) );
  NAND2_X1 U853 ( .A1(n770), .A2(G559), .ZN(n771) );
  NAND2_X1 U854 ( .A1(n771), .A2(n937), .ZN(n772) );
  XNOR2_X1 U855 ( .A(n772), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U856 ( .A1(G868), .A2(n936), .ZN(n775) );
  NAND2_X1 U857 ( .A1(G868), .A2(n937), .ZN(n773) );
  NOR2_X1 U858 ( .A1(G559), .A2(n773), .ZN(n774) );
  NOR2_X1 U859 ( .A1(n775), .A2(n774), .ZN(G282) );
  NAND2_X1 U860 ( .A1(G123), .A2(n710), .ZN(n776) );
  XOR2_X1 U861 ( .A(KEYINPUT18), .B(n776), .Z(n777) );
  XNOR2_X1 U862 ( .A(n777), .B(KEYINPUT71), .ZN(n779) );
  NAND2_X1 U863 ( .A1(G135), .A2(n890), .ZN(n778) );
  NAND2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U865 ( .A(KEYINPUT72), .B(n780), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G99), .A2(n891), .ZN(n781) );
  XNOR2_X1 U867 ( .A(KEYINPUT73), .B(n781), .ZN(n782) );
  NOR2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U869 ( .A1(n894), .A2(G111), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n1006) );
  XNOR2_X1 U871 ( .A(G2096), .B(n1006), .ZN(n786) );
  NOR2_X1 U872 ( .A1(G2100), .A2(n786), .ZN(n787) );
  XOR2_X1 U873 ( .A(KEYINPUT74), .B(n787), .Z(G156) );
  XOR2_X1 U874 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n788) );
  XNOR2_X1 U875 ( .A(G305), .B(n788), .ZN(n791) );
  XNOR2_X1 U876 ( .A(G166), .B(G299), .ZN(n789) );
  XNOR2_X1 U877 ( .A(n789), .B(G288), .ZN(n790) );
  XNOR2_X1 U878 ( .A(n791), .B(n790), .ZN(n807) );
  NAND2_X1 U879 ( .A1(n792), .A2(G55), .ZN(n793) );
  XNOR2_X1 U880 ( .A(n793), .B(KEYINPUT78), .ZN(n796) );
  NAND2_X1 U881 ( .A1(G67), .A2(n794), .ZN(n795) );
  NAND2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U883 ( .A(n797), .B(KEYINPUT79), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G80), .A2(n798), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U886 ( .A1(G93), .A2(n801), .ZN(n802) );
  XNOR2_X1 U887 ( .A(KEYINPUT77), .B(n802), .ZN(n803) );
  NOR2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U889 ( .A(KEYINPUT80), .B(n805), .Z(n835) );
  XNOR2_X1 U890 ( .A(G290), .B(n835), .ZN(n806) );
  XNOR2_X1 U891 ( .A(n807), .B(n806), .ZN(n838) );
  XNOR2_X1 U892 ( .A(n936), .B(KEYINPUT75), .ZN(n809) );
  NAND2_X1 U893 ( .A1(n937), .A2(G559), .ZN(n808) );
  XNOR2_X1 U894 ( .A(n809), .B(n808), .ZN(n832) );
  XOR2_X1 U895 ( .A(n838), .B(n832), .Z(n810) );
  NOR2_X1 U896 ( .A1(n811), .A2(n810), .ZN(n813) );
  NOR2_X1 U897 ( .A1(n835), .A2(G868), .ZN(n812) );
  NOR2_X1 U898 ( .A1(n813), .A2(n812), .ZN(G295) );
  NAND2_X1 U899 ( .A1(G2084), .A2(G2078), .ZN(n814) );
  XOR2_X1 U900 ( .A(KEYINPUT20), .B(n814), .Z(n815) );
  NAND2_X1 U901 ( .A1(G2090), .A2(n815), .ZN(n816) );
  XNOR2_X1 U902 ( .A(KEYINPUT21), .B(n816), .ZN(n817) );
  NAND2_X1 U903 ( .A1(n817), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U904 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U905 ( .A1(G69), .A2(G120), .ZN(n818) );
  NOR2_X1 U906 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U907 ( .A1(G108), .A2(n819), .ZN(n836) );
  NAND2_X1 U908 ( .A1(n836), .A2(G567), .ZN(n825) );
  NOR2_X1 U909 ( .A1(G220), .A2(G219), .ZN(n820) );
  XNOR2_X1 U910 ( .A(KEYINPUT22), .B(n820), .ZN(n821) );
  NAND2_X1 U911 ( .A1(n821), .A2(G96), .ZN(n822) );
  NOR2_X1 U912 ( .A1(G218), .A2(n822), .ZN(n823) );
  XOR2_X1 U913 ( .A(KEYINPUT86), .B(n823), .Z(n837) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n837), .ZN(n824) );
  NAND2_X1 U915 ( .A1(n825), .A2(n824), .ZN(n910) );
  NAND2_X1 U916 ( .A1(G661), .A2(G483), .ZN(n826) );
  XOR2_X1 U917 ( .A(KEYINPUT87), .B(n826), .Z(n827) );
  NOR2_X1 U918 ( .A1(n910), .A2(n827), .ZN(n831) );
  NAND2_X1 U919 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U922 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(G188) );
  XOR2_X1 U925 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  XOR2_X1 U927 ( .A(n832), .B(KEYINPUT76), .Z(n833) );
  NOR2_X1 U928 ( .A1(G860), .A2(n833), .ZN(n834) );
  XOR2_X1 U929 ( .A(n835), .B(n834), .Z(G145) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G69), .ZN(G235) );
  NOR2_X1 U932 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XOR2_X1 U934 ( .A(KEYINPUT112), .B(n838), .Z(n840) );
  XNOR2_X1 U935 ( .A(n937), .B(G286), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n936), .B(G171), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n843) );
  NOR2_X1 U939 ( .A1(G37), .A2(n843), .ZN(G397) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2078), .Z(n845) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2084), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U943 ( .A(n846), .B(G2100), .Z(n848) );
  XNOR2_X1 U944 ( .A(G2090), .B(G2072), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n850) );
  XNOR2_X1 U947 ( .A(KEYINPUT107), .B(G2678), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n852), .B(n851), .Z(G227) );
  XNOR2_X1 U950 ( .A(G1961), .B(KEYINPUT108), .ZN(n862) );
  XOR2_X1 U951 ( .A(G1976), .B(G1971), .Z(n854) );
  XNOR2_X1 U952 ( .A(G1986), .B(G1956), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U954 ( .A(G1981), .B(G1966), .Z(n856) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U957 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U958 ( .A(G2474), .B(KEYINPUT41), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U961 ( .A1(n710), .A2(G124), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G100), .A2(n891), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U965 ( .A1(G136), .A2(n890), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G112), .A2(n894), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U969 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n872) );
  XNOR2_X1 U970 ( .A(n870), .B(KEYINPUT46), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(n873), .B(G162), .Z(n876) );
  XOR2_X1 U973 ( .A(G160), .B(n874), .Z(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n888) );
  NAND2_X1 U975 ( .A1(G130), .A2(n710), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G118), .A2(n894), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n884) );
  NAND2_X1 U978 ( .A1(n890), .A2(G142), .ZN(n879) );
  XOR2_X1 U979 ( .A(KEYINPUT109), .B(n879), .Z(n881) );
  NAND2_X1 U980 ( .A1(n891), .A2(G106), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U982 ( .A(n882), .B(KEYINPUT45), .Z(n883) );
  NOR2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n886) );
  XOR2_X1 U984 ( .A(n886), .B(n885), .Z(n887) );
  XOR2_X1 U985 ( .A(n888), .B(n887), .Z(n889) );
  XNOR2_X1 U986 ( .A(G164), .B(n889), .ZN(n902) );
  NAND2_X1 U987 ( .A1(G139), .A2(n890), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G103), .A2(n891), .ZN(n892) );
  NAND2_X1 U989 ( .A1(n893), .A2(n892), .ZN(n899) );
  NAND2_X1 U990 ( .A1(G127), .A2(n710), .ZN(n896) );
  NAND2_X1 U991 ( .A1(G115), .A2(n894), .ZN(n895) );
  NAND2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n897), .Z(n898) );
  NOR2_X1 U994 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U995 ( .A(KEYINPUT110), .B(n900), .Z(n993) );
  XNOR2_X1 U996 ( .A(n1006), .B(n993), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U998 ( .A1(G37), .A2(n903), .ZN(G395) );
  NOR2_X1 U999 ( .A1(G401), .A2(n910), .ZN(n907) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n904), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G397), .A2(n905), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n907), .A2(n906), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(n908), .A2(G395), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n909), .B(KEYINPUT113), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(n910), .ZN(G319) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  INV_X1 U1009 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U1010 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1022) );
  XOR2_X1 U1011 ( .A(G2090), .B(G35), .Z(n927) );
  XOR2_X1 U1012 ( .A(n911), .B(G25), .Z(n914) );
  XOR2_X1 U1013 ( .A(n912), .B(G27), .Z(n913) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n923) );
  XNOR2_X1 U1015 ( .A(G32), .B(n915), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n916), .A2(G28), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(G2067), .B(G26), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(G2072), .B(G33), .ZN(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(n919), .B(KEYINPUT115), .ZN(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(n924), .B(KEYINPUT116), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n925), .B(KEYINPUT53), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(G34), .B(G2084), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(KEYINPUT54), .B(n928), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1029 ( .A(KEYINPUT55), .B(n931), .Z(n932) );
  NOR2_X1 U1030 ( .A1(G29), .A2(n932), .ZN(n990) );
  XNOR2_X1 U1031 ( .A(G16), .B(KEYINPUT56), .ZN(n958) );
  XNOR2_X1 U1032 ( .A(G1966), .B(G168), .ZN(n934) );
  NAND2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(KEYINPUT57), .B(n935), .ZN(n956) );
  XOR2_X1 U1035 ( .A(n936), .B(G1341), .Z(n953) );
  XOR2_X1 U1036 ( .A(G1348), .B(n937), .Z(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(G301), .B(G1961), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G299), .B(G1956), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n950) );
  XOR2_X1 U1044 ( .A(G1971), .B(G303), .Z(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT117), .B(n948), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(KEYINPUT118), .B(n951), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(KEYINPUT119), .B(n954), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n988) );
  INV_X1 U1052 ( .A(G16), .ZN(n986) );
  XNOR2_X1 U1053 ( .A(G1986), .B(G24), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(G1976), .B(KEYINPUT122), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(n959), .B(G23), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(G22), .B(G1971), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(KEYINPUT123), .B(n962), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT58), .B(n965), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n966), .B(KEYINPUT124), .ZN(n980) );
  XNOR2_X1 U1062 ( .A(G20), .B(n967), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G1341), .B(G19), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(G6), .B(G1981), .ZN(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(KEYINPUT120), .B(n972), .ZN(n975) );
  XOR2_X1 U1068 ( .A(KEYINPUT59), .B(G1348), .Z(n973) );
  XNOR2_X1 U1069 ( .A(G4), .B(n973), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1071 ( .A(KEYINPUT60), .B(n976), .Z(n978) );
  XNOR2_X1 U1072 ( .A(G1961), .B(G5), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n983) );
  XOR2_X1 U1075 ( .A(KEYINPUT121), .B(G1966), .Z(n981) );
  XNOR2_X1 U1076 ( .A(G21), .B(n981), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(KEYINPUT61), .B(n984), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(G11), .A2(n991), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(n992), .B(KEYINPUT125), .ZN(n1020) );
  XOR2_X1 U1084 ( .A(G164), .B(G2078), .Z(n995) );
  XNOR2_X1 U1085 ( .A(G2072), .B(n993), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1087 ( .A(KEYINPUT50), .B(n996), .Z(n1001) );
  XOR2_X1 U1088 ( .A(G2090), .B(G162), .Z(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(KEYINPUT51), .B(n999), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1014) );
  XOR2_X1 U1093 ( .A(G160), .B(G2084), .Z(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(KEYINPUT114), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(KEYINPUT52), .B(n1015), .ZN(n1017) );
  INV_X1 U1101 ( .A(KEYINPUT55), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(G29), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(n1022), .B(n1021), .ZN(G150) );
  INV_X1 U1106 ( .A(G150), .ZN(G311) );
endmodule

