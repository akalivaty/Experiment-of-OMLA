

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U553 ( .A1(n523), .A2(G2104), .ZN(n870) );
  INV_X1 U554 ( .A(KEYINPUT28), .ZN(n637) );
  OR2_X1 U555 ( .A1(n923), .A2(n662), .ZN(n669) );
  NOR2_X1 U556 ( .A1(G164), .A2(G1384), .ZN(n621) );
  NOR2_X1 U557 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U558 ( .A1(n551), .A2(n541), .ZN(n777) );
  XNOR2_X1 U559 ( .A(KEYINPUT30), .B(KEYINPUT98), .ZN(n684) );
  XNOR2_X1 U560 ( .A(n685), .B(n684), .ZN(n686) );
  INV_X1 U561 ( .A(n914), .ZN(n713) );
  NOR2_X1 U562 ( .A1(n724), .A2(n713), .ZN(n714) );
  AND2_X1 U563 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U564 ( .A1(n621), .A2(n620), .ZN(n695) );
  NAND2_X1 U565 ( .A1(G8), .A2(n695), .ZN(n724) );
  NOR2_X1 U566 ( .A1(G651), .A2(n551), .ZN(n781) );
  XOR2_X1 U567 ( .A(KEYINPUT1), .B(n542), .Z(n782) );
  NOR2_X1 U568 ( .A1(n535), .A2(n534), .ZN(G160) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XOR2_X2 U570 ( .A(KEYINPUT17), .B(n520), .Z(n869) );
  NAND2_X1 U571 ( .A1(G138), .A2(n869), .ZN(n522) );
  INV_X1 U572 ( .A(G2105), .ZN(n523) );
  NAND2_X1 U573 ( .A1(G102), .A2(n870), .ZN(n521) );
  NAND2_X1 U574 ( .A1(n522), .A2(n521), .ZN(n527) );
  NOR2_X1 U575 ( .A1(G2104), .A2(n523), .ZN(n873) );
  NAND2_X1 U576 ( .A1(G126), .A2(n873), .ZN(n525) );
  AND2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n874) );
  NAND2_X1 U578 ( .A1(G114), .A2(n874), .ZN(n524) );
  NAND2_X1 U579 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U580 ( .A1(n527), .A2(n526), .ZN(G164) );
  NAND2_X1 U581 ( .A1(n873), .A2(G125), .ZN(n531) );
  INV_X1 U582 ( .A(KEYINPUT23), .ZN(n529) );
  NAND2_X1 U583 ( .A1(G101), .A2(n870), .ZN(n528) );
  XNOR2_X1 U584 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U586 ( .A1(G137), .A2(n869), .ZN(n533) );
  NAND2_X1 U587 ( .A1(G113), .A2(n874), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U589 ( .A(G543), .B(KEYINPUT0), .Z(n551) );
  INV_X1 U590 ( .A(G651), .ZN(n541) );
  NAND2_X1 U591 ( .A1(G73), .A2(n777), .ZN(n536) );
  XOR2_X1 U592 ( .A(KEYINPUT77), .B(n536), .Z(n537) );
  XNOR2_X1 U593 ( .A(n537), .B(KEYINPUT2), .ZN(n540) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n538) );
  XNOR2_X1 U595 ( .A(n538), .B(KEYINPUT64), .ZN(n778) );
  NAND2_X1 U596 ( .A1(G86), .A2(n778), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n546) );
  NAND2_X1 U598 ( .A1(G48), .A2(n781), .ZN(n544) );
  NOR2_X1 U599 ( .A1(G543), .A2(n541), .ZN(n542) );
  NAND2_X1 U600 ( .A1(G61), .A2(n782), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U603 ( .A(KEYINPUT78), .B(n547), .Z(G305) );
  NAND2_X1 U604 ( .A1(G49), .A2(n781), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G74), .A2(G651), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U607 ( .A1(n782), .A2(n550), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n551), .A2(G87), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n553), .A2(n552), .ZN(G288) );
  NAND2_X1 U610 ( .A1(G52), .A2(n781), .ZN(n555) );
  NAND2_X1 U611 ( .A1(G64), .A2(n782), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U613 ( .A1(n777), .A2(G77), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G90), .A2(n778), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U617 ( .A1(n560), .A2(n559), .ZN(G171) );
  NAND2_X1 U618 ( .A1(n781), .A2(G51), .ZN(n561) );
  XNOR2_X1 U619 ( .A(n561), .B(KEYINPUT72), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G63), .A2(n782), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U622 ( .A(KEYINPUT6), .B(n564), .ZN(n572) );
  NAND2_X1 U623 ( .A1(n778), .A2(G89), .ZN(n565) );
  XNOR2_X1 U624 ( .A(n565), .B(KEYINPUT4), .ZN(n566) );
  XNOR2_X1 U625 ( .A(n566), .B(KEYINPUT70), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G76), .A2(n777), .ZN(n567) );
  NAND2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U628 ( .A(KEYINPUT71), .B(n569), .ZN(n570) );
  XNOR2_X1 U629 ( .A(KEYINPUT5), .B(n570), .ZN(n571) );
  NOR2_X1 U630 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U631 ( .A(KEYINPUT7), .B(n573), .Z(G168) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U633 ( .A1(n777), .A2(G75), .ZN(n575) );
  NAND2_X1 U634 ( .A1(G88), .A2(n778), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G50), .A2(n781), .ZN(n577) );
  NAND2_X1 U637 ( .A1(G62), .A2(n782), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U639 ( .A1(n579), .A2(n578), .ZN(G166) );
  INV_X1 U640 ( .A(G166), .ZN(G303) );
  NAND2_X1 U641 ( .A1(n777), .A2(G72), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G85), .A2(n778), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U644 ( .A1(G47), .A2(n781), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G60), .A2(n782), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n584) );
  OR2_X1 U647 ( .A1(n585), .A2(n584), .ZN(G290) );
  NAND2_X1 U648 ( .A1(G105), .A2(n870), .ZN(n586) );
  XNOR2_X1 U649 ( .A(n586), .B(KEYINPUT38), .ZN(n593) );
  NAND2_X1 U650 ( .A1(G141), .A2(n869), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G117), .A2(n874), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U653 ( .A1(n873), .A2(G129), .ZN(n589) );
  XOR2_X1 U654 ( .A(KEYINPUT90), .B(n589), .Z(n590) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U656 ( .A1(n593), .A2(n592), .ZN(n866) );
  NAND2_X1 U657 ( .A1(G1996), .A2(n866), .ZN(n602) );
  NAND2_X1 U658 ( .A1(G131), .A2(n869), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G95), .A2(n870), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U661 ( .A1(G119), .A2(n873), .ZN(n596) );
  XNOR2_X1 U662 ( .A(KEYINPUT89), .B(n596), .ZN(n597) );
  NOR2_X1 U663 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U664 ( .A1(n874), .A2(G107), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n600), .A2(n599), .ZN(n867) );
  NAND2_X1 U666 ( .A1(G1991), .A2(n867), .ZN(n601) );
  NAND2_X1 U667 ( .A1(n602), .A2(n601), .ZN(n998) );
  NAND2_X1 U668 ( .A1(G160), .A2(G40), .ZN(n619) );
  NOR2_X1 U669 ( .A1(n621), .A2(n619), .ZN(n743) );
  NAND2_X1 U670 ( .A1(n998), .A2(n743), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n603), .B(KEYINPUT91), .ZN(n737) );
  XOR2_X1 U672 ( .A(KEYINPUT92), .B(n737), .Z(n618) );
  XNOR2_X1 U673 ( .A(KEYINPUT37), .B(G2067), .ZN(n734) );
  XNOR2_X1 U674 ( .A(KEYINPUT35), .B(KEYINPUT87), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n874), .A2(G116), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n604), .B(KEYINPUT86), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G128), .A2(n873), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n608), .B(n607), .ZN(n615) );
  NAND2_X1 U680 ( .A1(n870), .A2(G104), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n609), .B(KEYINPUT84), .ZN(n611) );
  NAND2_X1 U682 ( .A1(G140), .A2(n869), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U684 ( .A(KEYINPUT85), .B(n612), .Z(n613) );
  XNOR2_X1 U685 ( .A(KEYINPUT34), .B(n613), .ZN(n614) );
  NOR2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U687 ( .A(KEYINPUT36), .B(n616), .ZN(n888) );
  NOR2_X1 U688 ( .A1(n734), .A2(n888), .ZN(n1002) );
  NAND2_X1 U689 ( .A1(n1002), .A2(n743), .ZN(n617) );
  XNOR2_X1 U690 ( .A(n617), .B(KEYINPUT88), .ZN(n740) );
  NAND2_X1 U691 ( .A1(n618), .A2(n740), .ZN(n731) );
  INV_X1 U692 ( .A(n619), .ZN(n620) );
  NOR2_X1 U693 ( .A1(G1981), .A2(G305), .ZN(n622) );
  XOR2_X1 U694 ( .A(n622), .B(KEYINPUT24), .Z(n623) );
  NOR2_X1 U695 ( .A1(n724), .A2(n623), .ZN(n729) );
  NOR2_X1 U696 ( .A1(G1976), .A2(G288), .ZN(n712) );
  NAND2_X1 U697 ( .A1(n712), .A2(KEYINPUT33), .ZN(n624) );
  XOR2_X1 U698 ( .A(KEYINPUT101), .B(n624), .Z(n625) );
  NOR2_X1 U699 ( .A1(n724), .A2(n625), .ZN(n718) );
  NAND2_X1 U700 ( .A1(G53), .A2(n781), .ZN(n627) );
  NAND2_X1 U701 ( .A1(G65), .A2(n782), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n777), .A2(G78), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G91), .A2(n778), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n911) );
  INV_X1 U707 ( .A(G2072), .ZN(n990) );
  NOR2_X1 U708 ( .A1(n695), .A2(n990), .ZN(n633) );
  XOR2_X1 U709 ( .A(KEYINPUT95), .B(KEYINPUT27), .Z(n632) );
  XNOR2_X1 U710 ( .A(n633), .B(n632), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n695), .A2(G1956), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U713 ( .A(KEYINPUT96), .B(n636), .Z(n670) );
  NOR2_X1 U714 ( .A1(n911), .A2(n670), .ZN(n638) );
  XNOR2_X1 U715 ( .A(n638), .B(n637), .ZN(n674) );
  NAND2_X1 U716 ( .A1(n782), .A2(G66), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G92), .A2(n778), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U719 ( .A(KEYINPUT68), .B(n641), .ZN(n644) );
  NAND2_X1 U720 ( .A1(G54), .A2(n781), .ZN(n642) );
  XNOR2_X1 U721 ( .A(KEYINPUT69), .B(n642), .ZN(n643) );
  NOR2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n777), .A2(G79), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U725 ( .A(KEYINPUT15), .B(n647), .ZN(n923) );
  NAND2_X1 U726 ( .A1(G81), .A2(n778), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(KEYINPUT12), .ZN(n650) );
  NAND2_X1 U728 ( .A1(G68), .A2(n777), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n651), .B(KEYINPUT13), .ZN(n653) );
  NAND2_X1 U731 ( .A1(G43), .A2(n781), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n782), .A2(G56), .ZN(n654) );
  XOR2_X1 U734 ( .A(KEYINPUT14), .B(n654), .Z(n655) );
  XOR2_X2 U735 ( .A(KEYINPUT66), .B(n657), .Z(n912) );
  INV_X1 U736 ( .A(G1996), .ZN(n942) );
  NOR2_X1 U737 ( .A1(n695), .A2(n942), .ZN(n658) );
  XOR2_X1 U738 ( .A(n658), .B(KEYINPUT26), .Z(n660) );
  NAND2_X1 U739 ( .A1(n695), .A2(G1341), .ZN(n659) );
  NAND2_X1 U740 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U741 ( .A1(n912), .A2(n661), .ZN(n662) );
  NAND2_X1 U742 ( .A1(n923), .A2(n662), .ZN(n667) );
  INV_X1 U743 ( .A(n695), .ZN(n676) );
  INV_X1 U744 ( .A(G1348), .ZN(n971) );
  NOR2_X1 U745 ( .A1(n676), .A2(n971), .ZN(n663) );
  XNOR2_X1 U746 ( .A(n663), .B(KEYINPUT97), .ZN(n665) );
  NAND2_X1 U747 ( .A1(n676), .A2(G2067), .ZN(n664) );
  NAND2_X1 U748 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U749 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U750 ( .A1(n669), .A2(n668), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n911), .A2(n670), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U753 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U754 ( .A(KEYINPUT29), .B(n675), .Z(n681) );
  XNOR2_X1 U755 ( .A(G1961), .B(KEYINPUT93), .ZN(n968) );
  NAND2_X1 U756 ( .A1(n695), .A2(n968), .ZN(n678) );
  XNOR2_X1 U757 ( .A(G2078), .B(KEYINPUT25), .ZN(n948) );
  NAND2_X1 U758 ( .A1(n676), .A2(n948), .ZN(n677) );
  NAND2_X1 U759 ( .A1(n678), .A2(n677), .ZN(n688) );
  NAND2_X1 U760 ( .A1(G171), .A2(n688), .ZN(n679) );
  XNOR2_X1 U761 ( .A(KEYINPUT94), .B(n679), .ZN(n680) );
  NAND2_X1 U762 ( .A1(n681), .A2(n680), .ZN(n694) );
  NOR2_X1 U763 ( .A1(G1966), .A2(n724), .ZN(n706) );
  NOR2_X1 U764 ( .A1(G2084), .A2(n695), .ZN(n703) );
  INV_X1 U765 ( .A(n703), .ZN(n682) );
  NAND2_X1 U766 ( .A1(G8), .A2(n682), .ZN(n683) );
  OR2_X1 U767 ( .A1(n706), .A2(n683), .ZN(n685) );
  NOR2_X1 U768 ( .A1(G168), .A2(n686), .ZN(n687) );
  XNOR2_X1 U769 ( .A(n687), .B(KEYINPUT99), .ZN(n691) );
  NOR2_X1 U770 ( .A1(G171), .A2(n688), .ZN(n689) );
  XOR2_X1 U771 ( .A(KEYINPUT100), .B(n689), .Z(n690) );
  NAND2_X1 U772 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U773 ( .A(n692), .B(KEYINPUT31), .ZN(n693) );
  NAND2_X1 U774 ( .A1(n694), .A2(n693), .ZN(n704) );
  NAND2_X1 U775 ( .A1(n704), .A2(G286), .ZN(n700) );
  NOR2_X1 U776 ( .A1(G1971), .A2(n724), .ZN(n697) );
  NOR2_X1 U777 ( .A1(G2090), .A2(n695), .ZN(n696) );
  NOR2_X1 U778 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U779 ( .A1(n698), .A2(G303), .ZN(n699) );
  NAND2_X1 U780 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U781 ( .A1(n701), .A2(G8), .ZN(n702) );
  XNOR2_X1 U782 ( .A(n702), .B(KEYINPUT32), .ZN(n710) );
  NAND2_X1 U783 ( .A1(G8), .A2(n703), .ZN(n708) );
  INV_X1 U784 ( .A(n704), .ZN(n705) );
  NOR2_X1 U785 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U786 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U787 ( .A1(n710), .A2(n709), .ZN(n721) );
  NOR2_X1 U788 ( .A1(G1971), .A2(G303), .ZN(n711) );
  NOR2_X1 U789 ( .A1(n712), .A2(n711), .ZN(n918) );
  NAND2_X1 U790 ( .A1(n721), .A2(n918), .ZN(n715) );
  NAND2_X1 U791 ( .A1(G1976), .A2(G288), .ZN(n914) );
  NOR2_X1 U792 ( .A1(KEYINPUT33), .A2(n716), .ZN(n717) );
  NOR2_X1 U793 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U794 ( .A(n719), .B(KEYINPUT102), .ZN(n720) );
  XOR2_X1 U795 ( .A(G1981), .B(G305), .Z(n927) );
  NAND2_X1 U796 ( .A1(n720), .A2(n927), .ZN(n727) );
  NOR2_X1 U797 ( .A1(G2090), .A2(G303), .ZN(n722) );
  NAND2_X1 U798 ( .A1(G8), .A2(n722), .ZN(n723) );
  NAND2_X1 U799 ( .A1(n721), .A2(n723), .ZN(n725) );
  NAND2_X1 U800 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U801 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U802 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U803 ( .A1(n731), .A2(n730), .ZN(n733) );
  XNOR2_X1 U804 ( .A(G1986), .B(G290), .ZN(n920) );
  NAND2_X1 U805 ( .A1(n920), .A2(n743), .ZN(n732) );
  NAND2_X1 U806 ( .A1(n733), .A2(n732), .ZN(n746) );
  NAND2_X1 U807 ( .A1(n734), .A2(n888), .ZN(n1009) );
  NOR2_X1 U808 ( .A1(G1996), .A2(n866), .ZN(n1006) );
  NOR2_X1 U809 ( .A1(G1986), .A2(G290), .ZN(n735) );
  NOR2_X1 U810 ( .A1(G1991), .A2(n867), .ZN(n996) );
  NOR2_X1 U811 ( .A1(n735), .A2(n996), .ZN(n736) );
  NOR2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U813 ( .A1(n1006), .A2(n738), .ZN(n739) );
  XNOR2_X1 U814 ( .A(KEYINPUT39), .B(n739), .ZN(n741) );
  NAND2_X1 U815 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U816 ( .A1(n1009), .A2(n742), .ZN(n744) );
  NAND2_X1 U817 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U818 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U819 ( .A(n747), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U820 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U821 ( .A(G57), .ZN(G237) );
  INV_X1 U822 ( .A(G132), .ZN(G219) );
  INV_X1 U823 ( .A(G82), .ZN(G220) );
  XOR2_X1 U824 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n749) );
  NAND2_X1 U825 ( .A1(G7), .A2(G661), .ZN(n748) );
  XNOR2_X1 U826 ( .A(n749), .B(n748), .ZN(G223) );
  INV_X1 U827 ( .A(G223), .ZN(n818) );
  NAND2_X1 U828 ( .A1(n818), .A2(G567), .ZN(n750) );
  XOR2_X1 U829 ( .A(KEYINPUT11), .B(n750), .Z(G234) );
  XOR2_X1 U830 ( .A(G860), .B(KEYINPUT67), .Z(n758) );
  INV_X1 U831 ( .A(n912), .ZN(n751) );
  NAND2_X1 U832 ( .A1(n758), .A2(n751), .ZN(G153) );
  INV_X1 U833 ( .A(G171), .ZN(G301) );
  NAND2_X1 U834 ( .A1(G868), .A2(G301), .ZN(n753) );
  INV_X1 U835 ( .A(n923), .ZN(n762) );
  INV_X1 U836 ( .A(G868), .ZN(n800) );
  NAND2_X1 U837 ( .A1(n762), .A2(n800), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n753), .A2(n752), .ZN(G284) );
  NAND2_X1 U839 ( .A1(n911), .A2(n800), .ZN(n754) );
  XNOR2_X1 U840 ( .A(n754), .B(KEYINPUT73), .ZN(n756) );
  NOR2_X1 U841 ( .A1(n800), .A2(G286), .ZN(n755) );
  NOR2_X1 U842 ( .A1(n756), .A2(n755), .ZN(G297) );
  INV_X1 U843 ( .A(G559), .ZN(n757) );
  NOR2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U845 ( .A1(n762), .A2(n759), .ZN(n760) );
  XOR2_X1 U846 ( .A(KEYINPUT16), .B(n760), .Z(G148) );
  NOR2_X1 U847 ( .A1(n912), .A2(G868), .ZN(n761) );
  XNOR2_X1 U848 ( .A(KEYINPUT74), .B(n761), .ZN(n767) );
  NOR2_X1 U849 ( .A1(n762), .A2(n800), .ZN(n763) );
  XNOR2_X1 U850 ( .A(n763), .B(KEYINPUT75), .ZN(n764) );
  NOR2_X1 U851 ( .A1(G559), .A2(n764), .ZN(n765) );
  XNOR2_X1 U852 ( .A(KEYINPUT76), .B(n765), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(G282) );
  NAND2_X1 U854 ( .A1(G123), .A2(n873), .ZN(n768) );
  XNOR2_X1 U855 ( .A(n768), .B(KEYINPUT18), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n870), .A2(G99), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G135), .A2(n869), .ZN(n772) );
  NAND2_X1 U859 ( .A1(G111), .A2(n874), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n995) );
  XNOR2_X1 U862 ( .A(n995), .B(G2096), .ZN(n776) );
  INV_X1 U863 ( .A(G2100), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(G156) );
  NAND2_X1 U865 ( .A1(n777), .A2(G80), .ZN(n780) );
  NAND2_X1 U866 ( .A1(G93), .A2(n778), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n786) );
  NAND2_X1 U868 ( .A1(G55), .A2(n781), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G67), .A2(n782), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n785) );
  OR2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n799) );
  NAND2_X1 U872 ( .A1(n923), .A2(G559), .ZN(n796) );
  XNOR2_X1 U873 ( .A(n912), .B(n796), .ZN(n787) );
  NOR2_X1 U874 ( .A1(G860), .A2(n787), .ZN(n788) );
  XOR2_X1 U875 ( .A(n799), .B(n788), .Z(G145) );
  XNOR2_X1 U876 ( .A(n912), .B(G305), .ZN(n795) );
  XOR2_X1 U877 ( .A(KEYINPUT79), .B(KEYINPUT19), .Z(n790) );
  XNOR2_X1 U878 ( .A(n911), .B(G166), .ZN(n789) );
  XNOR2_X1 U879 ( .A(n790), .B(n789), .ZN(n791) );
  XNOR2_X1 U880 ( .A(n791), .B(G288), .ZN(n792) );
  XOR2_X1 U881 ( .A(n799), .B(n792), .Z(n793) );
  XNOR2_X1 U882 ( .A(n793), .B(G290), .ZN(n794) );
  XNOR2_X1 U883 ( .A(n795), .B(n794), .ZN(n891) );
  XNOR2_X1 U884 ( .A(n891), .B(n796), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n797), .A2(G868), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n798), .B(KEYINPUT80), .ZN(n802) );
  NAND2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U888 ( .A1(n802), .A2(n801), .ZN(G295) );
  NAND2_X1 U889 ( .A1(G2084), .A2(G2078), .ZN(n805) );
  XNOR2_X1 U890 ( .A(KEYINPUT81), .B(KEYINPUT20), .ZN(n803) );
  XNOR2_X1 U891 ( .A(n803), .B(KEYINPUT82), .ZN(n804) );
  XNOR2_X1 U892 ( .A(n805), .B(n804), .ZN(n806) );
  NAND2_X1 U893 ( .A1(n806), .A2(G2090), .ZN(n807) );
  XNOR2_X1 U894 ( .A(KEYINPUT21), .B(n807), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n808), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U896 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U897 ( .A1(G220), .A2(G219), .ZN(n809) );
  XNOR2_X1 U898 ( .A(KEYINPUT22), .B(n809), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n810), .A2(G96), .ZN(n811) );
  NOR2_X1 U900 ( .A1(n811), .A2(G218), .ZN(n812) );
  XNOR2_X1 U901 ( .A(n812), .B(KEYINPUT83), .ZN(n825) );
  NAND2_X1 U902 ( .A1(n825), .A2(G2106), .ZN(n816) );
  NAND2_X1 U903 ( .A1(G69), .A2(G120), .ZN(n813) );
  NOR2_X1 U904 ( .A1(G237), .A2(n813), .ZN(n814) );
  NAND2_X1 U905 ( .A1(G108), .A2(n814), .ZN(n826) );
  NAND2_X1 U906 ( .A1(n826), .A2(G567), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n827) );
  NAND2_X1 U908 ( .A1(G483), .A2(G661), .ZN(n817) );
  NOR2_X1 U909 ( .A1(n827), .A2(n817), .ZN(n822) );
  NAND2_X1 U910 ( .A1(n822), .A2(G36), .ZN(G176) );
  NAND2_X1 U911 ( .A1(n818), .A2(G2106), .ZN(n819) );
  XNOR2_X1 U912 ( .A(n819), .B(KEYINPUT104), .ZN(G217) );
  NAND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n820) );
  XNOR2_X1 U914 ( .A(KEYINPUT105), .B(n820), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n821), .A2(G661), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G1), .A2(G3), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U918 ( .A(n824), .B(KEYINPUT106), .ZN(G188) );
  INV_X1 U920 ( .A(G120), .ZN(G236) );
  INV_X1 U921 ( .A(G96), .ZN(G221) );
  INV_X1 U922 ( .A(G69), .ZN(G235) );
  NOR2_X1 U923 ( .A1(n826), .A2(n825), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  INV_X1 U925 ( .A(n827), .ZN(G319) );
  XOR2_X1 U926 ( .A(KEYINPUT109), .B(G1986), .Z(n829) );
  XNOR2_X1 U927 ( .A(G1996), .B(G1991), .ZN(n828) );
  XNOR2_X1 U928 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U929 ( .A(n830), .B(KEYINPUT41), .Z(n832) );
  XNOR2_X1 U930 ( .A(G1966), .B(G1981), .ZN(n831) );
  XNOR2_X1 U931 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U932 ( .A(G1976), .B(G1971), .Z(n834) );
  XNOR2_X1 U933 ( .A(G1956), .B(G1961), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U935 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U936 ( .A(KEYINPUT108), .B(G2474), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(G229) );
  XOR2_X1 U938 ( .A(G2678), .B(G2084), .Z(n840) );
  XNOR2_X1 U939 ( .A(G2072), .B(G2078), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U941 ( .A(n841), .B(G2100), .Z(n843) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2090), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U944 ( .A(G2096), .B(KEYINPUT107), .Z(n845) );
  XNOR2_X1 U945 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U947 ( .A(n847), .B(n846), .Z(G227) );
  NAND2_X1 U948 ( .A1(G124), .A2(n873), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U950 ( .A1(n870), .A2(G100), .ZN(n849) );
  NAND2_X1 U951 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U952 ( .A1(G136), .A2(n869), .ZN(n852) );
  NAND2_X1 U953 ( .A1(G112), .A2(n874), .ZN(n851) );
  NAND2_X1 U954 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U955 ( .A1(n854), .A2(n853), .ZN(G162) );
  XNOR2_X1 U956 ( .A(KEYINPUT111), .B(KEYINPUT45), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G142), .A2(n869), .ZN(n856) );
  NAND2_X1 U958 ( .A1(G106), .A2(n870), .ZN(n855) );
  NAND2_X1 U959 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n863) );
  NAND2_X1 U961 ( .A1(n874), .A2(G118), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n859), .B(KEYINPUT110), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G130), .A2(n873), .ZN(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n887) );
  XOR2_X1 U966 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n865) );
  XNOR2_X1 U967 ( .A(G164), .B(KEYINPUT113), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n865), .B(n864), .ZN(n885) );
  XNOR2_X1 U969 ( .A(n995), .B(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(n881) );
  NAND2_X1 U971 ( .A1(G139), .A2(n869), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G103), .A2(n870), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n880) );
  NAND2_X1 U974 ( .A1(G127), .A2(n873), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G115), .A2(n874), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  XNOR2_X1 U978 ( .A(KEYINPUT112), .B(n878), .ZN(n879) );
  NOR2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n991) );
  XOR2_X1 U980 ( .A(n881), .B(n991), .Z(n883) );
  XNOR2_X1 U981 ( .A(G160), .B(G162), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n889) );
  XOR2_X1 U985 ( .A(n889), .B(n888), .Z(n890) );
  NOR2_X1 U986 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U987 ( .A(G286), .B(G301), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n893), .B(n923), .ZN(n894) );
  NOR2_X1 U990 ( .A1(G37), .A2(n894), .ZN(G397) );
  XOR2_X1 U991 ( .A(KEYINPUT103), .B(G2446), .Z(n896) );
  XNOR2_X1 U992 ( .A(G2435), .B(G2438), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n896), .B(n895), .ZN(n903) );
  XOR2_X1 U994 ( .A(G2451), .B(G2430), .Z(n898) );
  XNOR2_X1 U995 ( .A(G2454), .B(G2427), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U997 ( .A(n899), .B(G2443), .Z(n901) );
  XNOR2_X1 U998 ( .A(G1348), .B(G1341), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(n904), .A2(G14), .ZN(n910) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n910), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  INV_X1 U1010 ( .A(n910), .ZN(G401) );
  INV_X1 U1011 ( .A(n911), .ZN(G299) );
  XOR2_X1 U1012 ( .A(n912), .B(G1341), .Z(n922) );
  NAND2_X1 U1013 ( .A1(G1971), .A2(G303), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(G1956), .B(G299), .ZN(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n933) );
  XNOR2_X1 U1020 ( .A(G171), .B(G1961), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(G1348), .B(n923), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(KEYINPUT121), .B(n926), .ZN(n931) );
  XNOR2_X1 U1024 ( .A(G1966), .B(G168), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n929), .B(KEYINPUT57), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1029 ( .A(KEYINPUT122), .B(n934), .Z(n936) );
  XNOR2_X1 U1030 ( .A(KEYINPUT56), .B(G16), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n1022) );
  XOR2_X1 U1032 ( .A(G29), .B(KEYINPUT120), .Z(n959) );
  XOR2_X1 U1033 ( .A(G2084), .B(G34), .Z(n937) );
  XNOR2_X1 U1034 ( .A(KEYINPUT54), .B(n937), .ZN(n955) );
  XNOR2_X1 U1035 ( .A(G2090), .B(G35), .ZN(n953) );
  XNOR2_X1 U1036 ( .A(KEYINPUT117), .B(G2067), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(n938), .B(G26), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(G1991), .B(G25), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(G33), .B(G2072), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1041 ( .A1(G28), .A2(n941), .ZN(n945) );
  XOR2_X1 U1042 ( .A(KEYINPUT118), .B(n942), .Z(n943) );
  XNOR2_X1 U1043 ( .A(G32), .B(n943), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n950) );
  XOR2_X1 U1046 ( .A(G27), .B(n948), .Z(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n951), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n956), .B(KEYINPUT119), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(n957), .B(KEYINPUT55), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(G11), .A2(n960), .ZN(n1020) );
  XOR2_X1 U1055 ( .A(G1986), .B(G24), .Z(n964) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G22), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G23), .B(G1976), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n966) );
  XOR2_X1 U1060 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n965) );
  XNOR2_X1 U1061 ( .A(n966), .B(n965), .ZN(n970) );
  XOR2_X1 U1062 ( .A(KEYINPUT123), .B(G5), .Z(n967) );
  XNOR2_X1 U1063 ( .A(n968), .B(n967), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n985) );
  XNOR2_X1 U1065 ( .A(G1966), .B(G21), .ZN(n982) );
  XNOR2_X1 U1066 ( .A(G4), .B(KEYINPUT59), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(n972), .B(n971), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(G19), .B(G1341), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G1956), .B(G20), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(G1981), .B(G6), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(n979), .B(KEYINPUT60), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n980), .B(KEYINPUT124), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(n983), .B(KEYINPUT125), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1079 ( .A(KEYINPUT61), .B(n986), .Z(n987) );
  NOR2_X1 U1080 ( .A1(G16), .A2(n987), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(KEYINPUT127), .B(n988), .ZN(n1018) );
  XNOR2_X1 U1082 ( .A(G164), .B(G2078), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(n989), .B(KEYINPUT115), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n991), .B(n990), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(KEYINPUT50), .B(n994), .ZN(n1004) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n1000) );
  XOR2_X1 U1088 ( .A(G160), .B(G2084), .Z(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1012) );
  XOR2_X1 U1093 ( .A(G2090), .B(G162), .Z(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(KEYINPUT51), .B(n1007), .Z(n1008) );
  XNOR2_X1 U1096 ( .A(n1008), .B(KEYINPUT114), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT52), .B(n1013), .Z(n1014) );
  NOR2_X1 U1100 ( .A1(KEYINPUT55), .A2(n1014), .ZN(n1015) );
  XOR2_X1 U1101 ( .A(KEYINPUT116), .B(n1015), .Z(n1016) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(G29), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

