

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U545 ( .A(KEYINPUT66), .B(G2104), .Z(n561) );
  NOR2_X1 U546 ( .A1(n561), .A2(G2105), .ZN(n563) );
  NOR2_X1 U547 ( .A1(G299), .A2(n725), .ZN(n710) );
  NOR2_X1 U548 ( .A1(n772), .A2(n784), .ZN(n777) );
  NAND2_X1 U549 ( .A1(n563), .A2(G101), .ZN(n515) );
  XNOR2_X1 U550 ( .A(n780), .B(KEYINPUT108), .ZN(n785) );
  NOR2_X1 U551 ( .A1(n569), .A2(n568), .ZN(n687) );
  BUF_X1 U552 ( .A(n563), .Z(n885) );
  INV_X1 U553 ( .A(n692), .ZN(n704) );
  OR2_X1 U554 ( .A1(n784), .A2(n783), .ZN(n510) );
  XNOR2_X1 U555 ( .A(KEYINPUT96), .B(n817), .ZN(n511) );
  AND2_X1 U556 ( .A1(n511), .A2(n818), .ZN(n512) );
  NOR2_X1 U557 ( .A1(n916), .A2(n715), .ZN(n718) );
  NOR2_X1 U558 ( .A1(G171), .A2(n730), .ZN(n696) );
  XNOR2_X1 U559 ( .A(n743), .B(KEYINPUT32), .ZN(n752) );
  NOR2_X1 U560 ( .A1(n687), .A2(G1384), .ZN(n688) );
  OR2_X1 U561 ( .A1(n768), .A2(n767), .ZN(n779) );
  XNOR2_X1 U562 ( .A(n688), .B(KEYINPUT65), .ZN(n786) );
  AND2_X1 U563 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n513) );
  INV_X1 U565 ( .A(n786), .ZN(n788) );
  BUF_X1 U566 ( .A(n559), .Z(n886) );
  NOR2_X1 U567 ( .A1(G651), .A2(n624), .ZN(n656) );
  BUF_X1 U568 ( .A(n689), .Z(G160) );
  XOR2_X1 U569 ( .A(KEYINPUT68), .B(n513), .Z(n514) );
  XNOR2_X1 U570 ( .A(n514), .B(KEYINPUT17), .ZN(n559) );
  NAND2_X1 U571 ( .A1(G137), .A2(n886), .ZN(n517) );
  XOR2_X1 U572 ( .A(KEYINPUT23), .B(n515), .Z(n516) );
  NAND2_X1 U573 ( .A1(n517), .A2(n516), .ZN(n522) );
  NAND2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XNOR2_X2 U575 ( .A(n518), .B(KEYINPUT67), .ZN(n889) );
  NAND2_X1 U576 ( .A1(G113), .A2(n889), .ZN(n520) );
  AND2_X1 U577 ( .A1(G2105), .A2(n561), .ZN(n890) );
  NAND2_X1 U578 ( .A1(G125), .A2(n890), .ZN(n519) );
  NAND2_X1 U579 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U580 ( .A1(n522), .A2(n521), .ZN(n689) );
  INV_X1 U581 ( .A(G651), .ZN(n527) );
  NOR2_X1 U582 ( .A1(G543), .A2(n527), .ZN(n524) );
  XNOR2_X1 U583 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n523) );
  XNOR2_X1 U584 ( .A(n524), .B(n523), .ZN(n644) );
  NAND2_X1 U585 ( .A1(G64), .A2(n644), .ZN(n526) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n624) );
  NAND2_X1 U587 ( .A1(G52), .A2(n656), .ZN(n525) );
  NAND2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n532) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U590 ( .A1(G90), .A2(n649), .ZN(n529) );
  NOR2_X1 U591 ( .A1(n624), .A2(n527), .ZN(n646) );
  NAND2_X1 U592 ( .A1(G77), .A2(n646), .ZN(n528) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U594 ( .A(KEYINPUT9), .B(n530), .Z(n531) );
  NOR2_X1 U595 ( .A1(n532), .A2(n531), .ZN(G171) );
  NAND2_X1 U596 ( .A1(G78), .A2(n646), .ZN(n534) );
  NAND2_X1 U597 ( .A1(G65), .A2(n644), .ZN(n533) );
  NAND2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n537) );
  NAND2_X1 U599 ( .A1(G91), .A2(n649), .ZN(n535) );
  XNOR2_X1 U600 ( .A(KEYINPUT71), .B(n535), .ZN(n536) );
  NOR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n539) );
  NAND2_X1 U602 ( .A1(n656), .A2(G53), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(G299) );
  XOR2_X1 U604 ( .A(G2446), .B(G2430), .Z(n541) );
  XNOR2_X1 U605 ( .A(G2451), .B(KEYINPUT110), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U607 ( .A(n542), .B(G2427), .Z(n544) );
  XNOR2_X1 U608 ( .A(G1348), .B(G1341), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n548) );
  XOR2_X1 U610 ( .A(G2443), .B(G2435), .Z(n546) );
  XNOR2_X1 U611 ( .A(G2438), .B(G2454), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U613 ( .A(n548), .B(n547), .Z(n549) );
  AND2_X1 U614 ( .A1(G14), .A2(n549), .ZN(G401) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  AND2_X1 U616 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U617 ( .A1(n890), .A2(G123), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(KEYINPUT18), .ZN(n552) );
  NAND2_X1 U619 ( .A1(G135), .A2(n886), .ZN(n551) );
  NAND2_X1 U620 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(KEYINPUT77), .B(n553), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G99), .A2(n885), .ZN(n555) );
  NAND2_X1 U623 ( .A1(G111), .A2(n889), .ZN(n554) );
  AND2_X1 U624 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n988) );
  XNOR2_X1 U626 ( .A(G2096), .B(n988), .ZN(n558) );
  OR2_X1 U627 ( .A1(G2100), .A2(n558), .ZN(G156) );
  INV_X1 U628 ( .A(G108), .ZN(G238) );
  INV_X1 U629 ( .A(G120), .ZN(G236) );
  INV_X1 U630 ( .A(G132), .ZN(G219) );
  AND2_X1 U631 ( .A1(G138), .A2(n559), .ZN(n569) );
  AND2_X1 U632 ( .A1(G2105), .A2(G126), .ZN(n560) );
  NAND2_X1 U633 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U634 ( .A(n562), .B(KEYINPUT92), .ZN(n565) );
  NAND2_X1 U635 ( .A1(n563), .A2(G102), .ZN(n564) );
  AND2_X1 U636 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U637 ( .A1(n889), .A2(G114), .ZN(n566) );
  NAND2_X1 U638 ( .A1(n567), .A2(n566), .ZN(n568) );
  BUF_X1 U639 ( .A(n687), .Z(G164) );
  NAND2_X1 U640 ( .A1(G63), .A2(n644), .ZN(n571) );
  NAND2_X1 U641 ( .A1(G51), .A2(n656), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U643 ( .A(KEYINPUT6), .B(n572), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n649), .A2(G89), .ZN(n573) );
  XNOR2_X1 U645 ( .A(n573), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U646 ( .A1(G76), .A2(n646), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U648 ( .A(n576), .B(KEYINPUT5), .Z(n577) );
  NOR2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U650 ( .A(KEYINPUT76), .B(n579), .Z(n580) );
  XNOR2_X1 U651 ( .A(KEYINPUT7), .B(n580), .ZN(G168) );
  XOR2_X1 U652 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U653 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U654 ( .A(n581), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U655 ( .A(G223), .B(KEYINPUT73), .ZN(n835) );
  AND2_X1 U656 ( .A1(G567), .A2(n835), .ZN(n582) );
  XNOR2_X1 U657 ( .A(n582), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U658 ( .A1(G56), .A2(n644), .ZN(n583) );
  XOR2_X1 U659 ( .A(KEYINPUT14), .B(n583), .Z(n589) );
  NAND2_X1 U660 ( .A1(n649), .A2(G81), .ZN(n584) );
  XNOR2_X1 U661 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U662 ( .A1(G68), .A2(n646), .ZN(n585) );
  NAND2_X1 U663 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U664 ( .A(KEYINPUT13), .B(n587), .Z(n588) );
  NOR2_X1 U665 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n656), .A2(G43), .ZN(n590) );
  NAND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n916) );
  INV_X1 U668 ( .A(G860), .ZN(n605) );
  OR2_X1 U669 ( .A1(n916), .A2(n605), .ZN(G153) );
  INV_X1 U670 ( .A(G171), .ZN(G301) );
  NAND2_X1 U671 ( .A1(G868), .A2(G301), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G79), .A2(n646), .ZN(n593) );
  NAND2_X1 U673 ( .A1(G54), .A2(n656), .ZN(n592) );
  NAND2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U675 ( .A(n594), .B(KEYINPUT75), .ZN(n596) );
  NAND2_X1 U676 ( .A1(G66), .A2(n644), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n649), .A2(G92), .ZN(n597) );
  XOR2_X1 U679 ( .A(KEYINPUT74), .B(n597), .Z(n598) );
  NOR2_X1 U680 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U681 ( .A(KEYINPUT15), .B(n600), .Z(n921) );
  OR2_X1 U682 ( .A1(n921), .A2(G868), .ZN(n601) );
  NAND2_X1 U683 ( .A1(n602), .A2(n601), .ZN(G284) );
  NAND2_X1 U684 ( .A1(G868), .A2(G286), .ZN(n604) );
  INV_X1 U685 ( .A(G868), .ZN(n668) );
  NAND2_X1 U686 ( .A1(G299), .A2(n668), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U688 ( .A1(n605), .A2(G559), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n606), .A2(n921), .ZN(n607) );
  XNOR2_X1 U690 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U691 ( .A1(G868), .A2(n916), .ZN(n610) );
  NAND2_X1 U692 ( .A1(G868), .A2(n921), .ZN(n608) );
  NOR2_X1 U693 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U694 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G559), .A2(n921), .ZN(n611) );
  XNOR2_X1 U696 ( .A(n611), .B(n916), .ZN(n665) );
  NOR2_X1 U697 ( .A1(G860), .A2(n665), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G93), .A2(n649), .ZN(n613) );
  NAND2_X1 U699 ( .A1(G67), .A2(n644), .ZN(n612) );
  NAND2_X1 U700 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U701 ( .A1(G80), .A2(n646), .ZN(n615) );
  NAND2_X1 U702 ( .A1(G55), .A2(n656), .ZN(n614) );
  NAND2_X1 U703 ( .A1(n615), .A2(n614), .ZN(n616) );
  OR2_X1 U704 ( .A1(n617), .A2(n616), .ZN(n667) );
  XOR2_X1 U705 ( .A(n667), .B(KEYINPUT78), .Z(n618) );
  XNOR2_X1 U706 ( .A(n619), .B(n618), .ZN(G145) );
  NAND2_X1 U707 ( .A1(G49), .A2(n656), .ZN(n621) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n620) );
  NAND2_X1 U709 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U710 ( .A1(n644), .A2(n622), .ZN(n623) );
  XOR2_X1 U711 ( .A(KEYINPUT79), .B(n623), .Z(n626) );
  NAND2_X1 U712 ( .A1(n624), .A2(G87), .ZN(n625) );
  NAND2_X1 U713 ( .A1(n626), .A2(n625), .ZN(G288) );
  NAND2_X1 U714 ( .A1(G85), .A2(n649), .ZN(n628) );
  NAND2_X1 U715 ( .A1(G72), .A2(n646), .ZN(n627) );
  NAND2_X1 U716 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U717 ( .A1(G47), .A2(n656), .ZN(n629) );
  XOR2_X1 U718 ( .A(KEYINPUT70), .B(n629), .Z(n630) );
  NOR2_X1 U719 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n644), .A2(G60), .ZN(n632) );
  NAND2_X1 U721 ( .A1(n633), .A2(n632), .ZN(G290) );
  NAND2_X1 U722 ( .A1(G88), .A2(n649), .ZN(n634) );
  XNOR2_X1 U723 ( .A(n634), .B(KEYINPUT86), .ZN(n637) );
  NAND2_X1 U724 ( .A1(G75), .A2(n646), .ZN(n635) );
  XOR2_X1 U725 ( .A(KEYINPUT87), .B(n635), .Z(n636) );
  NAND2_X1 U726 ( .A1(n637), .A2(n636), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(G62), .ZN(n638) );
  XNOR2_X1 U728 ( .A(n638), .B(KEYINPUT84), .ZN(n640) );
  NAND2_X1 U729 ( .A1(G50), .A2(n656), .ZN(n639) );
  NAND2_X1 U730 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U731 ( .A(KEYINPUT85), .B(n641), .Z(n642) );
  NOR2_X1 U732 ( .A1(n643), .A2(n642), .ZN(G166) );
  INV_X1 U733 ( .A(G166), .ZN(G303) );
  NAND2_X1 U734 ( .A1(n644), .A2(G61), .ZN(n645) );
  XNOR2_X1 U735 ( .A(KEYINPUT80), .B(n645), .ZN(n654) );
  XOR2_X1 U736 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n648) );
  NAND2_X1 U737 ( .A1(G73), .A2(n646), .ZN(n647) );
  XNOR2_X1 U738 ( .A(n648), .B(n647), .ZN(n652) );
  NAND2_X1 U739 ( .A1(G86), .A2(n649), .ZN(n650) );
  XNOR2_X1 U740 ( .A(KEYINPUT81), .B(n650), .ZN(n651) );
  NOR2_X1 U741 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U742 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U743 ( .A(n655), .B(KEYINPUT83), .ZN(n658) );
  NAND2_X1 U744 ( .A1(G48), .A2(n656), .ZN(n657) );
  NAND2_X1 U745 ( .A1(n658), .A2(n657), .ZN(G305) );
  XNOR2_X1 U746 ( .A(KEYINPUT88), .B(G299), .ZN(n659) );
  XNOR2_X1 U747 ( .A(n659), .B(G288), .ZN(n660) );
  XNOR2_X1 U748 ( .A(KEYINPUT19), .B(n660), .ZN(n662) );
  XOR2_X1 U749 ( .A(G290), .B(n667), .Z(n661) );
  XNOR2_X1 U750 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U751 ( .A(n663), .B(G303), .ZN(n664) );
  XNOR2_X1 U752 ( .A(n664), .B(G305), .ZN(n901) );
  XNOR2_X1 U753 ( .A(n665), .B(n901), .ZN(n666) );
  NAND2_X1 U754 ( .A1(n666), .A2(G868), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U756 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n672), .ZN(n674) );
  XOR2_X1 U760 ( .A(KEYINPUT21), .B(KEYINPUT89), .Z(n673) );
  XNOR2_X1 U761 ( .A(n674), .B(n673), .ZN(n675) );
  NAND2_X1 U762 ( .A1(G2072), .A2(n675), .ZN(G158) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U764 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U765 ( .A1(G220), .A2(G219), .ZN(n676) );
  XNOR2_X1 U766 ( .A(KEYINPUT22), .B(n676), .ZN(n677) );
  NAND2_X1 U767 ( .A1(n677), .A2(G96), .ZN(n678) );
  NOR2_X1 U768 ( .A1(G218), .A2(n678), .ZN(n679) );
  XOR2_X1 U769 ( .A(KEYINPUT90), .B(n679), .Z(n839) );
  NAND2_X1 U770 ( .A1(n839), .A2(G2106), .ZN(n680) );
  XNOR2_X1 U771 ( .A(n680), .B(KEYINPUT91), .ZN(n684) );
  NOR2_X1 U772 ( .A1(G236), .A2(G238), .ZN(n681) );
  NAND2_X1 U773 ( .A1(G69), .A2(n681), .ZN(n682) );
  OR2_X1 U774 ( .A1(G237), .A2(n682), .ZN(n840) );
  AND2_X1 U775 ( .A1(G567), .A2(n840), .ZN(n683) );
  NOR2_X1 U776 ( .A1(n684), .A2(n683), .ZN(G319) );
  INV_X1 U777 ( .A(G319), .ZN(n686) );
  NAND2_X1 U778 ( .A1(G483), .A2(G661), .ZN(n685) );
  NOR2_X1 U779 ( .A1(n686), .A2(n685), .ZN(n838) );
  NAND2_X1 U780 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U781 ( .A1(n689), .A2(G40), .ZN(n787) );
  NOR2_X1 U782 ( .A1(n786), .A2(n787), .ZN(n690) );
  XNOR2_X1 U783 ( .A(n690), .B(KEYINPUT64), .ZN(n692) );
  BUF_X1 U784 ( .A(n692), .Z(n711) );
  INV_X1 U785 ( .A(G1961), .ZN(n691) );
  OR2_X1 U786 ( .A1(n711), .A2(n691), .ZN(n694) );
  XOR2_X1 U787 ( .A(G2078), .B(KEYINPUT25), .Z(n970) );
  NAND2_X1 U788 ( .A1(n970), .A2(n711), .ZN(n693) );
  NAND2_X1 U789 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U790 ( .A(KEYINPUT98), .B(n695), .Z(n730) );
  XOR2_X1 U791 ( .A(KEYINPUT102), .B(n696), .Z(n702) );
  NAND2_X1 U792 ( .A1(n704), .A2(G8), .ZN(n784) );
  NOR2_X1 U793 ( .A1(G1966), .A2(n784), .ZN(n750) );
  NOR2_X1 U794 ( .A1(n704), .A2(G2084), .ZN(n746) );
  NOR2_X1 U795 ( .A1(n750), .A2(n746), .ZN(n697) );
  NAND2_X1 U796 ( .A1(G8), .A2(n697), .ZN(n698) );
  XNOR2_X1 U797 ( .A(n698), .B(KEYINPUT30), .ZN(n699) );
  NOR2_X1 U798 ( .A1(G168), .A2(n699), .ZN(n700) );
  XNOR2_X1 U799 ( .A(n700), .B(KEYINPUT101), .ZN(n701) );
  NAND2_X1 U800 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U801 ( .A(n703), .B(KEYINPUT31), .ZN(n734) );
  INV_X1 U802 ( .A(G2072), .ZN(n965) );
  NOR2_X1 U803 ( .A1(n704), .A2(n965), .ZN(n706) );
  XOR2_X1 U804 ( .A(KEYINPUT27), .B(KEYINPUT99), .Z(n705) );
  XNOR2_X1 U805 ( .A(n706), .B(n705), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n704), .A2(G1956), .ZN(n707) );
  NAND2_X1 U807 ( .A1(n708), .A2(n707), .ZN(n725) );
  INV_X1 U808 ( .A(KEYINPUT100), .ZN(n709) );
  XNOR2_X1 U809 ( .A(n710), .B(n709), .ZN(n717) );
  NAND2_X1 U810 ( .A1(n711), .A2(G1996), .ZN(n712) );
  XNOR2_X1 U811 ( .A(n712), .B(KEYINPUT26), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n704), .A2(G1341), .ZN(n713) );
  NAND2_X1 U813 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U814 ( .A1(n921), .A2(n718), .ZN(n716) );
  NAND2_X1 U815 ( .A1(n717), .A2(n716), .ZN(n724) );
  NOR2_X1 U816 ( .A1(n921), .A2(n718), .ZN(n722) );
  NAND2_X1 U817 ( .A1(G2067), .A2(n711), .ZN(n720) );
  NAND2_X1 U818 ( .A1(n704), .A2(G1348), .ZN(n719) );
  NAND2_X1 U819 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U820 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U821 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U822 ( .A1(G299), .A2(n725), .ZN(n726) );
  XOR2_X1 U823 ( .A(KEYINPUT28), .B(n726), .Z(n727) );
  NOR2_X1 U824 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U825 ( .A(n729), .B(KEYINPUT29), .ZN(n732) );
  NAND2_X1 U826 ( .A1(G171), .A2(n730), .ZN(n731) );
  NAND2_X1 U827 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U828 ( .A1(n734), .A2(n733), .ZN(n745) );
  AND2_X1 U829 ( .A1(G286), .A2(G8), .ZN(n735) );
  NAND2_X1 U830 ( .A1(n745), .A2(n735), .ZN(n742) );
  INV_X1 U831 ( .A(G8), .ZN(n740) );
  NOR2_X1 U832 ( .A1(n704), .A2(G2090), .ZN(n737) );
  NOR2_X1 U833 ( .A1(G1971), .A2(n784), .ZN(n736) );
  NOR2_X1 U834 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U835 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U836 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U837 ( .A1(n742), .A2(n741), .ZN(n743) );
  INV_X1 U838 ( .A(KEYINPUT103), .ZN(n744) );
  XNOR2_X1 U839 ( .A(n745), .B(n744), .ZN(n748) );
  NAND2_X1 U840 ( .A1(n746), .A2(G8), .ZN(n747) );
  NAND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U842 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U844 ( .A(n753), .B(KEYINPUT104), .ZN(n771) );
  NAND2_X1 U845 ( .A1(G166), .A2(G8), .ZN(n754) );
  NOR2_X1 U846 ( .A1(G2090), .A2(n754), .ZN(n762) );
  XOR2_X1 U847 ( .A(G1981), .B(KEYINPUT107), .Z(n755) );
  XNOR2_X1 U848 ( .A(G305), .B(n755), .ZN(n928) );
  INV_X1 U849 ( .A(KEYINPUT33), .ZN(n759) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n756) );
  XNOR2_X1 U851 ( .A(KEYINPUT105), .B(n756), .ZN(n770) );
  OR2_X1 U852 ( .A1(n784), .A2(n770), .ZN(n757) );
  NOR2_X1 U853 ( .A1(n759), .A2(n757), .ZN(n758) );
  XOR2_X1 U854 ( .A(n758), .B(KEYINPUT106), .Z(n773) );
  INV_X1 U855 ( .A(n773), .ZN(n760) );
  OR2_X1 U856 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U857 ( .A1(n928), .A2(n761), .ZN(n764) );
  OR2_X1 U858 ( .A1(n762), .A2(n764), .ZN(n763) );
  NOR2_X1 U859 ( .A1(n771), .A2(n763), .ZN(n768) );
  INV_X1 U860 ( .A(n764), .ZN(n766) );
  INV_X1 U861 ( .A(n784), .ZN(n765) );
  AND2_X1 U862 ( .A1(n766), .A2(n765), .ZN(n767) );
  OR2_X1 U863 ( .A1(G303), .A2(G1971), .ZN(n769) );
  NAND2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n935) );
  NOR2_X1 U865 ( .A1(n771), .A2(n935), .ZN(n772) );
  NAND2_X1 U866 ( .A1(G1976), .A2(G288), .ZN(n919) );
  AND2_X1 U867 ( .A1(n919), .A2(n773), .ZN(n775) );
  INV_X1 U868 ( .A(n928), .ZN(n774) );
  AND2_X1 U869 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U871 ( .A1(G1981), .A2(G305), .ZN(n781) );
  XNOR2_X1 U872 ( .A(n781), .B(KEYINPUT97), .ZN(n782) );
  XNOR2_X1 U873 ( .A(KEYINPUT24), .B(n782), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n785), .A2(n510), .ZN(n819) );
  NOR2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n830) );
  XNOR2_X1 U876 ( .A(KEYINPUT37), .B(G2067), .ZN(n828) );
  NAND2_X1 U877 ( .A1(n885), .A2(G104), .ZN(n790) );
  NAND2_X1 U878 ( .A1(G140), .A2(n886), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U880 ( .A(KEYINPUT34), .B(n791), .ZN(n796) );
  NAND2_X1 U881 ( .A1(G116), .A2(n889), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G128), .A2(n890), .ZN(n792) );
  NAND2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U884 ( .A(n794), .B(KEYINPUT35), .Z(n795) );
  NOR2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U886 ( .A(KEYINPUT36), .B(n797), .Z(n798) );
  XNOR2_X1 U887 ( .A(KEYINPUT93), .B(n798), .ZN(n898) );
  NOR2_X1 U888 ( .A1(n828), .A2(n898), .ZN(n991) );
  NAND2_X1 U889 ( .A1(n830), .A2(n991), .ZN(n826) );
  INV_X1 U890 ( .A(n826), .ZN(n816) );
  NAND2_X1 U891 ( .A1(G107), .A2(n889), .ZN(n800) );
  NAND2_X1 U892 ( .A1(G119), .A2(n890), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U894 ( .A(KEYINPUT94), .B(n801), .ZN(n805) );
  NAND2_X1 U895 ( .A1(n885), .A2(G95), .ZN(n803) );
  NAND2_X1 U896 ( .A1(G131), .A2(n886), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n881) );
  XNOR2_X1 U899 ( .A(KEYINPUT95), .B(G1991), .ZN(n969) );
  NOR2_X1 U900 ( .A1(n881), .A2(n969), .ZN(n814) );
  NAND2_X1 U901 ( .A1(n890), .A2(G129), .ZN(n807) );
  NAND2_X1 U902 ( .A1(G141), .A2(n886), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n885), .A2(G105), .ZN(n808) );
  XOR2_X1 U905 ( .A(KEYINPUT38), .B(n808), .Z(n809) );
  NOR2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n889), .A2(G117), .ZN(n811) );
  NAND2_X1 U908 ( .A1(n812), .A2(n811), .ZN(n868) );
  AND2_X1 U909 ( .A1(n868), .A2(G1996), .ZN(n813) );
  NOR2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n993) );
  INV_X1 U911 ( .A(n830), .ZN(n815) );
  NOR2_X1 U912 ( .A1(n993), .A2(n815), .ZN(n823) );
  NOR2_X1 U913 ( .A1(n816), .A2(n823), .ZN(n817) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n913) );
  NAND2_X1 U915 ( .A1(n913), .A2(n830), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n819), .A2(n512), .ZN(n833) );
  NOR2_X1 U917 ( .A1(G1996), .A2(n868), .ZN(n998) );
  AND2_X1 U918 ( .A1(n969), .A2(n881), .ZN(n987) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U920 ( .A1(n987), .A2(n820), .ZN(n821) );
  XOR2_X1 U921 ( .A(KEYINPUT109), .B(n821), .Z(n822) );
  NOR2_X1 U922 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U923 ( .A1(n998), .A2(n824), .ZN(n825) );
  XNOR2_X1 U924 ( .A(KEYINPUT39), .B(n825), .ZN(n827) );
  NAND2_X1 U925 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U926 ( .A1(n828), .A2(n898), .ZN(n995) );
  NAND2_X1 U927 ( .A1(n829), .A2(n995), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U929 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U930 ( .A(n834), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U933 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U935 ( .A1(n838), .A2(n837), .ZN(G188) );
  XNOR2_X1 U936 ( .A(G96), .B(KEYINPUT111), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  XOR2_X1 U940 ( .A(KEYINPUT41), .B(G1956), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1981), .B(G1966), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n843), .B(KEYINPUT113), .Z(n845) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n847) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1961), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U950 ( .A(KEYINPUT114), .B(G2474), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(G229) );
  XOR2_X1 U952 ( .A(G2096), .B(KEYINPUT43), .Z(n853) );
  XNOR2_X1 U953 ( .A(G2090), .B(KEYINPUT112), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(n854), .B(G2678), .Z(n856) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U958 ( .A(KEYINPUT42), .B(G2100), .Z(n858) );
  XNOR2_X1 U959 ( .A(G2084), .B(G2078), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(G227) );
  NAND2_X1 U962 ( .A1(G124), .A2(n890), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n885), .A2(G100), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U966 ( .A1(n889), .A2(G112), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G136), .A2(n886), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U969 ( .A1(n867), .A2(n866), .ZN(G162) );
  XOR2_X1 U970 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n870) );
  XOR2_X1 U971 ( .A(G160), .B(n868), .Z(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n880) );
  NAND2_X1 U973 ( .A1(n885), .A2(G106), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G142), .A2(n886), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n873), .B(KEYINPUT45), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G118), .A2(n889), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G130), .A2(n890), .ZN(n876) );
  XNOR2_X1 U980 ( .A(KEYINPUT115), .B(n876), .ZN(n877) );
  NOR2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U982 ( .A(n880), .B(n879), .Z(n883) );
  XNOR2_X1 U983 ( .A(G164), .B(n881), .ZN(n882) );
  XNOR2_X1 U984 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n988), .B(n884), .ZN(n897) );
  NAND2_X1 U986 ( .A1(n885), .A2(G103), .ZN(n888) );
  NAND2_X1 U987 ( .A1(G139), .A2(n886), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n895) );
  NAND2_X1 U989 ( .A1(G115), .A2(n889), .ZN(n892) );
  NAND2_X1 U990 ( .A1(G127), .A2(n890), .ZN(n891) );
  NAND2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n893), .Z(n894) );
  NOR2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n1003) );
  XNOR2_X1 U994 ( .A(n1003), .B(G162), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n899) );
  XOR2_X1 U996 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U997 ( .A1(G37), .A2(n900), .ZN(G395) );
  XNOR2_X1 U998 ( .A(n916), .B(n901), .ZN(n903) );
  XNOR2_X1 U999 ( .A(G171), .B(n921), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1001 ( .A(n904), .B(G286), .Z(n905) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n905), .ZN(G397) );
  NOR2_X1 U1003 ( .A1(G229), .A2(G227), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n908), .ZN(n909) );
  AND2_X1 U1007 ( .A1(G319), .A2(n909), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1012 ( .A(G1956), .B(G299), .ZN(n912) );
  NOR2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(G1971), .A2(G303), .ZN(n914) );
  NAND2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(G1341), .B(n916), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n926) );
  XOR2_X1 U1019 ( .A(G1348), .B(n921), .Z(n923) );
  XOR2_X1 U1020 ( .A(G171), .B(G1961), .Z(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(n924), .B(KEYINPUT123), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n933) );
  XNOR2_X1 U1024 ( .A(G1966), .B(KEYINPUT121), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(n927), .B(G168), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n931) );
  XOR2_X1 U1027 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n930) );
  XNOR2_X1 U1028 ( .A(n931), .B(n930), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1031 ( .A(KEYINPUT124), .B(n936), .Z(n938) );
  XNOR2_X1 U1032 ( .A(G16), .B(KEYINPUT56), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n1017) );
  XOR2_X1 U1034 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n945) );
  XNOR2_X1 U1035 ( .A(G1971), .B(G22), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(G23), .B(G1976), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1038 ( .A(G1986), .B(KEYINPUT126), .Z(n941) );
  XNOR2_X1 U1039 ( .A(G24), .B(n941), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(n945), .B(n944), .ZN(n960) );
  XOR2_X1 U1042 ( .A(G1348), .B(KEYINPUT59), .Z(n946) );
  XNOR2_X1 U1043 ( .A(G4), .B(n946), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G6), .B(G1981), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G1341), .B(G19), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(G1956), .B(G20), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(n953), .B(KEYINPUT60), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(KEYINPUT125), .B(n954), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G1966), .B(G21), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(G5), .B(G1961), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(KEYINPUT61), .B(n961), .ZN(n963) );
  INV_X1 U1058 ( .A(G16), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1060 ( .A1(n964), .A2(G11), .ZN(n1015) );
  XNOR2_X1 U1061 ( .A(G33), .B(n965), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n966), .A2(G28), .ZN(n976) );
  XNOR2_X1 U1063 ( .A(G2067), .B(G26), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(G32), .B(G1996), .ZN(n967) );
  NOR2_X1 U1065 ( .A1(n968), .A2(n967), .ZN(n974) );
  XOR2_X1 U1066 ( .A(n969), .B(G25), .Z(n972) );
  XNOR2_X1 U1067 ( .A(G27), .B(n970), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1071 ( .A(KEYINPUT53), .B(n977), .Z(n980) );
  XOR2_X1 U1072 ( .A(G34), .B(KEYINPUT54), .Z(n978) );
  XNOR2_X1 U1073 ( .A(G2084), .B(n978), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(G35), .B(G2090), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT120), .B(n983), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(G29), .A2(n984), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n985), .B(KEYINPUT55), .ZN(n1013) );
  XOR2_X1 U1080 ( .A(G160), .B(G2084), .Z(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(n994), .B(KEYINPUT117), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n1001) );
  XOR2_X1 U1087 ( .A(G2090), .B(G162), .Z(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(n999), .B(KEYINPUT51), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(KEYINPUT118), .B(n1002), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(G2072), .B(n1003), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(n1004), .B(KEYINPUT119), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(G2078), .B(G164), .Z(n1005) );
  NOR2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT52), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(G29), .A2(n1011), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1018), .Z(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

