//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(G355));
  XNOR2_X1  g0007(.A(KEYINPUT66), .B(G238), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(new_n203), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G87), .A2(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n214), .B1(new_n201), .B2(new_n215), .ZN(new_n216));
  NOR3_X1   g0016(.A1(new_n209), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT67), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n217), .A2(new_n219), .B1(G1), .B2(G20), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G20), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n229), .B1(new_n230), .B2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G13), .ZN(new_n232));
  NAND4_X1  g0032(.A1(new_n232), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT0), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n222), .A2(new_n228), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g0037(.A(new_n237), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G250), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n212), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT2), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G226), .ZN(new_n245));
  INV_X1    g0045(.A(G232), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n242), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G68), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n225), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n259), .A2(new_n201), .B1(new_n226), .B2(G68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n226), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G77), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n257), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT11), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT76), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n266), .B1(new_n268), .B2(G68), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT12), .ZN(new_n270));
  INV_X1    g0070(.A(new_n268), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n257), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n203), .B1(new_n267), .B2(G20), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n265), .A2(new_n274), .A3(KEYINPUT77), .ZN(new_n275));
  AOI21_X1  g0075(.A(KEYINPUT77), .B1(new_n265), .B2(new_n274), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT14), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G97), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT75), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT75), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G33), .A3(G97), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n246), .A2(G1698), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n284), .B1(G226), .B2(G1698), .ZN(new_n285));
  AND2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n283), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G238), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  AND2_X1   g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  OAI21_X1  g0099(.A(G274), .B1(new_n299), .B2(new_n225), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT69), .B1(new_n300), .B2(new_n294), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  AND2_X1   g0102(.A1(G1), .A2(G13), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n290), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT69), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(new_n295), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n298), .A2(new_n307), .A3(KEYINPUT13), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT13), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n289), .A2(new_n292), .B1(new_n296), .B2(G238), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n301), .A2(new_n306), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n278), .B(G169), .C1(new_n308), .C2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT13), .B1(new_n298), .B2(new_n307), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(new_n309), .A3(new_n311), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(G179), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n315), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n278), .B1(new_n318), .B2(G169), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n277), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(G200), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n314), .A2(G190), .A3(new_n315), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n321), .A2(new_n274), .A3(new_n265), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT78), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n256), .A2(new_n225), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT8), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G58), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n261), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n330), .A2(new_n331), .B1(G150), .B2(new_n258), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n204), .A2(G20), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n326), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT70), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n201), .B1(new_n267), .B2(G20), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n272), .A2(new_n336), .B1(new_n201), .B2(new_n271), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT9), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n334), .A2(KEYINPUT70), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT9), .B1(new_n338), .B2(new_n341), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT3), .B(G33), .ZN(new_n346));
  INV_X1    g0146(.A(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G222), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G223), .A2(G1698), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n292), .C1(G77), .C2(new_n346), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n296), .A2(G226), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n311), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G200), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n354), .B2(G190), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n345), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT74), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT10), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n345), .A2(new_n357), .A3(new_n360), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n339), .A2(new_n342), .B1(new_n364), .B2(new_n353), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n365), .A2(KEYINPUT71), .ZN(new_n366));
  INV_X1    g0166(.A(G179), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n365), .A2(KEYINPUT71), .B1(new_n367), .B2(new_n354), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n362), .A2(new_n363), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n346), .B1(new_n246), .B2(G1698), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n208), .A2(new_n347), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n292), .B1(G107), .B2(new_n346), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n296), .A2(G244), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(G190), .A3(new_n311), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT72), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n311), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G200), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n374), .A2(new_n307), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(KEYINPUT72), .A3(G190), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n267), .A2(G20), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n272), .A2(G77), .A3(new_n383), .ZN(new_n384));
  XOR2_X1   g0184(.A(new_n384), .B(KEYINPUT73), .Z(new_n385));
  NAND2_X1  g0185(.A1(new_n271), .A2(new_n262), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT15), .B(G87), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n387), .A2(new_n261), .B1(new_n226), .B2(new_n262), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n259), .B1(new_n327), .B2(new_n329), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n257), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n385), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n378), .A2(new_n380), .A3(new_n382), .A4(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n385), .A2(new_n386), .A3(new_n390), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n379), .B2(G179), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n381), .A2(G169), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n325), .A2(new_n369), .A3(new_n392), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n346), .B2(G20), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n203), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n202), .A2(new_n203), .ZN(new_n403));
  NOR2_X1   g0203(.A1(G58), .A2(G68), .ZN(new_n404));
  OAI21_X1  g0204(.A(G20), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n258), .A2(G159), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n398), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT7), .B1(new_n288), .B2(new_n226), .ZN(new_n409));
  NOR4_X1   g0209(.A1(new_n286), .A2(new_n287), .A3(new_n399), .A4(G20), .ZN(new_n410));
  OAI21_X1  g0210(.A(G68), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n407), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(KEYINPUT16), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n408), .A2(new_n413), .A3(new_n257), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n326), .A2(new_n268), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n330), .A2(new_n383), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n415), .A2(new_n416), .B1(new_n268), .B2(new_n330), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT79), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  OR2_X1    g0219(.A1(G223), .A2(G1698), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n215), .A2(G1698), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(new_n286), .C2(new_n287), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G87), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n306), .A2(new_n301), .B1(new_n424), .B2(new_n292), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n291), .A2(G232), .A3(new_n294), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT80), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n291), .A2(new_n294), .A3(KEYINPUT80), .A4(G232), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(G169), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n424), .A2(new_n292), .ZN(new_n432));
  AND4_X1   g0232(.A1(new_n367), .A2(new_n430), .A3(new_n311), .A4(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n419), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n419), .B2(new_n434), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(G200), .B1(new_n425), .B2(new_n430), .ZN(new_n440));
  INV_X1    g0240(.A(G190), .ZN(new_n441));
  AND4_X1   g0241(.A1(new_n441), .A2(new_n430), .A3(new_n311), .A4(new_n432), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT17), .B1(new_n419), .B2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n430), .A2(new_n311), .A3(new_n432), .A4(new_n441), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n430), .A2(new_n311), .A3(new_n432), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n445), .B1(new_n446), .B2(G200), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT17), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n414), .A4(new_n418), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n444), .A2(KEYINPUT81), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT81), .B1(new_n444), .B2(new_n449), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n439), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n324), .A2(KEYINPUT78), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n397), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n267), .A2(G33), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n272), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G107), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT88), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n268), .A2(G107), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(KEYINPUT25), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT25), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n268), .B2(G107), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n456), .A2(new_n457), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n460), .A2(new_n462), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n226), .B(G87), .C1(new_n286), .C2(new_n287), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT22), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT22), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n346), .A2(new_n468), .A3(new_n226), .A4(G87), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(KEYINPUT86), .A2(KEYINPUT23), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT85), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT86), .B1(new_n473), .B2(KEYINPUT23), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n226), .A2(G107), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n471), .B(new_n472), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  OR2_X1    g0276(.A1(KEYINPUT86), .A2(KEYINPUT23), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n457), .A2(G20), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n470), .A2(new_n480), .A3(KEYINPUT87), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(KEYINPUT24), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT87), .B1(new_n470), .B2(new_n480), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT24), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n326), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n465), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G45), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G1), .ZN(new_n491));
  INV_X1    g0291(.A(G41), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT5), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT5), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G41), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n496), .A2(G264), .A3(new_n291), .ZN(new_n497));
  AND2_X1   g0297(.A1(G257), .A2(G1698), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n286), .B2(new_n287), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT89), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n346), .A2(G250), .A3(new_n347), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G294), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT89), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n498), .C1(new_n286), .C2(new_n287), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n497), .B1(new_n505), .B2(new_n292), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n304), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n367), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n496), .A2(new_n300), .ZN(new_n510));
  AOI211_X1 g0310(.A(new_n510), .B(new_n497), .C1(new_n505), .C2(new_n292), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n509), .B1(new_n511), .B2(G169), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n484), .A2(KEYINPUT24), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(new_n486), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n481), .A2(new_n482), .A3(new_n487), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n257), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n505), .A2(new_n292), .ZN(new_n518));
  INV_X1    g0318(.A(new_n497), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n518), .A2(G190), .A3(new_n508), .A4(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n463), .A2(new_n464), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n521), .C1(new_n511), .C2(new_n355), .ZN(new_n522));
  OAI22_X1  g0322(.A1(new_n489), .A2(new_n512), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G116), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n271), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n326), .A2(G116), .A3(new_n268), .A4(new_n455), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n256), .A2(new_n225), .B1(G20), .B2(new_n525), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G283), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n529), .B(new_n226), .C1(G33), .C2(new_n211), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n528), .A2(KEYINPUT20), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT20), .B1(new_n528), .B2(new_n530), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n526), .B(new_n527), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n347), .A2(G257), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G264), .A2(G1698), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n534), .B(new_n535), .C1(new_n286), .C2(new_n287), .ZN(new_n536));
  OR2_X1    g0336(.A1(KEYINPUT3), .A2(G33), .ZN(new_n537));
  INV_X1    g0337(.A(G303), .ZN(new_n538));
  NAND2_X1  g0338(.A1(KEYINPUT3), .A2(G33), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n536), .A2(new_n292), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n496), .A2(G270), .A3(new_n291), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n508), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n533), .A2(KEYINPUT21), .A3(G169), .A4(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT84), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n291), .B1(new_n288), .B2(new_n538), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n536), .B1(new_n507), .B2(new_n304), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n364), .B1(new_n548), .B2(new_n542), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n549), .A2(KEYINPUT84), .A3(KEYINPUT21), .A4(new_n533), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n533), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT21), .ZN(new_n553));
  AND4_X1   g0353(.A1(G179), .A2(new_n508), .A3(new_n541), .A4(new_n542), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n552), .A2(new_n553), .B1(new_n533), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n533), .B1(G200), .B2(new_n543), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n441), .B2(new_n543), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n551), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n346), .A2(new_n226), .A3(G68), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n261), .A2(new_n211), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n560), .B1(KEYINPUT19), .B2(new_n561), .ZN(new_n562));
  NOR3_X1   g0362(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n280), .A2(new_n282), .A3(KEYINPUT19), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n563), .B1(new_n564), .B2(new_n226), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n257), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n387), .A2(new_n271), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n566), .B(new_n567), .C1(new_n387), .C2(new_n456), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n267), .A2(G45), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n291), .A2(G250), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G238), .A2(G1698), .ZN(new_n571));
  INV_X1    g0371(.A(G244), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(G1698), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n346), .B1(G33), .B2(G116), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n570), .B1(new_n574), .B2(new_n291), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT82), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n304), .B2(new_n491), .ZN(new_n577));
  AND4_X1   g0377(.A1(new_n576), .A2(new_n291), .A3(G274), .A4(new_n491), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT83), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n570), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G116), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n572), .A2(G1698), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(G238), .B2(G1698), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n582), .B1(new_n584), .B2(new_n288), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n581), .B1(new_n585), .B2(new_n292), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT83), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT82), .B1(new_n300), .B2(new_n569), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n304), .A2(new_n576), .A3(new_n491), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n580), .A2(new_n367), .A3(new_n591), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n575), .A2(new_n579), .A3(KEYINPUT83), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n587), .B1(new_n586), .B2(new_n590), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n568), .B(new_n592), .C1(new_n595), .C2(G169), .ZN(new_n596));
  OAI21_X1  g0396(.A(G200), .B1(new_n593), .B2(new_n594), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n580), .A2(G190), .A3(new_n591), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n272), .A2(G87), .A3(new_n455), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n566), .A2(new_n567), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT4), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(G1698), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n603), .B(G244), .C1(new_n287), .C2(new_n286), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n572), .B1(new_n537), .B2(new_n539), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n604), .B(new_n529), .C1(new_n605), .C2(KEYINPUT4), .ZN(new_n606));
  OAI21_X1  g0406(.A(G250), .B1(new_n286), .B2(new_n287), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n347), .B1(new_n607), .B2(KEYINPUT4), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n292), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n507), .A2(new_n292), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n510), .B1(new_n610), .B2(G257), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n355), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n611), .A3(new_n441), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n268), .A2(G97), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n456), .B2(new_n211), .ZN(new_n618));
  OAI21_X1  g0418(.A(G107), .B1(new_n409), .B2(new_n410), .ZN(new_n619));
  XNOR2_X1  g0419(.A(G97), .B(G107), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT6), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n621), .A2(new_n211), .A3(G107), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G20), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n258), .A2(G77), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n619), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n618), .B1(new_n628), .B2(new_n257), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n615), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n623), .B1(new_n621), .B2(new_n620), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n627), .B1(new_n631), .B2(new_n226), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n457), .B1(new_n400), .B2(new_n401), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n257), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n618), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n609), .A2(new_n611), .A3(G179), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n364), .B1(new_n609), .B2(new_n611), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n596), .A2(new_n601), .A3(new_n630), .A4(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n454), .A2(new_n524), .A3(new_n559), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT90), .ZN(G372));
  NAND2_X1  g0444(.A1(new_n586), .A2(new_n590), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n364), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n592), .A2(new_n568), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(G200), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n598), .A2(new_n600), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n551), .B(new_n555), .C1(new_n489), .C2(new_n512), .ZN(new_n651));
  INV_X1    g0451(.A(new_n522), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n485), .A2(new_n488), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n612), .A2(G169), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n629), .B1(new_n655), .B2(new_n637), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n636), .B1(new_n613), .B2(new_n614), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n650), .A2(new_n651), .A3(new_n654), .A4(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT91), .B1(new_n638), .B2(new_n639), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT91), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n655), .A2(new_n661), .A3(new_n637), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n629), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT26), .B1(new_n650), .B2(new_n663), .ZN(new_n664));
  AND4_X1   g0464(.A1(KEYINPUT26), .A2(new_n596), .A3(new_n656), .A4(new_n601), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n659), .B(new_n647), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n454), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n396), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n323), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(new_n320), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT81), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT79), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n417), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n411), .A2(new_n412), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n326), .B1(new_n674), .B2(new_n398), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n673), .B1(new_n413), .B2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n448), .B1(new_n676), .B2(new_n447), .ZN(new_n677));
  INV_X1    g0477(.A(new_n449), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n671), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n444), .A2(KEYINPUT81), .A3(new_n449), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n439), .B1(new_n670), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n362), .A2(new_n363), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n683), .A2(new_n685), .B1(new_n366), .B2(new_n368), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n667), .A2(new_n686), .ZN(G369));
  AND2_X1   g0487(.A1(new_n551), .A2(new_n555), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n267), .A2(new_n226), .A3(G13), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n512), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n521), .B1(new_n514), .B2(new_n516), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(new_n694), .ZN(new_n699));
  INV_X1    g0499(.A(new_n694), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n489), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n699), .B1(new_n523), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT92), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT92), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n704), .B(new_n699), .C1(new_n523), .C2(new_n701), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n696), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n697), .A2(new_n698), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n694), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT93), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n705), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n698), .A2(new_n694), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n654), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n704), .B1(new_n712), .B2(new_n699), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n695), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT93), .ZN(new_n715));
  INV_X1    g0515(.A(new_n708), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n709), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n710), .A2(new_n713), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n533), .A2(new_n694), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n559), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n688), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n718), .A2(new_n725), .ZN(G399));
  NAND2_X1  g0526(.A1(new_n563), .A2(new_n525), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT94), .ZN(new_n728));
  INV_X1    g0528(.A(new_n234), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G41), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n728), .A2(new_n730), .A3(new_n267), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n224), .B2(new_n730), .ZN(new_n732));
  XNOR2_X1  g0532(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n666), .A2(new_n700), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT29), .ZN(new_n737));
  INV_X1    g0537(.A(new_n650), .ZN(new_n738));
  INV_X1    g0538(.A(new_n663), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT26), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT26), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n596), .A2(new_n601), .A3(new_n741), .A4(new_n656), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n740), .A2(new_n742), .A3(new_n647), .A4(new_n659), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n737), .B1(new_n743), .B2(new_n700), .ZN(new_n744));
  INV_X1    g0544(.A(G330), .ZN(new_n745));
  AND4_X1   g0545(.A1(new_n506), .A2(new_n554), .A3(new_n609), .A4(new_n611), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n595), .A2(new_n746), .A3(KEYINPUT30), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n580), .A2(new_n591), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n506), .A2(new_n554), .A3(new_n609), .A4(new_n611), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n506), .A2(new_n508), .ZN(new_n752));
  AOI21_X1  g0552(.A(G179), .B1(new_n548), .B2(new_n542), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n752), .A2(new_n612), .A3(new_n645), .A4(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n747), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n694), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(KEYINPUT31), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n755), .A2(new_n758), .A3(new_n694), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n642), .A2(new_n524), .A3(new_n559), .A4(new_n700), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n745), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OR3_X1    g0562(.A1(new_n736), .A2(new_n744), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n734), .B1(new_n764), .B2(G1), .ZN(G364));
  INV_X1    g0565(.A(new_n723), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n226), .A2(G13), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT96), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n490), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n267), .B1(new_n770), .B2(KEYINPUT97), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(KEYINPUT97), .B2(new_n770), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n730), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(G330), .B2(new_n722), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n225), .B1(G20), .B2(new_n364), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n729), .A2(new_n346), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G45), .B2(new_n223), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(G45), .B2(new_n251), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n729), .A2(new_n288), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G355), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G116), .B2(new_n234), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n780), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n773), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n226), .A2(G190), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(new_n367), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT100), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G107), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G179), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n789), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n789), .A2(G179), .A3(new_n355), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT98), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n796), .B(new_n802), .C1(new_n262), .C2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G190), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT101), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n810), .A2(new_n811), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n203), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n226), .A2(new_n441), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n817), .A2(new_n367), .A3(G200), .ZN(new_n818));
  INV_X1    g0618(.A(G87), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n817), .A2(G179), .A3(new_n355), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n346), .B1(new_n818), .B2(new_n819), .C1(new_n202), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n809), .A2(new_n441), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n226), .B1(new_n797), .B2(G190), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n823), .A2(new_n201), .B1(new_n824), .B2(new_n211), .ZN(new_n825));
  NOR4_X1   g0625(.A1(new_n808), .A2(new_n816), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n827), .A2(KEYINPUT102), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(KEYINPUT102), .ZN(new_n829));
  INV_X1    g0629(.A(new_n815), .ZN(new_n830));
  XNOR2_X1  g0630(.A(KEYINPUT33), .B(G317), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n798), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G329), .ZN(new_n834));
  INV_X1    g0634(.A(new_n820), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n346), .B1(new_n835), .B2(G322), .ZN(new_n836));
  INV_X1    g0636(.A(new_n824), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G294), .B1(G326), .B2(new_n822), .ZN(new_n838));
  AND4_X1   g0638(.A1(new_n832), .A2(new_n834), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n807), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n818), .B(KEYINPUT103), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n840), .A2(G311), .B1(new_n841), .B2(G303), .ZN(new_n842));
  INV_X1    g0642(.A(G283), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n839), .B(new_n842), .C1(new_n843), .C2(new_n794), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n828), .A2(new_n829), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n788), .B1(new_n845), .B2(new_n779), .ZN(new_n846));
  INV_X1    g0646(.A(new_n778), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n722), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n775), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G396));
  NOR3_X1   g0650(.A1(new_n394), .A2(new_n395), .A3(new_n694), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n393), .A2(new_n694), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n392), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n851), .B1(new_n853), .B2(new_n396), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n735), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n396), .A2(new_n392), .A3(new_n700), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n666), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n762), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n773), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  INV_X1    g0662(.A(new_n773), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n779), .A2(new_n776), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n262), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n795), .A2(G87), .ZN(new_n866));
  INV_X1    g0666(.A(new_n841), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n866), .B1(new_n457), .B2(new_n867), .C1(new_n525), .C2(new_n807), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n815), .A2(new_n843), .ZN(new_n869));
  INV_X1    g0669(.A(G311), .ZN(new_n870));
  INV_X1    g0670(.A(G294), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n288), .B1(new_n798), .B2(new_n870), .C1(new_n820), .C2(new_n871), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n823), .A2(new_n538), .B1(new_n824), .B2(new_n211), .ZN(new_n873));
  NOR4_X1   g0673(.A1(new_n868), .A2(new_n869), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(G132), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n346), .B1(new_n798), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n795), .A2(G68), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n201), .B2(new_n867), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT104), .Z(new_n879));
  AOI211_X1 g0679(.A(new_n876), .B(new_n879), .C1(G58), .C2(new_n837), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n835), .A2(G143), .B1(G137), .B2(new_n822), .ZN(new_n881));
  INV_X1    g0681(.A(G150), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n881), .B1(new_n815), .B2(new_n882), .C1(new_n807), .C2(new_n799), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT34), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n874), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n779), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n865), .B1(new_n777), .B2(new_n854), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n862), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(G384));
  AND3_X1   g0689(.A1(new_n755), .A2(new_n758), .A3(new_n694), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n758), .B1(new_n755), .B2(new_n694), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR4_X1   g0692(.A1(new_n641), .A2(new_n523), .A3(new_n558), .A4(new_n694), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT109), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT109), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n760), .A2(new_n761), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n454), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT110), .Z(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n277), .A2(new_n694), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n320), .A2(new_n323), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(new_n320), .B2(new_n323), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n854), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n900), .B(new_n904), .C1(new_n894), .C2(new_n896), .ZN(new_n905));
  INV_X1    g0705(.A(new_n692), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n419), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n452), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n419), .A2(new_n434), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT37), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n447), .A2(new_n414), .A3(new_n418), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n910), .A2(new_n907), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT105), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n910), .A2(new_n907), .A3(new_n912), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT37), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n915), .A2(KEYINPUT105), .A3(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n677), .A2(new_n678), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n910), .A2(KEYINPUT18), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n436), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n908), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT107), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n916), .A2(new_n925), .A3(new_n913), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n913), .A2(new_n925), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT38), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n920), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n905), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n904), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT109), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n895), .B1(new_n760), .B2(new_n761), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT106), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n919), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n909), .B2(new_n919), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n917), .A2(new_n918), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n907), .B1(new_n681), .B2(new_n439), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n929), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(KEYINPUT106), .A3(new_n920), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n936), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n932), .B1(new_n945), .B2(KEYINPUT40), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n899), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n899), .A2(new_n946), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(G330), .A3(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT111), .Z(new_n950));
  AOI21_X1  g0750(.A(new_n851), .B1(new_n666), .B2(new_n857), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n902), .A2(new_n903), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n938), .A2(new_n939), .A3(new_n937), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT106), .B1(new_n943), .B2(new_n920), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n320), .A2(new_n694), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT39), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n943), .B2(new_n920), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n920), .A2(new_n930), .A3(new_n959), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n923), .A2(new_n692), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n956), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT108), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n956), .A2(new_n962), .A3(KEYINPUT108), .A4(new_n963), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n454), .B1(new_n736), .B2(new_n744), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n686), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n968), .B(new_n970), .Z(new_n971));
  OR2_X1    g0771(.A1(new_n950), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n768), .A2(G1), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n950), .A2(new_n971), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n976), .A2(G116), .A3(new_n227), .A4(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT36), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n403), .A2(new_n223), .A3(new_n262), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n203), .A2(G50), .ZN(new_n981));
  OAI211_X1 g0781(.A(G1), .B(new_n232), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n975), .A2(new_n979), .A3(new_n982), .ZN(G367));
  OAI21_X1  g0783(.A(new_n658), .B1(new_n629), .B2(new_n700), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n663), .A2(new_n694), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n714), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT42), .ZN(new_n989));
  INV_X1    g0789(.A(new_n707), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n656), .B1(new_n986), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n989), .B1(new_n694), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n650), .B1(new_n600), .B2(new_n700), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n600), .A2(new_n700), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n647), .B2(new_n994), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n992), .A2(KEYINPUT43), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT112), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n995), .B(KEYINPUT43), .Z(new_n999));
  NAND2_X1  g0799(.A1(new_n992), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n725), .A2(new_n987), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n998), .A2(new_n1002), .A3(new_n1000), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n730), .B(KEYINPUT41), .Z(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT45), .B1(new_n718), .B2(new_n986), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT45), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1008), .B(new_n987), .C1(new_n709), .C2(new_n717), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(KEYINPUT44), .B1(new_n718), .B2(new_n986), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n709), .A2(new_n717), .A3(new_n1012), .A4(new_n987), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n724), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n706), .A2(KEYINPUT93), .A3(new_n708), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n715), .B1(new_n714), .B2(new_n716), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n986), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n1008), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n718), .A2(KEYINPUT45), .A3(new_n986), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1021), .A2(new_n725), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n719), .A2(new_n696), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n714), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(new_n766), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n764), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1015), .A2(new_n1022), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT113), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1015), .A2(new_n1022), .A3(new_n1027), .A4(KEYINPUT113), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1006), .B1(new_n1032), .B2(new_n764), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1004), .B(new_n1005), .C1(new_n1033), .C2(new_n772), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n780), .B1(new_n234), .B2(new_n387), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n242), .B2(new_n781), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n824), .A2(new_n203), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n835), .A2(G150), .B1(new_n833), .B2(G137), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(new_n346), .C1(new_n202), .C2(new_n818), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1037), .B(new_n1039), .C1(G143), .C2(new_n822), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n795), .A2(G77), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n807), .A2(new_n201), .B1(new_n815), .B2(new_n799), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1042), .B1(new_n1043), .B2(KEYINPUT115), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(KEYINPUT115), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n841), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n818), .A2(new_n525), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1046), .B1(KEYINPUT46), .B2(new_n1047), .C1(new_n815), .C2(new_n871), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT114), .Z(new_n1049));
  NAND2_X1  g0849(.A1(new_n795), .A2(G97), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n843), .B2(new_n807), .ZN(new_n1051));
  INV_X1    g0851(.A(G317), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n288), .B1(new_n798), .B2(new_n1052), .C1(new_n820), .C2(new_n538), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n823), .A2(new_n870), .B1(new_n824), .B2(new_n457), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1044), .A2(new_n1045), .B1(new_n1049), .B2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT47), .Z(new_n1057));
  AOI211_X1 g0857(.A(new_n863), .B(new_n1036), .C1(new_n1057), .C2(new_n779), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n847), .B2(new_n995), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1034), .A2(new_n1059), .ZN(G387));
  NAND2_X1  g0860(.A1(new_n247), .A2(G45), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1061), .A2(new_n781), .B1(new_n728), .B2(new_n784), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n330), .A2(new_n201), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT50), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n490), .B1(new_n203), .B2(new_n262), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1064), .A2(new_n728), .A3(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1062), .A2(new_n1066), .B1(G107), .B2(new_n234), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n863), .B1(new_n1067), .B2(new_n780), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n824), .A2(new_n387), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n288), .B1(new_n833), .B2(G150), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n818), .A2(new_n262), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n201), .C2(new_n820), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1069), .B(new_n1072), .C1(G159), .C2(new_n822), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n830), .A2(new_n330), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n840), .A2(G68), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1073), .A2(new_n1050), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n346), .B1(new_n833), .B2(G326), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n818), .A2(new_n871), .B1(new_n824), .B2(new_n843), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n835), .A2(G317), .B1(G322), .B2(new_n822), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n815), .B2(new_n870), .C1(new_n807), .C2(new_n538), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT48), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n1081), .B2(new_n1080), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT49), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1077), .B1(new_n525), .B2(new_n794), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1076), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n779), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1068), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n719), .B2(new_n778), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n1025), .B2(new_n772), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1026), .A2(new_n730), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n764), .A2(new_n1025), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(G393));
  INV_X1    g0894(.A(new_n730), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1015), .A2(new_n1022), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1095), .B1(new_n1096), .B2(new_n1026), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1032), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(KEYINPUT116), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT116), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1015), .A2(new_n1022), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1099), .A2(new_n772), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n986), .A2(new_n847), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT117), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n780), .B1(new_n211), .B2(new_n234), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n254), .B2(new_n781), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n815), .A2(new_n538), .B1(new_n525), .B2(new_n824), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT118), .Z(new_n1108));
  OAI22_X1  g0908(.A1(new_n1052), .A2(new_n823), .B1(new_n820), .B2(new_n870), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT52), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n840), .A2(G294), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n818), .A2(new_n843), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n346), .B(new_n1112), .C1(G322), .C2(new_n833), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1110), .A2(new_n1111), .A3(new_n796), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n840), .A2(new_n330), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n818), .A2(new_n203), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n288), .B(new_n1116), .C1(G143), .C2(new_n833), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n837), .A2(G77), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1115), .A2(new_n866), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n835), .A2(G159), .B1(G150), .B2(new_n822), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n830), .A2(G50), .B1(KEYINPUT51), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(KEYINPUT51), .B2(new_n1120), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1108), .A2(new_n1114), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n863), .B(new_n1106), .C1(new_n1123), .C2(new_n779), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1104), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1102), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1098), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(G390));
  OAI21_X1  g0928(.A(new_n957), .B1(new_n951), .B2(new_n952), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT119), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT39), .B1(new_n938), .B2(new_n939), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n920), .A2(new_n930), .A3(new_n959), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT119), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1133), .B(new_n957), .C1(new_n951), .C2(new_n952), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n743), .A2(new_n700), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n853), .A2(new_n396), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n851), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n931), .B(new_n957), .C1(new_n1138), .C2(new_n952), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n897), .A2(G330), .A3(new_n933), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n952), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n762), .A2(new_n1144), .A3(new_n854), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1135), .A2(new_n1139), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n454), .A2(G330), .A3(new_n897), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n969), .A2(new_n1147), .A3(new_n686), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n952), .B1(new_n860), .B2(new_n855), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1141), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n951), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n745), .B(new_n855), .C1(new_n894), .C2(new_n896), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1138), .B(new_n1145), .C1(new_n1153), .C2(new_n1144), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1148), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1143), .A2(new_n1146), .A3(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1156), .A2(new_n730), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1148), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT120), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1146), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1141), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1160), .B(new_n1161), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1161), .B1(new_n1166), .B2(new_n1160), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1157), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1166), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1131), .A2(new_n776), .A3(new_n1132), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n864), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n773), .B1(new_n330), .B2(new_n1171), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n288), .B1(new_n798), .B2(new_n871), .C1(new_n820), .C2(new_n525), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1118), .B1(new_n823), .B2(new_n843), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n830), .C2(G107), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n840), .A2(G97), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n841), .A2(G87), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1175), .A2(new_n877), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n818), .A2(new_n882), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT121), .Z(new_n1180));
  INV_X1    g0980(.A(KEYINPUT53), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1180), .A2(new_n1181), .B1(G137), .B2(new_n830), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n1181), .B2(new_n1180), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n346), .B1(new_n820), .B2(new_n875), .ZN(new_n1184));
  INV_X1    g0984(.A(G128), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n823), .A2(new_n1185), .B1(new_n824), .B2(new_n799), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1184), .B(new_n1186), .C1(G125), .C2(new_n833), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT54), .B(G143), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1187), .B1(new_n201), .B2(new_n794), .C1(new_n807), .C2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1178), .B1(new_n1183), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1172), .B1(new_n1190), .B2(new_n779), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT122), .Z(new_n1192));
  AOI22_X1  g0992(.A1(new_n1169), .A2(new_n772), .B1(new_n1170), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1168), .A2(new_n1193), .ZN(G378));
  NAND2_X1  g0994(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n745), .B1(new_n905), .B2(new_n931), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n945), .B2(KEYINPUT40), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n369), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n906), .B1(new_n338), .B2(new_n341), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n369), .A2(new_n1199), .ZN(new_n1203));
  OR3_X1    g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1202), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1197), .A2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1196), .B(new_n1206), .C1(new_n945), .C2(KEYINPUT40), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n968), .A2(new_n1210), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n966), .A2(new_n1208), .A3(new_n967), .A4(new_n1209), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1195), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT57), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1195), .A2(new_n1211), .A3(KEYINPUT57), .A4(new_n1212), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n730), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1211), .A2(new_n772), .A3(new_n1212), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n288), .A2(new_n492), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n387), .A2(new_n807), .B1(new_n794), .B2(new_n202), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1071), .B1(new_n843), .B2(new_n798), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1219), .B(new_n1222), .C1(G107), .C2(new_n835), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1037), .B1(new_n822), .B2(G116), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1221), .B(new_n1225), .C1(G97), .C2(new_n830), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1220), .B1(new_n1226), .B2(KEYINPUT58), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT123), .Z(new_n1228));
  NOR2_X1   g1028(.A1(new_n824), .A2(new_n882), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1185), .A2(new_n820), .B1(new_n818), .B2(new_n1188), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(G125), .C2(new_n822), .ZN(new_n1231));
  INV_X1    g1031(.A(G137), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1231), .B1(new_n875), .B2(new_n815), .C1(new_n1232), .C2(new_n807), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1234));
  AOI211_X1 g1034(.A(G33), .B(G41), .C1(new_n833), .C2(G124), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n794), .B2(new_n799), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1233), .B2(KEYINPUT59), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1226), .A2(KEYINPUT58), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n886), .B1(new_n1228), .B2(new_n1238), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n863), .B(new_n1239), .C1(new_n201), .C2(new_n864), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1206), .B2(new_n777), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1218), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1217), .A2(new_n1242), .ZN(G375));
  NAND2_X1  g1043(.A1(new_n952), .A2(new_n776), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n773), .B1(G68), .B2(new_n1171), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n807), .A2(new_n457), .B1(new_n815), .B2(new_n525), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT124), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n288), .B1(new_n798), .B2(new_n538), .C1(new_n820), .C2(new_n843), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1069), .B(new_n1248), .C1(G294), .C2(new_n822), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n841), .A2(G97), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1247), .A2(new_n1041), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1246), .A2(KEYINPUT124), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G150), .A2(new_n840), .B1(new_n795), .B2(G58), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n799), .B2(new_n867), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n346), .B1(new_n820), .B2(new_n1232), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G128), .B2(new_n833), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n837), .A2(G50), .B1(G132), .B2(new_n822), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(new_n815), .C2(new_n1188), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n1251), .A2(new_n1252), .B1(new_n1254), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1245), .B1(new_n1259), .B2(new_n779), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1158), .A2(new_n772), .B1(new_n1244), .B2(new_n1260), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1155), .A2(new_n1006), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1262), .B2(new_n1263), .ZN(G381));
  XNOR2_X1  g1064(.A(G375), .B(KEYINPUT125), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1168), .A2(new_n1193), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1034), .A2(new_n1059), .A3(new_n1127), .ZN(new_n1267));
  NOR4_X1   g1067(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(G407));
  NAND2_X1  g1069(.A1(new_n693), .A2(G213), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1265), .A2(new_n1266), .A3(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(G407), .A2(G213), .A3(new_n1272), .ZN(G409));
  NAND3_X1  g1073(.A1(new_n1217), .A2(G378), .A3(new_n1242), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1218), .B(new_n1241), .C1(new_n1213), .C2(new_n1006), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1266), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1271), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1263), .A2(KEYINPUT60), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1155), .A2(new_n1095), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1263), .A2(KEYINPUT60), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1283), .B2(new_n1261), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G384), .B(new_n1261), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1277), .A2(new_n1278), .A3(new_n1287), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1283), .A2(new_n1261), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n888), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1271), .A2(G2897), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1285), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1292), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1289), .B1(new_n1277), .B2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1278), .B1(new_n1277), .B2(new_n1287), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1288), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(G393), .B(new_n849), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1127), .B1(new_n1034), .B2(new_n1059), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1300), .B1(new_n1267), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G387), .A2(G390), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1034), .A2(new_n1059), .A3(new_n1127), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1300), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  OR2_X1    g1108(.A1(new_n1277), .A2(new_n1296), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT61), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1309), .A2(new_n1302), .A3(new_n1306), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1277), .A2(new_n1287), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1277), .A2(KEYINPUT63), .A3(new_n1287), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  OAI22_X1  g1116(.A1(new_n1299), .A2(new_n1308), .B1(new_n1311), .B2(new_n1316), .ZN(G405));
  NAND2_X1  g1117(.A1(G375), .A2(new_n1266), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1274), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1287), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1318), .B(new_n1274), .C1(new_n1284), .C2(new_n1286), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1307), .B(new_n1322), .ZN(G402));
endmodule


