//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n207), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n210), .B1(new_n214), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n234), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  AND2_X1   g0049(.A1(new_n249), .A2(new_n211), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(G20), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n250), .A2(G68), .A3(new_n252), .A4(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n254), .B(KEYINPUT72), .Z(new_n255));
  NAND2_X1  g0055(.A1(new_n249), .A2(new_n211), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G50), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n258), .A2(new_n259), .B1(new_n212), .B2(G68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n212), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n223), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n256), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT11), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n263), .A2(new_n264), .ZN(new_n266));
  INV_X1    g0066(.A(new_n252), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n217), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT12), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n255), .A2(new_n265), .A3(new_n266), .A4(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G169), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  OAI211_X1 g0073(.A(G1), .B(G13), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n272), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G226), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT70), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT70), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n278), .A2(new_n283), .A3(G226), .A4(new_n279), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n276), .A2(new_n277), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n236), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n287), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n274), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  AOI21_X1  g0090(.A(G1), .B1(new_n273), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G274), .ZN(new_n292));
  INV_X1    g0092(.A(new_n291), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n274), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(KEYINPUT71), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT71), .ZN(new_n297));
  OAI21_X1  g0097(.A(G238), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n292), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OR3_X1    g0099(.A1(new_n289), .A2(new_n299), .A3(KEYINPUT13), .ZN(new_n300));
  OAI21_X1  g0100(.A(KEYINPUT13), .B1(new_n289), .B2(new_n299), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n271), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT14), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(new_n301), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n302), .A2(new_n303), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n270), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(G200), .ZN(new_n310));
  INV_X1    g0110(.A(new_n270), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n300), .A2(G190), .A3(new_n301), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(G58), .A2(G68), .ZN(new_n315));
  OAI211_X1 g0115(.A(KEYINPUT73), .B(G20), .C1(new_n315), .C2(new_n201), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n257), .A2(G159), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(G58), .B(G68), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT73), .B1(new_n319), .B2(G20), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT74), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(G20), .B1(new_n315), .B2(new_n201), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT73), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT74), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(new_n316), .A4(new_n317), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n276), .A2(new_n212), .A3(new_n277), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT7), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT7), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n276), .A2(new_n329), .A3(new_n212), .A4(new_n277), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(G68), .A3(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n321), .A2(KEYINPUT16), .A3(new_n326), .A4(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT16), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n328), .A2(G68), .A3(new_n330), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n324), .A2(new_n316), .A3(new_n317), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(new_n336), .A3(new_n256), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT8), .ZN(new_n338));
  INV_X1    g0138(.A(G58), .ZN(new_n339));
  OR3_X1    g0139(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT67), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n338), .B1(new_n339), .B2(KEYINPUT67), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n267), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n250), .A2(new_n253), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(new_n342), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n337), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT75), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n281), .A2(G1698), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n278), .B(new_n349), .C1(G223), .C2(G1698), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G87), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n274), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n292), .B1(new_n294), .B2(new_n236), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n271), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n352), .A2(new_n354), .A3(new_n307), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT75), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n337), .A2(new_n360), .A3(new_n346), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n348), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT76), .B(KEYINPUT18), .Z(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT77), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n331), .A2(new_n324), .A3(new_n316), .A4(new_n317), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n250), .B1(new_n367), .B2(new_n333), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n345), .B1(new_n368), .B2(new_n332), .ZN(new_n369));
  INV_X1    g0169(.A(G190), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n353), .A2(new_n370), .A3(new_n355), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n352), .B2(new_n354), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT17), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  AND4_X1   g0175(.A1(KEYINPUT17), .A2(new_n374), .A3(new_n337), .A4(new_n346), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n366), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(new_n337), .A3(new_n346), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT17), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n369), .A2(KEYINPUT17), .A3(new_n374), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT77), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n348), .A2(new_n359), .A3(new_n361), .A4(new_n363), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n365), .A2(new_n377), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n292), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n295), .B2(G226), .ZN(new_n387));
  AND2_X1   g0187(.A1(KEYINPUT66), .A2(G223), .ZN(new_n388));
  NOR2_X1   g0188(.A1(KEYINPUT66), .A2(G223), .ZN(new_n389));
  OAI21_X1  g0189(.A(G1698), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(G222), .A2(G1698), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n286), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n274), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(new_n278), .B2(G77), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n387), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G190), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n342), .A2(new_n261), .ZN(new_n398));
  OAI21_X1  g0198(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n399));
  INV_X1    g0199(.A(G150), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(new_n258), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n256), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  MUX2_X1   g0202(.A(new_n252), .B(new_n344), .S(G50), .Z(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT9), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n402), .A2(KEYINPUT9), .A3(new_n403), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n397), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT10), .B1(new_n408), .B2(KEYINPUT69), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n372), .B2(new_n396), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n408), .B1(KEYINPUT69), .B2(KEYINPUT10), .C1(new_n372), .C2(new_n396), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n395), .A2(new_n271), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n413), .B(new_n404), .C1(G179), .C2(new_n395), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT15), .B(G87), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT68), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n417), .A2(new_n261), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT8), .B(G58), .Z(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n250), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n267), .A2(new_n223), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n344), .B2(new_n223), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n278), .A2(G1698), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n425), .A2(new_n218), .B1(new_n225), .B2(new_n278), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n279), .B2(new_n287), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n292), .B1(new_n224), .B2(new_n294), .C1(new_n427), .C2(new_n274), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n271), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G179), .B2(new_n428), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(G200), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(new_n424), .C1(new_n370), .C2(new_n428), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n415), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n314), .A2(new_n385), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n286), .A2(G303), .ZN(new_n437));
  INV_X1    g0237(.A(G257), .ZN(new_n438));
  OAI221_X1 g0238(.A(new_n437), .B1(new_n280), .B2(new_n438), .C1(new_n226), .C2(new_n425), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n393), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n251), .B(G45), .C1(new_n273), .C2(KEYINPUT5), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT80), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT5), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(G41), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(G270), .A3(new_n274), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n274), .B(G274), .C1(new_n443), .C2(G41), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT80), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n441), .B(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT81), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n442), .A2(KEYINPUT81), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n440), .A2(new_n445), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT20), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n455), .B(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G97), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n212), .B1(new_n458), .B2(G33), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n256), .B1(new_n212), .B2(G116), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n454), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n461), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(KEYINPUT20), .C1(new_n457), .C2(new_n459), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n250), .B(new_n252), .C1(G1), .C2(new_n272), .ZN(new_n466));
  MUX2_X1   g0266(.A(new_n252), .B(new_n466), .S(G116), .Z(new_n467));
  AOI21_X1  g0267(.A(new_n271), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n453), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT21), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n453), .A2(G200), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n465), .A2(new_n467), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n472), .B(new_n473), .C1(new_n370), .C2(new_n453), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n453), .A2(new_n468), .A3(KEYINPUT21), .ZN(new_n475));
  OR3_X1    g0275(.A1(new_n453), .A2(new_n473), .A3(new_n307), .ZN(new_n476));
  AND4_X1   g0276(.A1(new_n471), .A2(new_n474), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n278), .A2(new_n212), .A3(G87), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n478), .B(KEYINPUT22), .ZN(new_n479));
  INV_X1    g0279(.A(G116), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n272), .A2(new_n480), .A3(G20), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT23), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n212), .B2(G107), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n225), .A2(KEYINPUT23), .A3(G20), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT24), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n479), .A2(new_n488), .A3(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n256), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n466), .A2(KEYINPUT78), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n466), .A2(KEYINPUT78), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G107), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT25), .ZN(new_n496));
  AOI211_X1 g0296(.A(G107), .B(new_n252), .C1(KEYINPUT84), .C2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(KEYINPUT84), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n497), .B(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g0300(.A(KEYINPUT85), .B(G294), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G33), .ZN(new_n502));
  OAI221_X1 g0302(.A(new_n502), .B1(new_n280), .B2(new_n220), .C1(new_n438), .C2(new_n425), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n393), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n444), .A2(G264), .A3(new_n274), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(G200), .B1(new_n506), .B2(new_n452), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n505), .ZN(new_n508));
  INV_X1    g0308(.A(new_n452), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n508), .A2(new_n509), .A3(G190), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n491), .B(new_n500), .C1(new_n507), .C2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n280), .B2(new_n224), .ZN(new_n513));
  INV_X1    g0313(.A(new_n457), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n280), .A2(new_n512), .A3(new_n224), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n393), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n444), .A2(G257), .A3(new_n274), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n452), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n252), .A2(G97), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n492), .A2(new_n493), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n458), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n225), .A2(KEYINPUT6), .A3(G97), .ZN(new_n526));
  XOR2_X1   g0326(.A(G97), .B(G107), .Z(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(KEYINPUT6), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n328), .A2(G107), .A3(new_n330), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n250), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n521), .B(new_n532), .C1(new_n370), .C2(new_n520), .ZN(new_n533));
  INV_X1    g0333(.A(new_n532), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n520), .A2(new_n271), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n518), .A2(new_n452), .A3(new_n307), .A4(new_n519), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n511), .A2(new_n533), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n506), .A2(new_n307), .A3(new_n452), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n271), .B1(new_n508), .B2(new_n509), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n250), .B1(new_n487), .B2(new_n489), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n495), .A2(new_n499), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n278), .A2(G238), .A3(new_n279), .ZN(new_n544));
  OAI221_X1 g0344(.A(new_n544), .B1(new_n272), .B2(new_n480), .C1(new_n425), .C2(new_n224), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n393), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n290), .A2(G1), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(new_n220), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n274), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT82), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT82), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n551), .A3(new_n274), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n550), .A2(new_n552), .B1(G274), .B2(new_n547), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(G179), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n271), .ZN(new_n557));
  INV_X1    g0357(.A(new_n417), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n492), .A2(new_n558), .A3(new_n493), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n278), .A2(new_n212), .A3(G68), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n261), .A2(new_n458), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n560), .B1(KEYINPUT19), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n212), .A2(new_n563), .B1(new_n204), .B2(new_n219), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n256), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n417), .A2(new_n267), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n559), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n567), .A2(KEYINPUT83), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT83), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n565), .A2(new_n566), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(new_n570), .B2(new_n559), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n556), .B(new_n557), .C1(new_n568), .C2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n565), .B(new_n566), .C1(new_n524), .C2(new_n219), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n372), .B1(new_n546), .B2(new_n553), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n554), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G190), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n543), .A2(new_n572), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n538), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n436), .A2(new_n477), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n581), .B(KEYINPUT86), .ZN(G372));
  INV_X1    g0382(.A(new_n573), .ZN(new_n583));
  INV_X1    g0383(.A(new_n574), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(KEYINPUT87), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT87), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n573), .B2(new_n574), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n587), .A3(new_n577), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n572), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n538), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n543), .A2(new_n471), .A3(new_n475), .A4(new_n476), .ZN(new_n591));
  OR2_X1    g0391(.A1(new_n568), .A2(new_n571), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n555), .B1(new_n271), .B2(new_n554), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n590), .A2(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n595), .A2(KEYINPUT26), .A3(new_n572), .A4(new_n578), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT88), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n572), .A2(new_n578), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT88), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(new_n595), .A4(KEYINPUT26), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT26), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n589), .B2(new_n537), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n597), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n436), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n309), .A2(new_n430), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n313), .A2(new_n377), .A3(new_n382), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n369), .A2(new_n358), .ZN(new_n609));
  XNOR2_X1  g0409(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n610), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n369), .B2(new_n358), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n412), .B(new_n411), .C1(new_n608), .C2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n605), .A2(new_n414), .A3(new_n615), .ZN(G369));
  AND2_X1   g0416(.A1(new_n476), .A2(new_n475), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n471), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n251), .A2(new_n212), .A3(G13), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(G213), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(G343), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n473), .A2(new_n625), .ZN(new_n626));
  MUX2_X1   g0426(.A(new_n477), .B(new_n618), .S(new_n626), .Z(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G330), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n543), .A2(new_n624), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n624), .B1(new_n541), .B2(new_n542), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n511), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n631), .A2(new_n543), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n628), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n633), .B(KEYINPUT90), .ZN(new_n634));
  INV_X1    g0434(.A(new_n629), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n632), .A2(new_n629), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n618), .A2(new_n625), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n634), .A2(new_n635), .A3(new_n639), .ZN(G399));
  INV_X1    g0440(.A(new_n208), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(G41), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G1), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n215), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT28), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n624), .B1(new_n594), .B2(new_n603), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT29), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n511), .A2(new_n537), .A3(new_n533), .ZN(new_n651));
  INV_X1    g0451(.A(new_n589), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(new_n591), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n572), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT26), .B1(new_n589), .B2(new_n537), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n598), .A2(new_n601), .A3(new_n595), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n625), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT29), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n650), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT95), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n543), .A2(new_n578), .A3(new_n572), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n651), .A2(new_n477), .A3(new_n662), .A4(new_n625), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT94), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n520), .A2(new_n453), .A3(new_n307), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n504), .A2(new_n505), .A3(new_n546), .A4(new_n553), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT91), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT91), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT30), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n554), .B(KEYINPUT92), .ZN(new_n672));
  AOI21_X1  g0472(.A(G179), .B1(new_n506), .B2(new_n452), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(new_n453), .A4(new_n520), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n665), .A2(new_n667), .A3(KEYINPUT30), .A4(new_n668), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n624), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT31), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT94), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n580), .A2(new_n680), .A3(new_n477), .A4(new_n625), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n664), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n676), .A2(KEYINPUT31), .A3(new_n624), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT93), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT93), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n676), .A2(new_n685), .A3(KEYINPUT31), .A4(new_n624), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(G330), .B1(new_n682), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n660), .A2(new_n661), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n650), .A2(new_n659), .ZN(new_n690));
  INV_X1    g0490(.A(G330), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n664), .A2(new_n679), .A3(new_n681), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n684), .A2(new_n686), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT95), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n647), .B1(new_n696), .B2(G1), .ZN(G364));
  NOR2_X1   g0497(.A1(new_n627), .A2(G330), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT96), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT96), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n212), .A2(G13), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n251), .B1(new_n701), .B2(G45), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OR3_X1    g0503(.A1(new_n703), .A2(new_n642), .A3(KEYINPUT97), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT97), .B1(new_n703), .B2(new_n642), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n699), .A2(new_n628), .A3(new_n700), .A4(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n211), .B1(G20), .B2(new_n271), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  XOR2_X1   g0509(.A(KEYINPUT33), .B(G317), .Z(new_n710));
  NOR2_X1   g0510(.A1(new_n307), .A2(new_n372), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n212), .A2(G190), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n212), .A2(new_n370), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n372), .A2(G179), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G303), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n286), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G179), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n714), .B(new_n719), .C1(G329), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n715), .A2(new_n711), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(KEYINPUT99), .B(G326), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n212), .B1(new_n720), .B2(G190), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n725), .A2(new_n727), .B1(new_n729), .B2(new_n501), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT100), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n307), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n715), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G322), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n712), .A2(new_n716), .ZN(new_n737));
  INV_X1    g0537(.A(G283), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n734), .A2(new_n712), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n739), .B1(G311), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n723), .A2(new_n732), .A3(new_n733), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n717), .A2(new_n219), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n278), .B1(new_n735), .B2(new_n339), .ZN(new_n745));
  INV_X1    g0545(.A(new_n713), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n744), .B(new_n745), .C1(G68), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n729), .A2(G97), .ZN(new_n748));
  INV_X1    g0548(.A(G159), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n721), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT32), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n724), .A2(new_n259), .B1(new_n740), .B2(new_n223), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n737), .A2(new_n225), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n747), .A2(new_n748), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n709), .B1(new_n743), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n708), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n278), .A2(new_n208), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT98), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n762), .A2(G355), .B1(new_n480), .B2(new_n641), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n247), .A2(G45), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n641), .A2(new_n278), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G45), .B2(new_n215), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n763), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n706), .B(new_n756), .C1(new_n760), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n759), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n627), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n707), .A2(new_n770), .ZN(G396));
  INV_X1    g0571(.A(new_n706), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n430), .A2(new_n624), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n432), .B1(new_n424), .B2(new_n625), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n430), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n648), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n648), .A2(new_n778), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n772), .B1(new_n781), .B2(new_n688), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n694), .A2(new_n779), .A3(new_n780), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n778), .A2(new_n758), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G137), .A2(new_n725), .B1(new_n746), .B2(G150), .ZN(new_n786));
  INV_X1    g0586(.A(new_n735), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G143), .A2(new_n787), .B1(new_n741), .B2(G159), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT34), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(KEYINPUT34), .ZN(new_n791));
  INV_X1    g0591(.A(G132), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n278), .B1(new_n721), .B2(new_n792), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n717), .A2(new_n259), .B1(new_n737), .B2(new_n217), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n793), .B(new_n794), .C1(G58), .C2(new_n729), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n790), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n724), .A2(new_n718), .B1(new_n717), .B2(new_n225), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n278), .B(new_n797), .C1(G294), .C2(new_n787), .ZN(new_n798));
  INV_X1    g0598(.A(new_n737), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G87), .A2(new_n799), .B1(new_n722), .B2(G311), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n746), .A2(G283), .B1(new_n741), .B2(G116), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n798), .A2(new_n748), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n709), .B1(new_n796), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n708), .A2(new_n757), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n706), .B1(new_n223), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n785), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n784), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G384));
  AOI211_X1 g0609(.A(new_n480), .B(new_n214), .C1(new_n528), .C2(KEYINPUT35), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(KEYINPUT35), .B2(new_n528), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT36), .Z(new_n812));
  OR3_X1    g0612(.A1(new_n215), .A2(new_n223), .A3(new_n315), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n259), .A2(G68), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n251), .B(G13), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n664), .A2(new_n679), .A3(new_n681), .A4(new_n683), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n311), .A2(new_n625), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n309), .A2(new_n313), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n305), .A2(new_n308), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n821), .B2(new_n819), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n817), .A2(new_n778), .A3(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT40), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n321), .A2(new_n326), .A3(new_n331), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n333), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n332), .A2(new_n256), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n346), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n622), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n384), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT103), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n348), .A2(new_n361), .A3(new_n830), .ZN(new_n834));
  XOR2_X1   g0634(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n835));
  AND2_X1   g0635(.A1(new_n378), .A2(new_n835), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n362), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n829), .A2(new_n830), .B1(new_n369), .B2(new_n374), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n829), .A2(new_n359), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n833), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n362), .A2(new_n834), .A3(new_n836), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n839), .A2(new_n840), .ZN(new_n844));
  OAI211_X1 g0644(.A(KEYINPUT103), .B(new_n843), .C1(new_n844), .C2(new_n838), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n832), .A2(new_n842), .A3(new_n845), .A4(KEYINPUT38), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n609), .B1(new_n369), .B2(new_n374), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n835), .B1(new_n847), .B2(new_n834), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n380), .A2(new_n381), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n614), .A2(new_n849), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n837), .A2(new_n848), .B1(new_n850), .B2(new_n834), .ZN(new_n851));
  XNOR2_X1  g0651(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n824), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n823), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT108), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT108), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n823), .A2(new_n857), .A3(new_n854), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n832), .A2(new_n842), .A3(new_n845), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT104), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n862), .A2(new_n863), .A3(new_n846), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n860), .A2(KEYINPUT104), .A3(new_n861), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n823), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n824), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n436), .A2(new_n817), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n691), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n774), .B1(new_n648), .B2(new_n778), .ZN(new_n873));
  INV_X1    g0673(.A(new_n822), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n875), .A2(new_n866), .B1(new_n614), .B2(new_n622), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT39), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n846), .A2(new_n853), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT107), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n864), .A2(KEYINPUT39), .A3(new_n865), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT105), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n864), .A2(KEYINPUT105), .A3(KEYINPUT39), .A4(new_n865), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n821), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(new_n270), .A3(new_n625), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n876), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n435), .B1(new_n650), .B2(new_n659), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n615), .A2(new_n414), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n887), .A2(new_n890), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n872), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n251), .B2(new_n701), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n872), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n816), .B1(new_n894), .B2(new_n895), .ZN(G367));
  NOR2_X1   g0696(.A1(new_n583), .A2(new_n625), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n589), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n592), .A2(new_n593), .A3(new_n897), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n759), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n233), .A2(new_n765), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n760), .C1(new_n208), .C2(new_n417), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n772), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(KEYINPUT112), .B(G317), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n740), .A2(new_n738), .B1(new_n721), .B2(new_n904), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n278), .B(new_n905), .C1(G303), .C2(new_n787), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n225), .B2(new_n728), .ZN(new_n907));
  INV_X1    g0707(.A(new_n717), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(G116), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT46), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n725), .A2(G311), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n799), .A2(G97), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n746), .A2(new_n501), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(G143), .A2(new_n725), .B1(new_n908), .B2(G58), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n729), .A2(G68), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n286), .B1(new_n787), .B2(G150), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(KEYINPUT113), .B(G137), .Z(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n722), .A2(new_n920), .B1(new_n799), .B2(G77), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n921), .B1(new_n259), .B2(new_n740), .C1(new_n749), .C2(new_n713), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n907), .A2(new_n914), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT47), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n903), .B1(new_n924), .B2(new_n708), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n900), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT111), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT110), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n637), .B1(new_n632), .B2(new_n629), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n639), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(G330), .A3(new_n627), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n628), .A2(new_n639), .A3(new_n929), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n928), .B1(new_n696), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n933), .ZN(new_n935));
  AOI211_X1 g0735(.A(KEYINPUT110), .B(new_n935), .C1(new_n689), .C2(new_n695), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n537), .B(new_n533), .C1(new_n532), .C2(new_n625), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n595), .A2(new_n624), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n639), .A2(new_n635), .A3(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT45), .Z(new_n942));
  AOI21_X1  g0742(.A(new_n940), .B1(new_n639), .B2(new_n635), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT44), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n942), .A2(new_n634), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n634), .B1(new_n942), .B2(new_n944), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n927), .B1(new_n937), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n689), .A2(new_n695), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT110), .B1(new_n949), .B2(new_n935), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n696), .A2(new_n928), .A3(new_n933), .ZN(new_n951));
  AND4_X1   g0751(.A1(new_n927), .A2(new_n950), .A3(new_n951), .A4(new_n947), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n696), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n642), .B(KEYINPUT41), .Z(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n703), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n636), .A2(new_n638), .A3(new_n940), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(KEYINPUT42), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(KEYINPUT42), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n537), .B1(new_n938), .B2(new_n543), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n625), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n898), .A2(new_n899), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(new_n962), .C2(new_n964), .ZN(new_n969));
  INV_X1    g0769(.A(new_n940), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n634), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n969), .B(new_n971), .Z(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n926), .B1(new_n956), .B2(new_n973), .ZN(G387));
  OAI21_X1  g0774(.A(new_n286), .B1(new_n737), .B2(new_n480), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n724), .A2(new_n736), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n735), .A2(new_n904), .B1(new_n740), .B2(new_n718), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(G311), .C2(new_n746), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT48), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(KEYINPUT48), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n908), .A2(new_n501), .B1(new_n729), .B2(G283), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n982), .B(new_n983), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n975), .B(new_n984), .C1(new_n722), .C2(new_n727), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n417), .A2(new_n728), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n724), .A2(new_n749), .B1(new_n735), .B2(new_n259), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G77), .B2(new_n908), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n342), .A2(new_n713), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G68), .A2(new_n741), .B1(new_n722), .B2(G150), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(new_n278), .A3(new_n912), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n708), .B1(new_n985), .B2(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n239), .A2(new_n290), .ZN(new_n996));
  INV_X1    g0796(.A(new_n644), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n996), .A2(new_n765), .B1(new_n997), .B2(new_n762), .ZN(new_n998));
  INV_X1    g0798(.A(new_n419), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n999), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n644), .B(new_n290), .C1(new_n217), .C2(new_n223), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n419), .B2(new_n259), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n998), .A2(new_n1004), .B1(G107), .B2(new_n208), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n706), .B1(new_n1005), .B2(new_n760), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n995), .B(new_n1006), .C1(new_n636), .C2(new_n769), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n933), .A2(new_n703), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT114), .Z(new_n1009));
  OAI21_X1  g0809(.A(new_n642), .B1(new_n696), .B2(new_n933), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1007), .B(new_n1009), .C1(new_n937), .C2(new_n1010), .ZN(G393));
  NAND2_X1  g0811(.A1(new_n947), .A2(KEYINPUT116), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT116), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n945), .B2(new_n946), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n703), .A3(new_n1014), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n244), .A2(new_n641), .A3(new_n278), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n760), .B1(new_n458), .B2(new_n208), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n772), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(G317), .A2(new_n725), .B1(new_n787), .B2(G311), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT52), .Z(new_n1020));
  AOI22_X1  g0820(.A1(new_n746), .A2(G303), .B1(new_n741), .B2(G294), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G283), .A2(new_n908), .B1(new_n722), .B2(G322), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n278), .B(new_n753), .C1(G116), .C2(new_n729), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G68), .A2(new_n908), .B1(new_n722), .B2(G143), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1025), .B(new_n278), .C1(new_n219), .C2(new_n737), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT118), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n728), .A2(new_n223), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n999), .A2(new_n740), .B1(new_n259), .B2(new_n713), .ZN(new_n1029));
  OR3_X1    g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n724), .A2(new_n400), .B1(new_n735), .B2(new_n749), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT117), .Z(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT51), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1024), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1018), .B1(new_n1034), .B2(new_n708), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n940), .B2(new_n769), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1015), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n950), .A2(new_n951), .A3(new_n947), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT111), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n937), .A2(new_n927), .A3(new_n947), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n937), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n947), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n643), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1037), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(G390));
  AND2_X1   g0846(.A1(new_n884), .A2(new_n757), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n706), .B1(new_n342), .B2(new_n804), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G132), .A2(new_n787), .B1(new_n799), .B2(G50), .ZN(new_n1049));
  INV_X1    g0849(.A(G125), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n721), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT53), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n717), .B2(new_n400), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n908), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(KEYINPUT54), .B(G143), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n278), .B1(new_n740), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(G128), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n713), .A2(new_n919), .B1(new_n724), .B2(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(G159), .C2(new_n729), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n713), .A2(new_n225), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n724), .A2(new_n738), .B1(new_n735), .B2(new_n480), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(G294), .C2(new_n722), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n217), .A2(new_n737), .B1(new_n740), .B2(new_n458), .ZN(new_n1064));
  NOR4_X1   g0864(.A1(new_n1064), .A2(new_n744), .A3(new_n1028), .A4(new_n278), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1055), .A2(new_n1060), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1048), .B1(new_n1066), .B2(new_n709), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1047), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n694), .A2(new_n778), .A3(new_n822), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n773), .B1(new_n658), .B2(new_n777), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n822), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n886), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n846), .B2(new_n853), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n886), .B1(new_n873), .B2(new_n874), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1070), .B(new_n1076), .C1(new_n884), .C2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n817), .A2(new_n822), .A3(G330), .A4(new_n778), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n882), .A2(new_n883), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n879), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n1081), .A3(new_n1077), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1079), .B1(new_n1082), .B2(new_n1075), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1078), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1068), .B1(new_n1084), .B2(new_n703), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT120), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n870), .A2(new_n691), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1087), .A2(new_n888), .A3(new_n889), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1071), .ZN(new_n1089));
  OAI211_X1 g0889(.A(G330), .B(new_n778), .C1(new_n682), .C2(new_n687), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n874), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n817), .A2(G330), .A3(new_n778), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n874), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1090), .A2(new_n874), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n873), .B1(new_n1096), .B2(new_n1079), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1088), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT119), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n643), .B1(new_n1084), .B2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(KEYINPUT119), .B(new_n1098), .C1(new_n1078), .C2(new_n1083), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1086), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1082), .A2(new_n1069), .A3(new_n1075), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1076), .B1(new_n884), .B2(new_n1077), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1099), .B(new_n1103), .C1(new_n1104), .C2(new_n1079), .ZN(new_n1105));
  AND4_X1   g0905(.A1(new_n1086), .A2(new_n1101), .A3(new_n1105), .A4(new_n642), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1085), .B1(new_n1102), .B2(new_n1106), .ZN(G378));
  NAND2_X1  g0907(.A1(new_n404), .A2(new_n830), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n415), .B(new_n1108), .Z(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1109), .B(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n887), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1111), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n876), .C1(new_n884), .C2(new_n886), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n869), .A2(new_n691), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1112), .A2(new_n1116), .A3(new_n1114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1111), .A2(new_n757), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G116), .A2(new_n725), .B1(new_n746), .B2(G97), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1122), .B(new_n916), .C1(new_n225), .C2(new_n735), .ZN(new_n1123));
  AOI211_X1 g0923(.A(G41), .B(new_n278), .C1(new_n908), .C2(G77), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1124), .B1(new_n339), .B2(new_n737), .C1(new_n738), .C2(new_n721), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT121), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1123), .B(new_n1126), .C1(new_n558), .C2(new_n741), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(KEYINPUT58), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n724), .A2(new_n1050), .B1(new_n713), .B2(new_n792), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n741), .A2(G137), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n1058), .B2(new_n735), .C1(new_n717), .C2(new_n1056), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1129), .B(new_n1131), .C1(G150), .C2(new_n729), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT59), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n799), .A2(G159), .ZN(new_n1136));
  AOI211_X1 g0936(.A(G33), .B(G41), .C1(new_n722), .C2(G124), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1128), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1127), .A2(KEYINPUT58), .B1(G50), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n708), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT122), .Z(new_n1143));
  AOI211_X1 g0943(.A(new_n706), .B(new_n1143), .C1(new_n259), .C2(new_n804), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1120), .A2(new_n703), .B1(new_n1121), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1069), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1096), .A2(new_n1079), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n873), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1103), .B(new_n1148), .C1(new_n1104), .C2(new_n1079), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1088), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1112), .A2(new_n1116), .A3(new_n1114), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1116), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1150), .B(KEYINPUT57), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n642), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT57), .B1(new_n1120), .B2(new_n1150), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1145), .B1(new_n1154), .B2(new_n1155), .ZN(G375));
  NAND2_X1  g0956(.A1(new_n874), .A2(new_n757), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT123), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n706), .B1(new_n217), .B2(new_n804), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G294), .A2(new_n725), .B1(new_n746), .B2(G116), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n458), .B2(new_n717), .C1(new_n225), .C2(new_n740), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G283), .A2(new_n787), .B1(new_n722), .B2(G303), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1162), .B(new_n286), .C1(new_n223), .C2(new_n737), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1161), .A2(new_n1163), .A3(new_n986), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n717), .A2(new_n749), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n713), .A2(new_n1056), .B1(new_n721), .B2(new_n1058), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(G150), .C2(new_n741), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n787), .A2(new_n920), .B1(new_n725), .B2(G132), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n286), .B1(new_n799), .B2(G58), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n259), .C2(new_n728), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1164), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1158), .B(new_n1159), .C1(new_n709), .C2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1148), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n702), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1148), .A2(new_n1088), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n955), .A3(new_n1098), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1176), .A2(new_n1178), .ZN(G381));
  OAI21_X1  g0979(.A(new_n703), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1144), .A2(new_n1121), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1118), .A2(new_n1119), .B1(new_n1088), .B2(new_n1149), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n643), .B1(new_n1183), .B2(KEYINPUT57), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1182), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1101), .A2(new_n1105), .A3(new_n642), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1085), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1045), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT124), .ZN(new_n1195));
  OR4_X1    g0995(.A1(G387), .A2(new_n1192), .A3(new_n1193), .A4(new_n1195), .ZN(G407));
  OAI211_X1 g0996(.A(G407), .B(G213), .C1(G343), .C2(new_n1192), .ZN(G409));
  XOR2_X1   g0997(.A(G393), .B(G396), .Z(new_n1198));
  NAND2_X1  g0998(.A1(G387), .A2(new_n1045), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n949), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n702), .B1(new_n1200), .B2(new_n954), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n972), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1202), .A2(new_n926), .A3(G390), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1198), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1199), .A2(new_n1198), .A3(new_n1203), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1088), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n642), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1148), .A2(new_n1088), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(KEYINPUT60), .B2(new_n1098), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1176), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n808), .ZN(new_n1214));
  OAI211_X1 g1014(.A(G384), .B(new_n1176), .C1(new_n1210), .C2(new_n1212), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n623), .A2(G213), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(G2897), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1216), .B(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1183), .A2(new_n955), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1190), .B1(new_n1145), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n1188), .B2(G378), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1220), .B1(new_n1223), .B2(new_n1218), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT61), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1185), .A2(new_n954), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1191), .B1(new_n1226), .B2(new_n1182), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1085), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1189), .A2(KEYINPUT120), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1100), .A2(new_n1086), .A3(new_n1101), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1227), .B1(G375), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT62), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1216), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1217), .A4(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1224), .A2(new_n1225), .A3(new_n1235), .ZN(new_n1236));
  XOR2_X1   g1036(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1237));
  NAND3_X1  g1037(.A1(new_n1187), .A2(new_n642), .A3(new_n1153), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(G378), .A3(new_n1145), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1218), .B1(new_n1239), .B2(new_n1227), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1237), .B1(new_n1240), .B2(new_n1234), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1207), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G390), .B1(new_n1202), .B2(new_n926), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n926), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1244), .B(new_n1045), .C1(new_n1201), .C2(new_n972), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1198), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1243), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(new_n1204), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT63), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1232), .A2(new_n1217), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1216), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT61), .B1(new_n1250), .B2(new_n1220), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1240), .A2(KEYINPUT63), .A3(new_n1234), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1248), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1242), .A2(new_n1254), .ZN(G405));
  NAND2_X1  g1055(.A1(G375), .A2(new_n1191), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT126), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1256), .A2(new_n1257), .A3(new_n1239), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1257), .B1(new_n1256), .B2(new_n1239), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1234), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G375), .A2(new_n1231), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1190), .B1(new_n1238), .B2(new_n1145), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT126), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1256), .A2(new_n1239), .A3(new_n1257), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1216), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1207), .B1(new_n1260), .B2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1234), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1263), .A2(new_n1216), .A3(new_n1264), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n1248), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(G402));
endmodule


