//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G146), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT0), .A3(G128), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT0), .B(G128), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G125), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT1), .B1(new_n187), .B2(G146), .ZN(new_n196));
  OAI211_X1 g010(.A(G128), .B(new_n196), .C1(new_n188), .C2(new_n190), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n189), .A2(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n187), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n198), .B(new_n199), .C1(KEYINPUT1), .C2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n195), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G953), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G224), .ZN(new_n207));
  XOR2_X1   g021(.A(new_n207), .B(KEYINPUT78), .Z(new_n208));
  XNOR2_X1  g022(.A(new_n205), .B(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n211), .A2(KEYINPUT3), .A3(G104), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT3), .B1(new_n211), .B2(G104), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT73), .B1(new_n211), .B2(G104), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT73), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n217), .A3(G107), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT74), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n217), .B2(G107), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n211), .A2(KEYINPUT3), .A3(G104), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT74), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n225), .A2(new_n226), .A3(new_n215), .A4(new_n218), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n220), .A2(new_n221), .A3(G101), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT2), .A2(G113), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n229), .B(KEYINPUT66), .ZN(new_n230));
  OR2_X1    g044(.A1(KEYINPUT2), .A2(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G116), .B(G119), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n228), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n220), .A2(G101), .A3(new_n227), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT75), .ZN(new_n240));
  INV_X1    g054(.A(G101), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n225), .A2(new_n241), .A3(new_n215), .A4(new_n218), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n242), .A2(KEYINPUT4), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n239), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n240), .B1(new_n239), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n238), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n217), .A2(G107), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n211), .A2(G104), .ZN(new_n248));
  OAI21_X1  g062(.A(G101), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT76), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT76), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n242), .A2(new_n252), .A3(new_n249), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n233), .A2(KEYINPUT5), .ZN(new_n255));
  INV_X1    g069(.A(G119), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G116), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n255), .B(G113), .C1(KEYINPUT5), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n254), .A2(new_n236), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G122), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n246), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n246), .A2(new_n259), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n260), .B(KEYINPUT77), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n261), .A2(KEYINPUT6), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n265));
  INV_X1    g079(.A(new_n263), .ZN(new_n266));
  AOI211_X1 g080(.A(new_n265), .B(new_n266), .C1(new_n246), .C2(new_n259), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n210), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n258), .A2(new_n236), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n250), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n259), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n260), .B(KEYINPUT8), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT79), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n194), .B2(G125), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n207), .A2(KEYINPUT7), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n205), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n195), .A2(new_n273), .A3(new_n204), .A4(new_n275), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n271), .A2(new_n272), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(G902), .B1(new_n279), .B2(new_n261), .ZN(new_n280));
  OAI21_X1  g094(.A(G210), .B1(G237), .B2(G902), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n268), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT81), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n268), .A2(KEYINPUT81), .A3(new_n280), .A4(new_n281), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n281), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n261), .A2(KEYINPUT6), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n262), .A2(new_n263), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n267), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n209), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n280), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT80), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n281), .B1(new_n268), .B2(new_n280), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT80), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n286), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G475), .A2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT84), .ZN(new_n302));
  OR2_X1    g116(.A1(KEYINPUT67), .A2(G953), .ZN(new_n303));
  INV_X1    g117(.A(G237), .ZN(new_n304));
  NAND2_X1  g118(.A1(KEYINPUT67), .A2(G953), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n303), .A2(G214), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n187), .ZN(new_n307));
  AND2_X1   g121(.A1(KEYINPUT67), .A2(G953), .ZN(new_n308));
  NOR2_X1   g122(.A1(KEYINPUT67), .A2(G953), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n310), .A2(G143), .A3(G214), .A4(new_n304), .ZN(new_n311));
  NAND2_X1  g125(.A1(KEYINPUT18), .A2(G131), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n307), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT82), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n307), .A2(new_n311), .A3(KEYINPUT82), .A4(new_n312), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n312), .B1(new_n307), .B2(new_n311), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(G146), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n307), .A2(new_n311), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT64), .B(G131), .Z(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT64), .B(G131), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n307), .A2(new_n311), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n203), .A2(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT83), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT19), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n319), .A2(KEYINPUT83), .A3(KEYINPUT19), .ZN(new_n334));
  AOI21_X1  g148(.A(G146), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT71), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n329), .B2(KEYINPUT16), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT16), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT16), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n339), .A2(new_n328), .A3(KEYINPUT71), .A4(G125), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n337), .A2(new_n338), .A3(G146), .A4(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n317), .A2(new_n321), .B1(new_n327), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G113), .B(G122), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(new_n217), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n302), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n346), .ZN(new_n348));
  AOI211_X1 g162(.A(new_n318), .B(new_n320), .C1(new_n315), .C2(new_n316), .ZN(new_n349));
  AOI211_X1 g163(.A(new_n335), .B(new_n342), .C1(new_n324), .C2(new_n326), .ZN(new_n350));
  OAI211_X1 g164(.A(KEYINPUT84), .B(new_n348), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n322), .A2(KEYINPUT17), .A3(new_n323), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n189), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n341), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT17), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n324), .A2(new_n358), .A3(new_n326), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n324), .A2(KEYINPUT85), .A3(new_n358), .A4(new_n326), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n357), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n349), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n346), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n301), .B1(new_n352), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT20), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT86), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT86), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n356), .B1(new_n360), .B2(new_n359), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n349), .B1(new_n370), .B2(new_n362), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n346), .A2(new_n371), .B1(new_n347), .B2(new_n351), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n369), .B(KEYINPUT20), .C1(new_n372), .C2(new_n301), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n352), .A2(new_n365), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n367), .A3(new_n300), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n368), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n348), .A2(KEYINPUT87), .ZN(new_n377));
  AOI21_X1  g191(.A(G902), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n378), .B1(new_n371), .B2(new_n377), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G475), .ZN(new_n380));
  INV_X1    g194(.A(G902), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n200), .A2(G143), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT89), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n187), .A2(G128), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT13), .ZN(new_n387));
  INV_X1    g201(.A(G134), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G116), .B(G122), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT88), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n391), .A2(G107), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n384), .A2(new_n385), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n384), .A2(new_n387), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(G134), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(G107), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n389), .A2(new_n392), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G122), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G116), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n211), .B1(new_n399), .B2(KEYINPUT14), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n390), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n386), .A2(new_n388), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n393), .A2(G134), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT9), .B(G234), .ZN(new_n405));
  INV_X1    g219(.A(G217), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n405), .A2(new_n406), .A3(G953), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n397), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n397), .B2(new_n404), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n381), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT15), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G478), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(G952), .ZN(new_n415));
  AOI211_X1 g229(.A(G953), .B(new_n415), .C1(G234), .C2(G237), .ZN(new_n416));
  AOI211_X1 g230(.A(new_n381), .B(new_n310), .C1(G234), .C2(G237), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT21), .B(G898), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n410), .A2(new_n412), .A3(G478), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n414), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n376), .A2(new_n380), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G469), .ZN(new_n424));
  INV_X1    g238(.A(new_n194), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n228), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n426), .B1(new_n244), .B2(new_n245), .ZN(new_n427));
  INV_X1    g241(.A(G137), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT11), .A3(G134), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n388), .A2(G137), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT65), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT11), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n388), .B2(G137), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n431), .A2(new_n432), .A3(new_n325), .A4(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n429), .A3(new_n430), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT65), .B1(new_n436), .B2(new_n323), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n435), .A2(new_n437), .B1(G131), .B2(new_n436), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT10), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n202), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n202), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n242), .A3(new_n249), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n254), .A2(new_n440), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n427), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n310), .A2(G227), .ZN(new_n445));
  XOR2_X1   g259(.A(G110), .B(G140), .Z(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n251), .A2(new_n202), .A3(new_n253), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n442), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n435), .A2(new_n437), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n436), .A2(G131), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT12), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT12), .ZN(new_n456));
  AOI211_X1 g270(.A(new_n456), .B(new_n438), .C1(new_n450), .C2(new_n442), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n449), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n228), .A2(new_n425), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n239), .A2(new_n243), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT75), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n239), .A2(new_n240), .A3(new_n243), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n242), .A2(new_n252), .A3(new_n249), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n252), .B1(new_n242), .B2(new_n249), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n440), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n442), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n467), .B1(new_n468), .B2(KEYINPUT10), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n454), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n448), .B1(new_n470), .B2(new_n444), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n424), .B(new_n381), .C1(new_n459), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(G469), .A2(G902), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n470), .A2(new_n444), .A3(new_n448), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n464), .A2(new_n469), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n465), .A2(new_n466), .A3(new_n441), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n454), .B1(new_n476), .B2(new_n468), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n456), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n451), .A2(KEYINPUT12), .A3(new_n454), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n475), .A2(new_n438), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(G469), .B(new_n474), .C1(new_n480), .C2(new_n448), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n472), .A2(new_n473), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G221), .B1(new_n405), .B2(G902), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n423), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G214), .B1(G237), .B2(G902), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n299), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n388), .A2(G137), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n428), .A2(G134), .ZN(new_n489));
  OAI21_X1  g303(.A(G131), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n197), .A2(new_n201), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n435), .B2(new_n437), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n492), .B1(new_n454), .B2(new_n425), .ZN(new_n493));
  INV_X1    g307(.A(new_n237), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n194), .B1(new_n452), .B2(new_n453), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n496), .A2(new_n237), .A3(new_n492), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT28), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT26), .B(G101), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n310), .A2(G210), .A3(new_n304), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT27), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n501), .A2(KEYINPUT27), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n502), .A3(new_n499), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n497), .A2(KEYINPUT28), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n498), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n496), .B2(new_n492), .ZN(new_n514));
  INV_X1    g328(.A(new_n491), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n452), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n516), .B(KEYINPUT30), .C1(new_n438), .C2(new_n194), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n237), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n497), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n508), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n511), .A2(new_n512), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n381), .B1(new_n511), .B2(new_n512), .ZN(new_n523));
  OAI21_X1  g337(.A(G472), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(G472), .A2(G902), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT31), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n508), .B1(new_n493), .B2(new_n494), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n518), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT69), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n518), .A2(new_n528), .A3(KEYINPUT69), .A4(new_n527), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n498), .A2(new_n510), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n508), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n518), .A2(new_n528), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT68), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT68), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n518), .A2(new_n537), .A3(new_n528), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(KEYINPUT31), .A3(new_n538), .ZN(new_n539));
  AOI211_X1 g353(.A(KEYINPUT32), .B(new_n526), .C1(new_n534), .C2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n531), .A2(new_n532), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n533), .A2(new_n508), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n541), .B1(new_n544), .B2(new_n525), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n524), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n256), .A2(G128), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT23), .B1(new_n200), .B2(G119), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n548), .A2(KEYINPUT23), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n549), .A2(new_n550), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT72), .B(G110), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G119), .B(G128), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT24), .B(G110), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n554), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n319), .A2(new_n189), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n341), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n355), .A2(new_n341), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n555), .ZN(new_n562));
  INV_X1    g376(.A(G110), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(new_n552), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n310), .A2(G221), .A3(G234), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT22), .B(G137), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n560), .A2(new_n564), .A3(new_n568), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n381), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT25), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n406), .B1(G234), .B2(new_n381), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n571), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n575), .A2(G902), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n574), .A2(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n546), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n487), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(new_n241), .ZN(G3));
  AOI21_X1  g396(.A(new_n526), .B1(new_n534), .B2(new_n539), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n544), .A2(new_n381), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(G472), .ZN(new_n585));
  INV_X1    g399(.A(new_n483), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n481), .A2(new_n473), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(new_n472), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT90), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n585), .A2(new_n588), .A3(new_n589), .A4(new_n579), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n482), .A2(new_n483), .A3(new_n579), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n544), .A2(new_n525), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n534), .B2(new_n539), .ZN(new_n593));
  INV_X1    g407(.A(G472), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT90), .B1(new_n591), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n292), .A2(new_n293), .A3(new_n287), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n486), .B1(new_n598), .B2(new_n297), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT91), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT92), .B1(new_n408), .B2(new_n409), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT33), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(KEYINPUT92), .B(KEYINPUT33), .C1(new_n408), .C2(new_n409), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G478), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(G902), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n605), .A2(new_n607), .B1(new_n606), .B2(new_n410), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n419), .B(new_n608), .C1(new_n376), .C2(new_n380), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n294), .A2(new_n282), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT91), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n486), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n600), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n597), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NAND2_X1  g430(.A1(new_n375), .A2(KEYINPUT93), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n366), .A2(new_n618), .A3(new_n367), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n617), .A2(new_n368), .A3(new_n373), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n410), .B(new_n413), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(G475), .B2(new_n379), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n620), .A2(new_n420), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n600), .A2(new_n623), .A3(new_n612), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n597), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT35), .B(G107), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NAND2_X1  g441(.A1(new_n574), .A2(new_n575), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n569), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n565), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n578), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n595), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n299), .A2(new_n485), .A3(new_n633), .A4(new_n486), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT37), .B(G110), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  AOI21_X1  g450(.A(new_n611), .B1(new_n610), .B2(new_n486), .ZN(new_n637));
  INV_X1    g451(.A(new_n486), .ZN(new_n638));
  AOI211_X1 g452(.A(KEYINPUT91), .B(new_n638), .C1(new_n294), .C2(new_n282), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n592), .A2(KEYINPUT32), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n583), .A2(new_n541), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n632), .B1(new_n643), .B2(new_n524), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT94), .B(G900), .Z(new_n645));
  NAND2_X1  g459(.A1(new_n417), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n416), .B1(new_n647), .B2(KEYINPUT95), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(KEYINPUT95), .B2(new_n647), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n620), .A2(new_n622), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n640), .A2(new_n644), .A3(new_n588), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  NAND2_X1  g466(.A1(new_n536), .A2(new_n538), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n495), .A2(new_n497), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n653), .B1(new_n508), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(G472), .B1(new_n655), .B2(G902), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n643), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n649), .B(KEYINPUT39), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n588), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n657), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n621), .B1(new_n376), .B2(new_n380), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n299), .B(KEYINPUT38), .Z(new_n664));
  OAI211_X1 g478(.A(new_n486), .B(new_n632), .C1(new_n660), .C2(new_n658), .ZN(new_n665));
  OR3_X1    g479(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  NAND2_X1  g481(.A1(new_n376), .A2(new_n380), .ZN(new_n668));
  INV_X1    g482(.A(new_n608), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n649), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n640), .A2(new_n644), .A3(new_n588), .A4(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT96), .B(G146), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G48));
  NOR2_X1   g488(.A1(new_n459), .A2(new_n471), .ZN(new_n675));
  OAI21_X1  g489(.A(G469), .B1(new_n675), .B2(G902), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n472), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n586), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n546), .A2(new_n678), .A3(new_n579), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n613), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT41), .B(G113), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT97), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n680), .B(new_n682), .ZN(G15));
  NOR2_X1   g497(.A1(new_n624), .A2(new_n679), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(G116), .Z(G18));
  NAND3_X1  g499(.A1(new_n600), .A2(new_n612), .A3(new_n678), .ZN(new_n686));
  INV_X1    g500(.A(new_n668), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n628), .A2(new_n631), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n546), .A2(new_n687), .A3(new_n422), .A4(new_n688), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  XOR2_X1   g505(.A(new_n525), .B(KEYINPUT98), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n544), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n693), .B(new_n579), .C1(new_n593), .C2(new_n594), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n676), .A2(new_n420), .A3(new_n483), .A4(new_n472), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n696), .A2(new_n600), .A3(new_n612), .A4(new_n662), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G122), .ZN(G24));
  OAI211_X1 g512(.A(new_n688), .B(new_n693), .C1(new_n593), .C2(new_n594), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n670), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n640), .A2(new_n700), .A3(new_n678), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT99), .B(G125), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G27));
  AND4_X1   g517(.A1(new_n486), .A2(new_n286), .A3(new_n296), .A4(new_n298), .ZN(new_n704));
  INV_X1    g518(.A(new_n579), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n643), .B2(new_n524), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT100), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n587), .A2(new_n707), .A3(new_n472), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n482), .A2(KEYINPUT100), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n708), .A2(new_n709), .A3(new_n483), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n704), .A2(new_n706), .A3(new_n671), .A4(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n286), .A2(new_n486), .A3(new_n296), .A4(new_n298), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n708), .A2(new_n709), .A3(new_n483), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(KEYINPUT42), .A3(new_n706), .A4(new_n671), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G131), .ZN(G33));
  NAND4_X1  g533(.A1(new_n704), .A2(new_n706), .A3(new_n650), .A4(new_n710), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT101), .B(G134), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G36));
  NAND2_X1  g536(.A1(new_n687), .A2(new_n669), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(KEYINPUT43), .Z(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(KEYINPUT103), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(KEYINPUT103), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n595), .A3(new_n688), .A4(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n474), .B1(new_n480), .B2(new_n448), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n424), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n732), .B2(new_n731), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n734), .A2(new_n473), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT102), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(KEYINPUT46), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n736), .A2(new_n472), .A3(new_n737), .ZN(new_n738));
  OR3_X1    g552(.A1(new_n735), .A2(KEYINPUT102), .A3(KEYINPUT46), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n586), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n659), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n714), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n729), .A2(new_n730), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G137), .ZN(G39));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(KEYINPUT104), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(KEYINPUT104), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n740), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n740), .A2(new_n748), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n670), .A2(new_n546), .A3(new_n579), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n704), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  OR2_X1    g569(.A1(new_n677), .A2(KEYINPUT49), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n677), .A2(KEYINPUT49), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n705), .A2(new_n638), .A3(new_n586), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n657), .A2(new_n756), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n664), .A2(new_n759), .A3(new_n687), .A4(new_n669), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n724), .A2(new_n416), .ZN(new_n761));
  INV_X1    g575(.A(new_n694), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n638), .A3(new_n664), .A4(new_n678), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(KEYINPUT50), .Z(new_n766));
  NAND3_X1  g580(.A1(new_n657), .A2(new_n416), .A3(new_n579), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n714), .A2(new_n586), .A3(new_n677), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(new_n687), .A3(new_n608), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n761), .A2(new_n769), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n766), .B(new_n770), .C1(new_n699), .C2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n752), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n676), .A2(new_n586), .A3(new_n472), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT112), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(KEYINPUT112), .A3(new_n776), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n704), .A3(new_n764), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n774), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n714), .B(new_n763), .C1(new_n775), .C2(new_n776), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n773), .B1(new_n772), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n771), .A2(new_n580), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT48), .Z(new_n784));
  NAND4_X1  g598(.A1(new_n768), .A2(new_n668), .A3(new_n669), .A4(new_n769), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n785), .A2(G952), .A3(new_n206), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n784), .B(new_n786), .C1(new_n686), .C2(new_n763), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT113), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n780), .A2(new_n782), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n704), .A2(new_n700), .A3(new_n710), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n380), .A2(new_n621), .A3(new_n649), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n588), .A2(new_n620), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n704), .A2(new_n644), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n720), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n679), .B1(new_n613), .B2(new_n624), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n697), .B1(new_n686), .B2(new_n689), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n621), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n376), .A2(new_n798), .A3(new_n380), .A4(new_n420), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n299), .A2(new_n486), .A3(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n634), .B(KEYINPUT105), .C1(new_n597), .C2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n299), .A2(new_n609), .A3(new_n486), .ZN(new_n802));
  OAI22_X1  g616(.A1(new_n597), .A2(new_n802), .B1(new_n487), .B2(new_n580), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT105), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n634), .B1(new_n597), .B2(new_n800), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n797), .A2(new_n718), .A3(new_n801), .A4(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT106), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT107), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n632), .A2(new_n649), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n643), .B2(new_n656), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n640), .A2(new_n811), .A3(new_n662), .A4(new_n710), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n651), .A2(new_n672), .A3(new_n812), .A4(new_n701), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(KEYINPUT52), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(KEYINPUT52), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n809), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n651), .A2(new_n701), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n818), .A3(new_n672), .A4(new_n812), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n813), .A2(KEYINPUT52), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT107), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n808), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT108), .B1(new_n824), .B2(KEYINPUT53), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT108), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n720), .A2(new_n790), .A3(new_n793), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n796), .A2(new_n795), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n718), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n805), .A2(new_n804), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n597), .A2(new_n802), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n581), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n832), .A2(new_n834), .A3(new_n801), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n831), .A2(new_n819), .A3(new_n820), .A4(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n825), .B(new_n828), .C1(new_n827), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT54), .ZN(new_n838));
  INV_X1    g652(.A(new_n679), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n839), .B(new_n640), .C1(new_n609), .C2(new_n623), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n690), .A3(KEYINPUT110), .A4(new_n697), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n796), .B2(new_n795), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n843), .A3(new_n718), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT111), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n841), .A2(new_n843), .A3(new_n718), .A4(KEYINPUT111), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n835), .A2(KEYINPUT53), .A3(new_n829), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n822), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT109), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n819), .A2(new_n820), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n852), .B(new_n827), .C1(new_n807), .C2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n852), .B1(new_n836), .B2(new_n827), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n850), .B(new_n851), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n838), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n789), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n415), .A2(new_n206), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT114), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n760), .B1(new_n859), .B2(new_n861), .ZN(G75));
  NOR2_X1   g676(.A1(new_n264), .A2(new_n267), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n209), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n268), .ZN(new_n865));
  XNOR2_X1  g679(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n865), .B(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n850), .B1(new_n855), .B2(new_n856), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(G902), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n869), .A2(G210), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n867), .B1(new_n870), .B2(KEYINPUT56), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT116), .Z(new_n872));
  NOR2_X1   g686(.A1(new_n310), .A2(G952), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n867), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n874), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n872), .A2(new_n877), .ZN(G51));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n868), .A2(KEYINPUT54), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n881), .A3(new_n857), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n868), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n473), .B(KEYINPUT57), .Z(new_n884));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n882), .A2(new_n887), .A3(new_n883), .A4(new_n884), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n879), .B1(new_n889), .B2(new_n675), .ZN(new_n890));
  INV_X1    g704(.A(new_n869), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n734), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n675), .B1(new_n886), .B2(new_n888), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n893), .B2(KEYINPUT120), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n873), .B1(new_n890), .B2(new_n894), .ZN(G54));
  AND3_X1   g709(.A1(new_n869), .A2(KEYINPUT58), .A3(G475), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n874), .B1(new_n896), .B2(new_n374), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n374), .B2(new_n896), .ZN(G60));
  NAND2_X1  g712(.A1(G478), .A2(G902), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT59), .Z(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n605), .B1(new_n858), .B2(new_n901), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n605), .A2(new_n882), .A3(new_n883), .A4(new_n901), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n873), .A3(new_n903), .ZN(G63));
  OAI21_X1  g718(.A(new_n874), .B1(KEYINPUT122), .B2(KEYINPUT61), .ZN(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n406), .A2(new_n381), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n906), .B(new_n907), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n868), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n909), .B2(new_n630), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n577), .B2(new_n909), .ZN(new_n911));
  NAND2_X1  g725(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(G66));
  INV_X1    g727(.A(G224), .ZN(new_n914));
  OAI21_X1  g728(.A(G953), .B1(new_n418), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n835), .A2(new_n830), .ZN(new_n916));
  INV_X1    g730(.A(new_n310), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n863), .B1(G898), .B2(new_n310), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(G69));
  NAND3_X1  g734(.A1(new_n754), .A2(new_n718), .A3(new_n720), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n817), .A2(new_n672), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT124), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n743), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n640), .A2(new_n706), .A3(new_n662), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n741), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT127), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n921), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n310), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n514), .A2(new_n517), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n333), .A2(new_n334), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT123), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n930), .B(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n917), .A2(G900), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n929), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n668), .A2(new_n669), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n668), .B2(new_n621), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n704), .A2(new_n706), .A3(new_n937), .A4(new_n660), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n743), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT126), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n923), .A2(new_n666), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n754), .B1(KEYINPUT62), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(KEYINPUT62), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT125), .Z(new_n945));
  AOI21_X1  g759(.A(new_n917), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n935), .B1(new_n946), .B2(new_n933), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n310), .B1(G227), .B2(G900), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n948), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n935), .B(new_n950), .C1(new_n946), .C2(new_n933), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(G72));
  NAND2_X1  g766(.A1(new_n520), .A2(new_n509), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n943), .A2(new_n916), .A3(new_n945), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT63), .Z(new_n956));
  AOI21_X1  g770(.A(new_n953), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n536), .A2(new_n521), .A3(new_n538), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n837), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n956), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n928), .B2(new_n916), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n518), .A2(new_n519), .A3(new_n508), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n874), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n957), .A2(new_n959), .A3(new_n963), .ZN(G57));
endmodule


