

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593;

  XNOR2_X1 U324 ( .A(KEYINPUT117), .B(KEYINPUT47), .ZN(n411) );
  XNOR2_X1 U325 ( .A(n329), .B(n328), .ZN(n334) );
  XNOR2_X1 U326 ( .A(n412), .B(n411), .ZN(n421) );
  XOR2_X1 U327 ( .A(n372), .B(n371), .Z(n292) );
  XNOR2_X1 U328 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U329 ( .A(n327), .B(KEYINPUT11), .ZN(n328) );
  XNOR2_X1 U330 ( .A(n383), .B(n382), .ZN(n385) );
  INV_X1 U331 ( .A(KEYINPUT106), .ZN(n414) );
  INV_X1 U332 ( .A(n337), .ZN(n338) );
  XNOR2_X1 U333 ( .A(n414), .B(KEYINPUT36), .ZN(n415) );
  XNOR2_X1 U334 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U335 ( .A(n564), .B(n415), .ZN(n590) );
  XNOR2_X1 U336 ( .A(n341), .B(n340), .ZN(n346) );
  NOR2_X1 U337 ( .A1(n462), .A2(n531), .ZN(n572) );
  XNOR2_X1 U338 ( .A(n463), .B(G190GAT), .ZN(n464) );
  XNOR2_X1 U339 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n294) );
  XNOR2_X1 U341 ( .A(KEYINPUT90), .B(KEYINPUT23), .ZN(n293) );
  XNOR2_X1 U342 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U343 ( .A(n295), .B(KEYINPUT22), .Z(n297) );
  XOR2_X1 U344 ( .A(G22GAT), .B(G155GAT), .Z(n349) );
  XNOR2_X1 U345 ( .A(n349), .B(KEYINPUT89), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n297), .B(n296), .ZN(n303) );
  XOR2_X1 U347 ( .A(G211GAT), .B(KEYINPUT21), .Z(n299) );
  XNOR2_X1 U348 ( .A(G197GAT), .B(G218GAT), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n317) );
  XOR2_X1 U350 ( .A(G50GAT), .B(G162GAT), .Z(n336) );
  XOR2_X1 U351 ( .A(n317), .B(n336), .Z(n301) );
  NAND2_X1 U352 ( .A1(G228GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U354 ( .A(n303), .B(n302), .Z(n311) );
  XOR2_X1 U355 ( .A(KEYINPUT88), .B(KEYINPUT2), .Z(n305) );
  XNOR2_X1 U356 ( .A(KEYINPUT3), .B(KEYINPUT87), .ZN(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U358 ( .A(G141GAT), .B(n306), .Z(n430) );
  XOR2_X1 U359 ( .A(G148GAT), .B(G106GAT), .Z(n308) );
  XNOR2_X1 U360 ( .A(G204GAT), .B(G78GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U362 ( .A(KEYINPUT73), .B(n309), .Z(n377) );
  XNOR2_X1 U363 ( .A(n430), .B(n377), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n473) );
  XOR2_X1 U365 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n313) );
  XNOR2_X1 U366 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U368 ( .A(n314), .B(KEYINPUT18), .Z(n316) );
  XNOR2_X1 U369 ( .A(G169GAT), .B(G183GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n461) );
  XOR2_X1 U371 ( .A(G36GAT), .B(KEYINPUT79), .Z(n337) );
  XOR2_X1 U372 ( .A(n337), .B(n317), .Z(n319) );
  NAND2_X1 U373 ( .A1(G226GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U375 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n321) );
  XNOR2_X1 U376 ( .A(G176GAT), .B(G204GAT), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U378 ( .A(n323), .B(n322), .Z(n325) );
  XOR2_X1 U379 ( .A(G8GAT), .B(KEYINPUT80), .Z(n350) );
  XOR2_X1 U380 ( .A(G92GAT), .B(G64GAT), .Z(n379) );
  XNOR2_X1 U381 ( .A(n350), .B(n379), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n461), .B(n326), .ZN(n528) );
  XOR2_X1 U384 ( .A(G43GAT), .B(G134GAT), .Z(n457) );
  XOR2_X1 U385 ( .A(G85GAT), .B(KEYINPUT74), .Z(n378) );
  XNOR2_X1 U386 ( .A(n457), .B(n378), .ZN(n329) );
  XOR2_X1 U387 ( .A(KEYINPUT10), .B(KEYINPUT66), .Z(n327) );
  XOR2_X1 U388 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n331) );
  XNOR2_X1 U389 ( .A(G190GAT), .B(KEYINPUT78), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U391 ( .A(G218GAT), .B(n332), .Z(n333) );
  XNOR2_X1 U392 ( .A(n334), .B(n333), .ZN(n341) );
  XNOR2_X1 U393 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n335), .B(KEYINPUT7), .ZN(n394) );
  XNOR2_X1 U395 ( .A(n394), .B(n336), .ZN(n339) );
  XOR2_X1 U396 ( .A(G92GAT), .B(G106GAT), .Z(n343) );
  NAND2_X1 U397 ( .A1(G232GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U399 ( .A(G99GAT), .B(n344), .Z(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n564) );
  XOR2_X1 U401 ( .A(KEYINPUT81), .B(G64GAT), .Z(n348) );
  XNOR2_X1 U402 ( .A(G78GAT), .B(G211GAT), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n364) );
  XOR2_X1 U404 ( .A(n350), .B(n349), .Z(n352) );
  XNOR2_X1 U405 ( .A(G71GAT), .B(G183GAT), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n357) );
  XOR2_X1 U407 ( .A(G15GAT), .B(G127GAT), .Z(n451) );
  XNOR2_X1 U408 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n353), .B(KEYINPUT13), .ZN(n373) );
  XOR2_X1 U410 ( .A(n451), .B(n373), .Z(n355) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U413 ( .A(n357), .B(n356), .Z(n362) );
  XOR2_X1 U414 ( .A(KEYINPUT70), .B(G1GAT), .Z(n391) );
  XOR2_X1 U415 ( .A(KEYINPUT82), .B(KEYINPUT14), .Z(n359) );
  XNOR2_X1 U416 ( .A(KEYINPUT15), .B(KEYINPUT12), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n391), .B(n360), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U420 ( .A(n364), .B(n363), .Z(n497) );
  INV_X1 U421 ( .A(n497), .ZN(n587) );
  INV_X1 U422 ( .A(G120GAT), .ZN(n365) );
  NAND2_X1 U423 ( .A1(n365), .A2(G71GAT), .ZN(n368) );
  INV_X1 U424 ( .A(G71GAT), .ZN(n366) );
  NAND2_X1 U425 ( .A1(n366), .A2(G120GAT), .ZN(n367) );
  NAND2_X1 U426 ( .A1(n368), .A2(n367), .ZN(n370) );
  XNOR2_X1 U427 ( .A(G99GAT), .B(G176GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n456) );
  XOR2_X1 U429 ( .A(n456), .B(KEYINPUT31), .Z(n372) );
  NAND2_X1 U430 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n292), .B(n373), .ZN(n383) );
  XOR2_X1 U432 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n375) );
  XNOR2_X1 U433 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  INV_X1 U437 ( .A(n385), .ZN(n413) );
  INV_X1 U438 ( .A(KEYINPUT41), .ZN(n384) );
  NAND2_X1 U439 ( .A1(n413), .A2(n384), .ZN(n387) );
  NAND2_X1 U440 ( .A1(n385), .A2(KEYINPUT41), .ZN(n386) );
  NAND2_X1 U441 ( .A1(n387), .A2(n386), .ZN(n512) );
  XOR2_X1 U442 ( .A(G15GAT), .B(G113GAT), .Z(n389) );
  XNOR2_X1 U443 ( .A(G36GAT), .B(G50GAT), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U445 ( .A(n390), .B(G43GAT), .Z(n393) );
  XNOR2_X1 U446 ( .A(G169GAT), .B(n391), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n398) );
  XOR2_X1 U448 ( .A(n394), .B(KEYINPUT69), .Z(n396) );
  NAND2_X1 U449 ( .A1(G229GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U451 ( .A(n398), .B(n397), .Z(n406) );
  XOR2_X1 U452 ( .A(G8GAT), .B(G197GAT), .Z(n400) );
  XNOR2_X1 U453 ( .A(G141GAT), .B(G22GAT), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U455 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n402) );
  XNOR2_X1 U456 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n406), .B(n405), .ZN(n579) );
  NAND2_X1 U460 ( .A1(n512), .A2(n579), .ZN(n407) );
  XOR2_X1 U461 ( .A(KEYINPUT46), .B(n407), .Z(n408) );
  NOR2_X1 U462 ( .A1(n587), .A2(n408), .ZN(n409) );
  XOR2_X1 U463 ( .A(KEYINPUT116), .B(n409), .Z(n410) );
  NOR2_X1 U464 ( .A1(n564), .A2(n410), .ZN(n412) );
  INV_X1 U465 ( .A(n413), .ZN(n582) );
  XNOR2_X1 U466 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n417) );
  NOR2_X1 U467 ( .A1(n497), .A2(n590), .ZN(n416) );
  XOR2_X1 U468 ( .A(n417), .B(n416), .Z(n418) );
  NAND2_X1 U469 ( .A1(n582), .A2(n418), .ZN(n419) );
  NOR2_X1 U470 ( .A1(n579), .A2(n419), .ZN(n420) );
  NOR2_X1 U471 ( .A1(n421), .A2(n420), .ZN(n422) );
  XNOR2_X1 U472 ( .A(n422), .B(KEYINPUT48), .ZN(n538) );
  NOR2_X1 U473 ( .A1(n528), .A2(n538), .ZN(n423) );
  XNOR2_X1 U474 ( .A(n423), .B(KEYINPUT54), .ZN(n448) );
  XOR2_X1 U475 ( .A(KEYINPUT96), .B(KEYINPUT94), .Z(n425) );
  XNOR2_X1 U476 ( .A(KEYINPUT92), .B(KEYINPUT95), .ZN(n424) );
  XNOR2_X1 U477 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U478 ( .A(KEYINPUT4), .B(n426), .Z(n428) );
  NAND2_X1 U479 ( .A1(G225GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U481 ( .A(n429), .B(KEYINPUT1), .Z(n432) );
  XNOR2_X1 U482 ( .A(n430), .B(KEYINPUT93), .ZN(n431) );
  XNOR2_X1 U483 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U484 ( .A(G155GAT), .B(G148GAT), .Z(n434) );
  XNOR2_X1 U485 ( .A(G1GAT), .B(G127GAT), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U487 ( .A(n436), .B(n435), .Z(n447) );
  XOR2_X1 U488 ( .A(KEYINPUT78), .B(G85GAT), .Z(n438) );
  XNOR2_X1 U489 ( .A(G134GAT), .B(G162GAT), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U491 ( .A(G113GAT), .B(KEYINPUT0), .Z(n454) );
  XOR2_X1 U492 ( .A(n439), .B(n454), .Z(n441) );
  XNOR2_X1 U493 ( .A(G29GAT), .B(G120GAT), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U495 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n443) );
  XNOR2_X1 U496 ( .A(G57GAT), .B(KEYINPUT91), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U499 ( .A(n447), .B(n446), .Z(n553) );
  INV_X1 U500 ( .A(n553), .ZN(n525) );
  NAND2_X1 U501 ( .A1(n448), .A2(n525), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n449), .B(KEYINPUT64), .ZN(n578) );
  NOR2_X1 U503 ( .A1(n473), .A2(n578), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n450), .B(KEYINPUT55), .ZN(n462) );
  XOR2_X1 U505 ( .A(KEYINPUT20), .B(n451), .Z(n453) );
  NAND2_X1 U506 ( .A1(G227GAT), .A2(G233GAT), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n455) );
  XOR2_X1 U508 ( .A(n455), .B(n454), .Z(n459) );
  XNOR2_X1 U509 ( .A(n456), .B(n457), .ZN(n458) );
  XNOR2_X1 U510 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U511 ( .A(n461), .B(n460), .Z(n540) );
  INV_X1 U512 ( .A(n540), .ZN(n531) );
  NAND2_X1 U513 ( .A1(n572), .A2(n564), .ZN(n465) );
  XOR2_X1 U514 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n463) );
  XOR2_X1 U515 ( .A(n473), .B(KEYINPUT28), .Z(n534) );
  XOR2_X1 U516 ( .A(KEYINPUT27), .B(n528), .Z(n470) );
  NAND2_X1 U517 ( .A1(n534), .A2(n470), .ZN(n466) );
  NOR2_X1 U518 ( .A1(n525), .A2(n466), .ZN(n539) );
  XNOR2_X1 U519 ( .A(KEYINPUT85), .B(n540), .ZN(n467) );
  NAND2_X1 U520 ( .A1(n539), .A2(n467), .ZN(n480) );
  XOR2_X1 U521 ( .A(KEYINPUT99), .B(KEYINPUT26), .Z(n469) );
  NAND2_X1 U522 ( .A1(n473), .A2(n531), .ZN(n468) );
  XNOR2_X1 U523 ( .A(n469), .B(n468), .ZN(n577) );
  INV_X1 U524 ( .A(n470), .ZN(n471) );
  NOR2_X1 U525 ( .A1(n577), .A2(n471), .ZN(n554) );
  XOR2_X1 U526 ( .A(n554), .B(KEYINPUT100), .Z(n477) );
  NOR2_X1 U527 ( .A1(n531), .A2(n528), .ZN(n472) );
  NOR2_X1 U528 ( .A1(n473), .A2(n472), .ZN(n475) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U531 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U532 ( .A1(n525), .A2(n478), .ZN(n479) );
  NAND2_X1 U533 ( .A1(n480), .A2(n479), .ZN(n496) );
  NOR2_X1 U534 ( .A1(n564), .A2(n497), .ZN(n481) );
  XNOR2_X1 U535 ( .A(n481), .B(KEYINPUT16), .ZN(n482) );
  XOR2_X1 U536 ( .A(KEYINPUT83), .B(n482), .Z(n483) );
  AND2_X1 U537 ( .A1(n496), .A2(n483), .ZN(n513) );
  NAND2_X1 U538 ( .A1(n582), .A2(n579), .ZN(n484) );
  XOR2_X1 U539 ( .A(KEYINPUT76), .B(n484), .Z(n501) );
  NAND2_X1 U540 ( .A1(n513), .A2(n501), .ZN(n493) );
  NOR2_X1 U541 ( .A1(n525), .A2(n493), .ZN(n486) );
  XNOR2_X1 U542 ( .A(KEYINPUT34), .B(KEYINPUT102), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U544 ( .A(G1GAT), .B(n487), .Z(G1324GAT) );
  NOR2_X1 U545 ( .A1(n528), .A2(n493), .ZN(n489) );
  XNOR2_X1 U546 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(G1325GAT) );
  NOR2_X1 U548 ( .A1(n531), .A2(n493), .ZN(n491) );
  XNOR2_X1 U549 ( .A(KEYINPUT35), .B(KEYINPUT104), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G15GAT), .B(n492), .ZN(G1326GAT) );
  NOR2_X1 U552 ( .A1(n534), .A2(n493), .ZN(n495) );
  XNOR2_X1 U553 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(G1327GAT) );
  NAND2_X1 U555 ( .A1(n497), .A2(n496), .ZN(n498) );
  NOR2_X1 U556 ( .A1(n590), .A2(n498), .ZN(n500) );
  XNOR2_X1 U557 ( .A(KEYINPUT107), .B(KEYINPUT37), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n500), .B(n499), .ZN(n524) );
  NAND2_X1 U559 ( .A1(n524), .A2(n501), .ZN(n502) );
  XNOR2_X1 U560 ( .A(n502), .B(KEYINPUT38), .ZN(n509) );
  NOR2_X1 U561 ( .A1(n509), .A2(n525), .ZN(n503) );
  XNOR2_X1 U562 ( .A(n503), .B(KEYINPUT39), .ZN(n504) );
  XNOR2_X1 U563 ( .A(G29GAT), .B(n504), .ZN(G1328GAT) );
  NOR2_X1 U564 ( .A1(n509), .A2(n528), .ZN(n505) );
  XOR2_X1 U565 ( .A(KEYINPUT108), .B(n505), .Z(n506) );
  XNOR2_X1 U566 ( .A(G36GAT), .B(n506), .ZN(G1329GAT) );
  NOR2_X1 U567 ( .A1(n509), .A2(n531), .ZN(n507) );
  XOR2_X1 U568 ( .A(KEYINPUT40), .B(n507), .Z(n508) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  XNOR2_X1 U570 ( .A(G50GAT), .B(KEYINPUT109), .ZN(n511) );
  NOR2_X1 U571 ( .A1(n534), .A2(n509), .ZN(n510) );
  XNOR2_X1 U572 ( .A(n511), .B(n510), .ZN(G1331GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT110), .B(n512), .Z(n543) );
  NOR2_X1 U574 ( .A1(n579), .A2(n543), .ZN(n523) );
  NAND2_X1 U575 ( .A1(n523), .A2(n513), .ZN(n520) );
  NOR2_X1 U576 ( .A1(n525), .A2(n520), .ZN(n514) );
  XOR2_X1 U577 ( .A(G57GAT), .B(n514), .Z(n515) );
  XNOR2_X1 U578 ( .A(KEYINPUT42), .B(n515), .ZN(G1332GAT) );
  NOR2_X1 U579 ( .A1(n528), .A2(n520), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(KEYINPUT111), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1333GAT) );
  NOR2_X1 U582 ( .A1(n531), .A2(n520), .ZN(n518) );
  XOR2_X1 U583 ( .A(KEYINPUT112), .B(n518), .Z(n519) );
  XNOR2_X1 U584 ( .A(G71GAT), .B(n519), .ZN(G1334GAT) );
  NOR2_X1 U585 ( .A1(n534), .A2(n520), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  NAND2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n533) );
  NOR2_X1 U589 ( .A1(n525), .A2(n533), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(KEYINPUT113), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(G1336GAT) );
  NOR2_X1 U592 ( .A1(n528), .A2(n533), .ZN(n529) );
  XOR2_X1 U593 ( .A(KEYINPUT114), .B(n529), .Z(n530) );
  XNOR2_X1 U594 ( .A(G92GAT), .B(n530), .ZN(G1337GAT) );
  NOR2_X1 U595 ( .A1(n531), .A2(n533), .ZN(n532) );
  XOR2_X1 U596 ( .A(G99GAT), .B(n532), .Z(G1338GAT) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X1 U598 ( .A(KEYINPUT44), .B(KEYINPUT115), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n537), .ZN(G1339GAT) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U602 ( .A1(n538), .A2(n541), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n579), .A2(n549), .ZN(n542) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n545) );
  INV_X1 U606 ( .A(n543), .ZN(n568) );
  NAND2_X1 U607 ( .A1(n549), .A2(n568), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n547) );
  NAND2_X1 U610 ( .A1(n549), .A2(n587), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U612 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U614 ( .A1(n549), .A2(n564), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U616 ( .A(G134GAT), .B(n552), .Z(G1343GAT) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U618 ( .A1(n538), .A2(n555), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n579), .A2(n563), .ZN(n556) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n558) );
  NAND2_X1 U623 ( .A1(n563), .A2(n512), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  XOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT121), .Z(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n587), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G162GAT), .B(n566), .ZN(G1347GAT) );
  NAND2_X1 U632 ( .A1(n572), .A2(n579), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n572), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n587), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n575) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U643 ( .A(KEYINPUT59), .B(n576), .Z(n581) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n586) );
  NAND2_X1 U645 ( .A1(n586), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U648 ( .A(n586), .ZN(n589) );
  OR2_X1 U649 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U655 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

