//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT2), .B(G113), .Z(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G116), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n200), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(new_n194), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n206), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(KEYINPUT11), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(G134), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT11), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G137), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n213), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n211), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G134), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G134), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n216), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n212), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n209), .A2(new_n210), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n218), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n230));
  INV_X1    g044(.A(G143), .ZN(new_n231));
  INV_X1    g045(.A(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT64), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G146), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n231), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n232), .A2(G143), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n232), .A2(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n233), .A2(new_n235), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G143), .ZN(new_n242));
  XOR2_X1   g056(.A(KEYINPUT0), .B(G128), .Z(new_n243));
  AOI22_X1  g057(.A1(new_n239), .A2(KEYINPUT0), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n229), .A2(new_n230), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n230), .B1(new_n229), .B2(new_n244), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(new_n223), .B2(G137), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n214), .A2(KEYINPUT68), .A3(new_n206), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n249), .B(new_n250), .C1(G134), .C2(new_n206), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G131), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n241), .B2(G143), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n253), .B(new_n242), .C1(new_n255), .C2(new_n237), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n241), .A2(G143), .ZN(new_n257));
  INV_X1    g071(.A(new_n238), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n254), .A3(G128), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(G128), .B1(new_n236), .B2(new_n254), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n253), .B1(new_n261), .B2(new_n242), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n228), .B(new_n252), .C1(new_n260), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n205), .B1(new_n247), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n229), .A2(new_n244), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n204), .B(KEYINPUT70), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT28), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n267), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n265), .A3(new_n263), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n193), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n226), .B1(new_n225), .B2(new_n227), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n242), .A2(new_n243), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n257), .A2(KEYINPUT0), .A3(G128), .A4(new_n258), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT67), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n229), .A2(new_n230), .A3(new_n244), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n263), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n263), .A2(KEYINPUT30), .A3(new_n265), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n204), .A3(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n287), .A2(new_n271), .A3(new_n193), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n187), .B1(new_n274), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n266), .A2(new_n267), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n271), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n266), .A2(KEYINPUT72), .A3(new_n267), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(KEYINPUT28), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n193), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n295), .A2(KEYINPUT29), .A3(new_n273), .A4(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n289), .A2(new_n290), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G472), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n287), .A2(new_n271), .A3(new_n296), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT31), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n283), .A2(new_n204), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n272), .B1(new_n302), .B2(new_n271), .ZN(new_n303));
  INV_X1    g117(.A(new_n273), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n193), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n287), .A2(new_n306), .A3(new_n271), .A4(new_n296), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n301), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(G472), .A2(G902), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT32), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n308), .A2(KEYINPUT32), .A3(new_n309), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n299), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT16), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT73), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G125), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n319), .A3(G140), .ZN(new_n320));
  NOR2_X1   g134(.A1(G125), .A2(G140), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n315), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT73), .B(G125), .ZN(new_n324));
  NOR2_X1   g138(.A1(KEYINPUT16), .A2(G140), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n232), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n325), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n321), .B1(new_n324), .B2(G140), .ZN(new_n329));
  OAI211_X1 g143(.A(G146), .B(new_n328), .C1(new_n329), .C2(new_n315), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n330), .A3(KEYINPUT74), .ZN(new_n331));
  INV_X1    g145(.A(new_n323), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n332), .A2(new_n333), .A3(G146), .A4(new_n328), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(G119), .B2(new_n237), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n196), .A2(KEYINPUT23), .A3(G128), .ZN(new_n338));
  OAI22_X1  g152(.A1(new_n337), .A2(new_n338), .B1(G119), .B2(new_n237), .ZN(new_n339));
  XNOR2_X1  g153(.A(G119), .B(G128), .ZN(new_n340));
  XOR2_X1   g154(.A(KEYINPUT24), .B(G110), .Z(new_n341));
  AOI22_X1  g155(.A1(new_n339), .A2(G110), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  OAI22_X1  g157(.A1(new_n339), .A2(G110), .B1(new_n340), .B2(new_n341), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n241), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n330), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  INV_X1    g163(.A(G953), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n350), .A2(G221), .A3(G234), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n349), .B(new_n351), .Z(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n343), .A2(new_n347), .A3(new_n352), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n290), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n357));
  INV_X1    g171(.A(G217), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(G234), .B2(new_n290), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT75), .B(KEYINPUT25), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n357), .B(new_n359), .C1(new_n356), .C2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n359), .A2(G902), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n354), .A2(new_n355), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n314), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g179(.A(KEYINPUT9), .B(G234), .Z(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n367), .A2(new_n358), .A3(G953), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT13), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n369), .B1(new_n237), .B2(G143), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT95), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT96), .ZN(new_n373));
  OAI211_X1 g187(.A(KEYINPUT95), .B(new_n369), .C1(new_n237), .C2(G143), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n237), .A2(G143), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n372), .A2(new_n373), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n231), .A2(G128), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n376), .B1(new_n369), .B2(new_n377), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n370), .A2(new_n371), .B1(new_n237), .B2(G143), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n373), .B1(new_n379), .B2(new_n374), .ZN(new_n380));
  OAI21_X1  g194(.A(G134), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n375), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(new_n214), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n198), .A2(G122), .ZN(new_n384));
  INV_X1    g198(.A(G122), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT94), .B1(new_n385), .B2(G116), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT94), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n198), .A3(G122), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  OR2_X1    g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n390), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n383), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n381), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT97), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT97), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n381), .A2(new_n396), .A3(new_n393), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n382), .A2(new_n214), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(new_n383), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n401));
  OAI21_X1  g215(.A(G107), .B1(new_n384), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n400), .B1(new_n389), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n389), .B2(new_n402), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n368), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n381), .A2(new_n396), .A3(new_n393), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n396), .B1(new_n381), .B2(new_n393), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n404), .B(new_n368), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n290), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G478), .ZN(new_n411));
  NOR2_X1   g225(.A1(KEYINPUT98), .A2(KEYINPUT15), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(KEYINPUT98), .A2(KEYINPUT15), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n417));
  INV_X1    g231(.A(new_n368), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n419), .B2(new_n408), .ZN(new_n420));
  INV_X1    g234(.A(new_n415), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT99), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n416), .A2(KEYINPUT99), .A3(new_n422), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G475), .A2(G902), .ZN(new_n428));
  XNOR2_X1  g242(.A(G113), .B(G122), .ZN(new_n429));
  INV_X1    g243(.A(G104), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(KEYINPUT18), .A2(G131), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G237), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n350), .A3(G214), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(G143), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n189), .B(G214), .C1(new_n437), .C2(G143), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n434), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n440), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n433), .B2(new_n432), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n443), .B2(new_n434), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT87), .B1(new_n329), .B2(G146), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n329), .A2(KEYINPUT87), .A3(G146), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n346), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n444), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(KEYINPUT17), .A3(G131), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n439), .A2(new_n440), .A3(new_n226), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT88), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n442), .A2(G131), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n439), .A2(new_n440), .A3(new_n453), .A4(new_n226), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n449), .B1(new_n455), .B2(KEYINPUT17), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n431), .B(new_n448), .C1(new_n335), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(KEYINPUT89), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n320), .A2(KEYINPUT19), .A3(new_n322), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT19), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n345), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n241), .A3(new_n461), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n330), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT89), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n451), .A2(new_n452), .A3(new_n464), .A4(new_n454), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n458), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n431), .B1(new_n466), .B2(new_n448), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n457), .B1(new_n467), .B2(KEYINPUT90), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n469), .B(new_n431), .C1(new_n466), .C2(new_n448), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n428), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT20), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n468), .A2(new_n470), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT20), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n428), .B(KEYINPUT92), .Z(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n475), .A3(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT93), .B(G475), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n448), .B1(new_n335), .B2(new_n456), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(new_n431), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n483), .B1(new_n485), .B2(G902), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n350), .A2(G952), .ZN(new_n488));
  NAND2_X1  g302(.A1(G234), .A2(G237), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g304(.A(KEYINPUT21), .B(G898), .Z(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(G902), .A3(G953), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT100), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n427), .A2(new_n487), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n257), .A2(new_n258), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n240), .A2(KEYINPUT1), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G128), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n254), .A2(new_n239), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n430), .A2(G107), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n390), .A2(G104), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G101), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT78), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT77), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n390), .B2(G104), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n430), .A2(KEYINPUT77), .A3(G107), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G101), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT3), .B1(new_n430), .B2(G107), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT3), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n390), .A3(G104), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n509), .A2(new_n510), .A3(new_n511), .A4(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n503), .A2(new_n515), .A3(G101), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n505), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n500), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT10), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n261), .A2(new_n242), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT69), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n256), .A3(new_n259), .ZN(new_n523));
  INV_X1    g337(.A(new_n517), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(KEYINPUT10), .A3(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n430), .A2(KEYINPUT77), .A3(G107), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT77), .B1(new_n430), .B2(G107), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n511), .B(new_n513), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G101), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(KEYINPUT4), .A3(new_n514), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT4), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n531), .A3(G101), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n244), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n520), .A2(new_n525), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n229), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n520), .A2(new_n525), .A3(new_n277), .A4(new_n533), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n350), .A2(G227), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT76), .ZN(new_n539));
  XNOR2_X1  g353(.A(G110), .B(G140), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n543), .A2(KEYINPUT12), .A3(new_n229), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT12), .B1(new_n543), .B2(new_n229), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n536), .A2(new_n542), .ZN(new_n547));
  OAI22_X1  g361(.A1(new_n537), .A2(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G469), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(new_n290), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT79), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n536), .A2(KEYINPUT79), .A3(new_n542), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n535), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n536), .B1(new_n544), .B2(new_n545), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n541), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n556), .A3(G469), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n549), .A2(new_n290), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n550), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G221), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n366), .B2(new_n290), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G214), .B1(G237), .B2(G902), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n324), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n280), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n523), .B2(new_n567), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT81), .B(G224), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n350), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT7), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n197), .A2(new_n199), .A3(KEYINPUT5), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(G113), .B1(new_n197), .B2(KEYINPUT5), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n574), .A2(new_n576), .B1(new_n202), .B2(new_n194), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n577), .A2(new_n514), .A3(new_n505), .A4(new_n516), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n203), .B1(new_n573), .B2(new_n575), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n517), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(G110), .B(G122), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT8), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n569), .A2(new_n572), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n567), .B1(new_n260), .B2(new_n262), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n244), .A2(new_n324), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT82), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n571), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n570), .A2(KEYINPUT82), .A3(new_n350), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(KEYINPUT7), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT83), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT83), .ZN(new_n594));
  AOI211_X1 g408(.A(new_n594), .B(new_n591), .C1(new_n585), .C2(new_n586), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n584), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT84), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n584), .B(KEYINPUT84), .C1(new_n593), .C2(new_n595), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n530), .A2(new_n204), .A3(new_n532), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n578), .A3(new_n582), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT80), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n600), .A2(new_n578), .A3(KEYINPUT80), .A4(new_n582), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n598), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G210), .B1(G237), .B2(G902), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n582), .B1(new_n600), .B2(new_n578), .ZN(new_n608));
  OR2_X1    g422(.A1(new_n608), .A2(KEYINPUT6), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n608), .B1(new_n603), .B2(new_n604), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT6), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n587), .B(new_n571), .ZN(new_n613));
  AOI21_X1  g427(.A(G902), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n606), .A2(new_n607), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n607), .B1(new_n606), .B2(new_n614), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n564), .A2(new_n566), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n365), .A2(new_n496), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  NAND2_X1  g434(.A1(new_n308), .A2(new_n290), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G472), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n310), .ZN(new_n623));
  NOR4_X1   g437(.A1(new_n623), .A2(new_n564), .A3(new_n364), .A4(new_n495), .ZN(new_n624));
  INV_X1    g438(.A(new_n607), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n585), .A2(new_n586), .A3(new_n572), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n581), .A2(new_n583), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n594), .B1(new_n569), .B2(new_n591), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n587), .A2(KEYINPUT83), .A3(new_n592), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n605), .B1(new_n631), .B2(KEYINPUT84), .ZN(new_n632));
  INV_X1    g446(.A(new_n599), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n612), .A2(new_n613), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n290), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n625), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n606), .A2(new_n607), .A3(new_n614), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(KEYINPUT101), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n606), .A2(new_n640), .A3(new_n607), .A4(new_n614), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n641), .A2(new_n565), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n639), .A2(new_n642), .A3(KEYINPUT102), .ZN(new_n643));
  AOI21_X1  g457(.A(KEYINPUT102), .B1(new_n639), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n410), .A2(KEYINPUT103), .A3(new_n411), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(new_n420), .B2(G478), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n650), .B1(new_n405), .B2(new_n409), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n419), .A2(KEYINPUT33), .A3(new_n408), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n651), .A2(G478), .A3(new_n290), .A4(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n481), .A2(new_n486), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n624), .A2(new_n645), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT34), .B(G104), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  NAND3_X1  g471(.A1(new_n425), .A2(new_n426), .A3(new_n486), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n477), .A2(new_n478), .A3(new_n428), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n474), .A2(new_n475), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n624), .A2(new_n645), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NOR2_X1   g478(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n348), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n362), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n361), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n623), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n618), .A2(new_n670), .A3(new_n496), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n615), .A2(new_n616), .A3(new_n640), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n641), .A2(new_n565), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n639), .A2(new_n642), .A3(KEYINPUT102), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n677), .A2(new_n678), .A3(new_n668), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n299), .A2(new_n312), .A3(new_n313), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT104), .B(G900), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(new_n492), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n490), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n658), .A2(new_n660), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n564), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n680), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n237), .ZN(G30));
  NAND2_X1  g503(.A1(new_n287), .A2(new_n271), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n296), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n290), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n296), .B1(new_n293), .B2(new_n294), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n312), .A2(new_n313), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(KEYINPUT105), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n427), .A2(new_n487), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n697), .A2(new_n566), .A3(new_n668), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n698), .B(KEYINPUT106), .Z(new_n699));
  XOR2_X1   g513(.A(new_n683), .B(KEYINPUT39), .Z(new_n700));
  NOR2_X1   g514(.A1(new_n564), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT40), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n617), .B(KEYINPUT38), .Z(new_n703));
  AND4_X1   g517(.A1(new_n696), .A2(new_n699), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n231), .ZN(G45));
  AOI221_X4 g519(.A(new_n684), .B1(new_n649), .B2(new_n653), .C1(new_n481), .C2(new_n486), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n680), .A2(new_n686), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n645), .A3(new_n708), .A4(new_n668), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n680), .A2(new_n706), .A3(new_n686), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT107), .B1(new_n679), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  NAND2_X1  g527(.A1(new_n548), .A2(new_n290), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G469), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n563), .A3(new_n550), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n654), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n718), .A2(new_n364), .A3(new_n495), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n645), .A2(new_n680), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  NAND3_X1  g536(.A1(new_n677), .A2(new_n678), .A3(new_n717), .ZN(new_n723));
  INV_X1    g537(.A(new_n364), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n680), .A2(new_n724), .A3(new_n494), .A4(new_n661), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT109), .B(G116), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G18));
  INV_X1    g544(.A(new_n679), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n496), .A2(new_n680), .A3(new_n717), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  NAND2_X1  g548(.A1(new_n677), .A2(new_n678), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n697), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n295), .A2(new_n273), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n301), .B(new_n307), .C1(new_n737), .C2(new_n296), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n621), .A2(G472), .B1(new_n738), .B2(new_n309), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n724), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n740), .A2(new_n495), .A3(new_n716), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  NAND3_X1  g557(.A1(new_n706), .A2(new_n668), .A3(new_n739), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n723), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n316), .ZN(G27));
  NAND2_X1  g560(.A1(new_n617), .A2(new_n565), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n564), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(new_n680), .A3(new_n724), .A4(new_n706), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT111), .B1(KEYINPUT110), .B2(KEYINPUT42), .ZN(new_n750));
  OR2_X1    g564(.A1(KEYINPUT111), .A2(KEYINPUT42), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n749), .A2(new_n750), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n226), .ZN(G33));
  NAND2_X1  g569(.A1(new_n365), .A2(new_n748), .ZN(new_n756));
  INV_X1    g570(.A(new_n685), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n219), .ZN(G36));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n554), .A2(new_n556), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(KEYINPUT45), .ZN(new_n762));
  OAI21_X1  g576(.A(G469), .B1(new_n761), .B2(KEYINPUT45), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n760), .B1(new_n765), .B2(new_n558), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(KEYINPUT46), .A3(new_n559), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n550), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n700), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n563), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n747), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n649), .A2(new_n653), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n481), .A3(new_n486), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT112), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT43), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n623), .A3(new_n668), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n771), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT113), .B(G137), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G39));
  NAND2_X1  g596(.A1(new_n768), .A2(new_n563), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT47), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(KEYINPUT47), .ZN(new_n785));
  INV_X1    g599(.A(new_n747), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n314), .A2(new_n364), .A3(new_n706), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT114), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n784), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  NAND2_X1  g604(.A1(new_n784), .A2(new_n785), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n715), .A2(new_n562), .A3(new_n550), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n740), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n775), .A2(new_n489), .A3(new_n488), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n786), .A3(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n794), .A2(new_n717), .A3(new_n786), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n668), .A3(new_n739), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n696), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n716), .A2(new_n364), .A3(new_n490), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n786), .A3(new_n800), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n801), .A2(new_n487), .A3(new_n772), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n794), .A2(new_n724), .A3(new_n717), .A4(new_n739), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n565), .A3(new_n703), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n798), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n796), .A2(new_n365), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT48), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(KEYINPUT48), .ZN(new_n815));
  OAI221_X1 g629(.A(new_n488), .B1(new_n801), .B2(new_n718), .C1(new_n803), .C2(new_n735), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n810), .A2(new_n811), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n687), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n643), .A2(new_n644), .A3(new_n716), .ZN(new_n820));
  INV_X1    g634(.A(new_n744), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n731), .A2(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n564), .A2(new_n668), .A3(new_n684), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n736), .A2(new_n695), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n712), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT117), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n712), .A2(new_n822), .A3(new_n828), .A4(new_n824), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n825), .A2(KEYINPUT52), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n617), .A2(new_n566), .ZN(new_n834));
  INV_X1    g648(.A(new_n423), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n718), .B1(new_n487), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n624), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n619), .A2(new_n837), .A3(new_n671), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n736), .A2(new_n741), .B1(new_n731), .B2(new_n732), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n728), .A2(new_n720), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n821), .A2(new_n748), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n835), .A2(new_n486), .A3(new_n683), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n669), .A2(new_n842), .A3(new_n660), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n786), .A2(new_n843), .A3(new_n680), .A4(new_n686), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  OAI221_X1 g660(.A(new_n846), .B1(new_n757), .B2(new_n756), .C1(new_n753), .C2(new_n752), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT116), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n754), .A2(new_n758), .A3(new_n845), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n838), .A2(new_n720), .A3(new_n839), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n728), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n832), .A2(new_n833), .A3(new_n848), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n852), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n827), .B1(new_n826), .B2(new_n829), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT118), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n679), .A2(new_n687), .B1(new_n723), .B2(new_n744), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n709), .B2(new_n711), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n828), .B1(new_n859), .B2(new_n824), .ZN(new_n860));
  INV_X1    g674(.A(new_n829), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT52), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n863), .A3(new_n830), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n854), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n853), .B(KEYINPUT54), .C1(new_n865), .C2(new_n833), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  INV_X1    g681(.A(new_n840), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n832), .A2(KEYINPUT53), .A3(new_n868), .A4(new_n849), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n867), .B(new_n869), .C1(new_n865), .C2(KEYINPUT53), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n818), .A2(new_n871), .B1(G952), .B2(G953), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n724), .A2(new_n563), .A3(new_n565), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n715), .A2(new_n550), .ZN(new_n874));
  AOI211_X1 g688(.A(new_n773), .B(new_n873), .C1(KEYINPUT49), .C2(new_n874), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT115), .Z(new_n876));
  NOR2_X1   g690(.A1(new_n874), .A2(KEYINPUT49), .ZN(new_n877));
  OR4_X1    g691(.A1(new_n696), .A2(new_n876), .A3(new_n703), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n872), .A2(new_n878), .ZN(G75));
  XNOR2_X1  g693(.A(new_n612), .B(new_n613), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT55), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n869), .B1(new_n865), .B2(KEYINPUT53), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(G210), .A3(G902), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT56), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n883), .A2(new_n887), .A3(new_n884), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n881), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n881), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n350), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n889), .A2(new_n893), .ZN(G51));
  NAND2_X1  g708(.A1(new_n882), .A2(KEYINPUT54), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(KEYINPUT120), .A3(new_n870), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n882), .A2(new_n897), .A3(KEYINPUT54), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n558), .B(KEYINPUT57), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n548), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n882), .A2(G902), .A3(new_n765), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n891), .B1(new_n901), .B2(new_n902), .ZN(G54));
  NAND4_X1  g717(.A1(new_n882), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n904), .A2(new_n905), .A3(new_n476), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n892), .B1(new_n904), .B2(new_n476), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n905), .B1(new_n904), .B2(new_n476), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G60));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT59), .Z(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n866), .B2(new_n870), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n651), .A2(new_n652), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n892), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n896), .A2(new_n898), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n913), .A2(new_n911), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(G63));
  NAND2_X1  g732(.A1(G217), .A2(G902), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT60), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n882), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n354), .A2(new_n355), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n891), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT61), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n666), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n923), .B1(new_n926), .B2(new_n921), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI221_X1 g742(.A(new_n923), .B1(new_n924), .B2(KEYINPUT61), .C1(new_n926), .C2(new_n921), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(G66));
  NAND2_X1  g744(.A1(new_n491), .A2(new_n570), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n868), .B2(G953), .ZN(new_n933));
  OAI221_X1 g747(.A(new_n609), .B1(G898), .B2(new_n350), .C1(new_n610), .C2(new_n611), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G69));
  AOI21_X1  g749(.A(new_n350), .B1(G227), .B2(G900), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(KEYINPUT126), .ZN(new_n937));
  INV_X1    g751(.A(new_n770), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(new_n365), .A3(new_n736), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(KEYINPUT125), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n754), .A2(new_n758), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(KEYINPUT125), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n940), .A2(new_n789), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n780), .ZN(new_n944));
  INV_X1    g758(.A(new_n859), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n350), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n285), .A2(new_n286), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n459), .A2(new_n461), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT123), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(G900), .B2(G953), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n365), .A2(new_n769), .A3(new_n748), .A4(new_n836), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT124), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n789), .A2(new_n780), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n704), .A2(new_n945), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n952), .B1(new_n962), .B2(G953), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n937), .B1(new_n954), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n936), .A2(KEYINPUT126), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n964), .B(new_n965), .Z(G72));
  AND2_X1   g780(.A1(new_n946), .A2(new_n868), .ZN(new_n967));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n288), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n970), .B1(new_n962), .B2(new_n868), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n971), .B(new_n892), .C1(new_n972), .C2(new_n691), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n865), .A2(new_n833), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(new_n853), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n288), .A2(new_n970), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n976), .A2(new_n691), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n975), .A2(KEYINPUT127), .A3(new_n977), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n973), .B1(new_n980), .B2(new_n981), .ZN(G57));
endmodule


