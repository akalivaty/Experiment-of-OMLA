//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT68), .B(G244), .ZN(new_n210));
  AND2_X1   g0010(.A1(new_n210), .A2(G77), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G87), .A2(G250), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n209), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n209), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT0), .Z(new_n221));
  AOI21_X1  g0021(.A(KEYINPUT65), .B1(G1), .B2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND3_X1  g0023(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n207), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(new_n227));
  NOR2_X1   g0027(.A1(G58), .A2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT67), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(KEYINPUT67), .B1(G58), .B2(G68), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n230), .A2(G50), .A3(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n218), .B(new_n221), .C1(new_n227), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(G97), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G68), .ZN(new_n247));
  INV_X1    g0047(.A(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n245), .B(new_n252), .ZN(G351));
  OAI211_X1 g0053(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  OAI211_X1 g0056(.A(G1), .B(G13), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G232), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n254), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n262), .A2(new_n264), .A3(G223), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT81), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT81), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n268), .A2(new_n269), .A3(G223), .A4(new_n265), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G87), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n268), .A2(G226), .A3(G1698), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n267), .A2(new_n270), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n223), .B(new_n224), .C1(new_n255), .C2(new_n256), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n261), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G169), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n278), .B1(G179), .B2(new_n276), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  AND3_X1   g0080(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(new_n222), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT72), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT72), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n286), .A2(new_n206), .A3(G13), .A4(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT70), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n289), .B(new_n280), .C1(new_n281), .C2(new_n222), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n283), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT71), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT8), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(new_n293), .A3(G58), .ZN(new_n294));
  INV_X1    g0094(.A(G58), .ZN(new_n295));
  AOI21_X1  g0095(.A(KEYINPUT71), .B1(new_n295), .B2(KEYINPUT8), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(KEYINPUT8), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n291), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT73), .B1(new_n207), .B2(G1), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT73), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(new_n206), .A3(G20), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n298), .A2(new_n303), .B1(new_n287), .B2(new_n285), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT79), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT80), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT79), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n299), .A2(new_n309), .A3(new_n305), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  AOI211_X1 g0111(.A(KEYINPUT79), .B(new_n304), .C1(new_n291), .C2(new_n298), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n309), .B1(new_n299), .B2(new_n305), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT80), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n295), .A2(new_n248), .ZN(new_n316));
  OAI21_X1  g0116(.A(G20), .B1(new_n316), .B2(new_n228), .ZN(new_n317));
  NOR2_X1   g0117(.A1(G20), .A2(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G159), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT7), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n268), .B2(G20), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n262), .A2(new_n264), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(KEYINPUT16), .B(new_n321), .C1(new_n326), .C2(new_n248), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT16), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n248), .B1(new_n323), .B2(new_n325), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(new_n320), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n283), .A2(new_n290), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n327), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n279), .B1(new_n315), .B2(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n334), .A2(KEYINPUT18), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(KEYINPUT18), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n273), .A2(new_n275), .ZN(new_n338));
  INV_X1    g0138(.A(new_n261), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(G190), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n276), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT80), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n308), .B1(new_n307), .B2(new_n310), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n333), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT17), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n337), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G222), .A2(G1698), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n265), .A2(G223), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n268), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(G77), .B2(new_n268), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n274), .B1(new_n352), .B2(KEYINPUT69), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(KEYINPUT69), .B2(new_n352), .ZN(new_n354));
  INV_X1    g0154(.A(new_n254), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n257), .A2(new_n258), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n355), .B1(new_n356), .B2(G226), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n207), .A2(G33), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n298), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G150), .ZN(new_n365));
  INV_X1    g0165(.A(new_n318), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n364), .B1(new_n365), .B2(new_n366), .C1(new_n202), .C2(new_n207), .ZN(new_n367));
  INV_X1    g0167(.A(new_n288), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n367), .A2(new_n331), .B1(new_n246), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n283), .A2(new_n290), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(new_n288), .A3(new_n303), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(new_n371), .B2(new_n246), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n358), .A2(new_n277), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n361), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n371), .A2(new_n203), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT74), .ZN(new_n376));
  XOR2_X1   g0176(.A(KEYINPUT15), .B(G87), .Z(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n376), .B1(new_n378), .B2(new_n362), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(KEYINPUT74), .A3(new_n363), .ZN(new_n380));
  XOR2_X1   g0180(.A(KEYINPUT8), .B(G58), .Z(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n318), .B1(G20), .B2(G77), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n331), .B1(new_n203), .B2(new_n368), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n375), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n268), .A2(G238), .A3(G1698), .ZN(new_n386));
  INV_X1    g0186(.A(G107), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n268), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n324), .A2(new_n260), .A3(G1698), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n275), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n355), .B1(new_n356), .B2(new_n210), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n277), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n385), .B(new_n393), .C1(G179), .C2(new_n392), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(G200), .ZN(new_n395));
  INV_X1    g0195(.A(G190), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(new_n392), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n394), .B1(new_n385), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT9), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n372), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n372), .A2(new_n399), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n358), .A2(G200), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n359), .A2(G190), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n400), .A2(new_n401), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT10), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n403), .A2(new_n402), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT10), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n406), .A2(new_n407), .A3(new_n400), .A4(new_n401), .ZN(new_n408));
  AOI211_X1 g0208(.A(new_n374), .B(new_n398), .C1(new_n405), .C2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT78), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n368), .A2(new_n248), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT12), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n363), .A2(G77), .B1(G20), .B2(new_n248), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n246), .B2(new_n366), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n331), .A2(new_n414), .A3(KEYINPUT11), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n371), .A2(new_n248), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT11), .B1(new_n331), .B2(new_n414), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT77), .ZN(new_n420));
  NOR2_X1   g0220(.A1(G226), .A2(G1698), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n260), .B2(G1698), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n268), .B1(G33), .B2(G97), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n423), .A2(new_n274), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT13), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n254), .B(KEYINPUT75), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n356), .A2(G238), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n424), .A2(new_n425), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n427), .B(new_n426), .C1(new_n274), .C2(new_n423), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT13), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G169), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n431), .A2(new_n434), .A3(G169), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n428), .A2(new_n430), .A3(KEYINPUT76), .ZN(new_n437));
  OR3_X1    g0237(.A1(new_n429), .A2(KEYINPUT76), .A3(KEYINPUT13), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n360), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n420), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n434), .B1(new_n431), .B2(G169), .ZN(new_n441));
  AOI211_X1 g0241(.A(KEYINPUT14), .B(new_n277), .C1(new_n428), .C2(new_n430), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n439), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(KEYINPUT77), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n419), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n431), .A2(G200), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n419), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n396), .B1(new_n437), .B2(new_n438), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n410), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n419), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n436), .A2(new_n420), .A3(new_n439), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT77), .B1(new_n443), .B2(new_n444), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n450), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT78), .ZN(new_n457));
  AND4_X1   g0257(.A1(new_n348), .A2(new_n409), .A3(new_n451), .A4(new_n457), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT5), .B(G41), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  INV_X1    g0260(.A(G274), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n460), .A2(new_n461), .A3(G1), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n257), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n460), .A2(G1), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(new_n459), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n463), .B1(new_n466), .B2(G270), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n268), .A2(G257), .A3(new_n265), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n268), .A2(G264), .A3(G1698), .ZN(new_n469));
  INV_X1    g0269(.A(G303), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n468), .B(new_n469), .C1(new_n470), .C2(new_n268), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n275), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n467), .A2(new_n472), .A3(G179), .ZN(new_n473));
  AOI21_X1  g0273(.A(G20), .B1(G33), .B2(G283), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n255), .A2(G97), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n474), .A2(new_n475), .B1(G20), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(new_n282), .A3(KEYINPUT20), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT20), .B1(new_n477), .B2(new_n282), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n479), .A2(new_n480), .B1(G116), .B2(new_n288), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n206), .A2(G33), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n283), .A2(new_n288), .A3(new_n290), .A4(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n476), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT85), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n370), .A2(G116), .A3(new_n288), .A4(new_n482), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT85), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n477), .A2(new_n282), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n490), .A2(new_n478), .B1(new_n476), .B2(new_n368), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n486), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n473), .B1(new_n485), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n485), .A2(new_n492), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n467), .A2(new_n472), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G169), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT21), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n496), .A2(new_n499), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n494), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT86), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n501), .A2(new_n494), .A3(KEYINPUT86), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n268), .A2(new_n207), .A3(G87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT22), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT22), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n268), .A2(new_n508), .A3(new_n207), .A4(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n387), .A2(G20), .ZN(new_n511));
  OAI22_X1  g0311(.A1(KEYINPUT23), .A2(new_n511), .B1(new_n362), .B2(new_n476), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(KEYINPUT23), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT88), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n511), .A2(new_n515), .A3(KEYINPUT23), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n512), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT24), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n510), .A2(KEYINPUT24), .A3(new_n517), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n331), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n483), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT25), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n288), .B2(G107), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n368), .A2(KEYINPUT25), .A3(new_n387), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n523), .A2(G107), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n268), .A2(G257), .A3(G1698), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n268), .A2(G250), .A3(new_n265), .ZN(new_n530));
  INV_X1    g0330(.A(G294), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n529), .B(new_n530), .C1(new_n255), .C2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(new_n275), .B1(new_n466), .B2(G264), .ZN(new_n533));
  INV_X1    g0333(.A(new_n463), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n277), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n528), .B(new_n536), .C1(G179), .C2(new_n535), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n500), .A2(new_n504), .A3(new_n505), .A4(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n268), .A2(G244), .A3(G1698), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n268), .A2(G238), .A3(new_n265), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G116), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n275), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n464), .A2(new_n465), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n462), .B1(new_n545), .B2(G250), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n544), .A2(KEYINPUT84), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT84), .B1(new_n544), .B2(new_n546), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n360), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n544), .A2(new_n546), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT84), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n544), .A2(KEYINPUT84), .A3(new_n546), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n277), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n268), .A2(new_n207), .A3(G68), .ZN(new_n555));
  NAND3_X1  g0355(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n207), .ZN(new_n557));
  INV_X1    g0357(.A(G87), .ZN(new_n558));
  INV_X1    g0358(.A(G97), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n559), .A3(new_n387), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n362), .A2(new_n559), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n555), .B(new_n561), .C1(KEYINPUT19), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n331), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n368), .A2(new_n378), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n483), .C2(new_n378), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n549), .A2(new_n554), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(G190), .B1(new_n547), .B2(new_n548), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n552), .A2(G200), .A3(new_n553), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n565), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(G87), .B2(new_n523), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n535), .A2(G200), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n533), .A2(G190), .A3(new_n534), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n573), .A2(new_n522), .A3(new_n527), .A4(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n567), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n494), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT87), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n495), .A2(G200), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n472), .A2(G190), .A3(new_n467), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n577), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n579), .B1(new_n396), .B2(new_n495), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT87), .B1(new_n583), .B2(new_n494), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n268), .A2(G244), .A3(new_n265), .ZN(new_n586));
  NAND2_X1  g0386(.A1(KEYINPUT82), .A2(KEYINPUT4), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n262), .A2(new_n264), .A3(G250), .A4(G1698), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT83), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n268), .A2(KEYINPUT83), .A3(G250), .A4(G1698), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n588), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(KEYINPUT82), .A2(KEYINPUT4), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(G33), .B2(G283), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n586), .B2(new_n587), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n275), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n463), .B1(new_n466), .B2(G257), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n360), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT6), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n600), .A2(new_n559), .A3(G107), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n600), .B2(new_n244), .ZN(new_n602));
  OAI22_X1  g0402(.A1(new_n602), .A2(new_n207), .B1(new_n203), .B2(new_n366), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n387), .B1(new_n323), .B2(new_n325), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n331), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n368), .A2(new_n559), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n523), .A2(G97), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n597), .A2(new_n598), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n607), .A2(new_n608), .B1(new_n609), .B2(new_n277), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n605), .A3(new_n606), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(G200), .B2(new_n609), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n597), .A2(new_n598), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G190), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n599), .A2(new_n610), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n576), .A2(new_n585), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n458), .A2(new_n539), .A3(new_n616), .ZN(G372));
  NAND2_X1  g0417(.A1(new_n405), .A2(new_n408), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n455), .B1(new_n394), .B2(new_n450), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n619), .A2(new_n347), .ZN(new_n620));
  INV_X1    g0420(.A(new_n337), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n618), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n374), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n458), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n550), .A2(new_n277), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n549), .A2(new_n566), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n609), .A2(new_n277), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n629), .A2(new_n599), .A3(new_n611), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(new_n567), .A3(new_n572), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n628), .B1(new_n631), .B2(KEYINPUT26), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n550), .A2(G200), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n568), .A2(new_n571), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n627), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT89), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n629), .A2(new_n599), .A3(new_n611), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT89), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n635), .A2(new_n637), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT90), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n632), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n627), .A2(new_n634), .A3(new_n575), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n538), .A2(new_n615), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n643), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n624), .B1(new_n625), .B2(new_n649), .ZN(G369));
  AND3_X1   g0450(.A1(new_n500), .A2(new_n504), .A3(new_n505), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT91), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT91), .ZN(new_n656));
  INV_X1    g0456(.A(G213), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n652), .B2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n651), .A2(new_n585), .B1(new_n494), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n661), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n577), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n651), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(G330), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n651), .A2(new_n661), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n537), .A2(new_n661), .ZN(new_n669));
  INV_X1    g0469(.A(new_n575), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n663), .B1(new_n522), .B2(new_n527), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n537), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n669), .ZN(G399));
  INV_X1    g0476(.A(new_n219), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n560), .A2(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n232), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n552), .A2(new_n553), .ZN(new_n684));
  INV_X1    g0484(.A(new_n473), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n684), .A2(new_n613), .A3(new_n685), .A4(new_n533), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  AND4_X1   g0487(.A1(new_n360), .A2(new_n535), .A3(new_n495), .A4(new_n550), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n686), .A2(new_n687), .B1(new_n688), .B2(new_n609), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n687), .B2(new_n686), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT92), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n661), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n616), .A2(new_n539), .A3(new_n663), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(KEYINPUT31), .ZN(new_n696));
  OAI21_X1  g0496(.A(G330), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n647), .A2(KEYINPUT93), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT93), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n538), .A2(new_n700), .A3(new_n615), .A4(new_n646), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n630), .A2(new_n638), .A3(new_n567), .A4(new_n572), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n627), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n635), .A2(new_n637), .A3(new_n640), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n703), .B1(KEYINPUT26), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n699), .A2(new_n701), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT94), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(new_n707), .A3(new_n663), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n707), .B1(new_n706), .B2(new_n663), .ZN(new_n710));
  OAI21_X1  g0510(.A(KEYINPUT29), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n648), .A2(new_n663), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n698), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n683), .B1(new_n715), .B2(G1), .ZN(G364));
  NAND2_X1  g0516(.A1(new_n207), .A2(G13), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n206), .B1(new_n718), .B2(G45), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n678), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n225), .B1(G20), .B2(new_n277), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT95), .Z(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n219), .A2(G355), .A3(new_n268), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n677), .A2(new_n268), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G45), .B2(new_n232), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n252), .A2(new_n460), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n732), .B1(G116), .B2(new_n219), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n722), .B1(new_n731), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n360), .A2(new_n341), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n207), .A2(G190), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(KEYINPUT33), .A2(G317), .ZN(new_n742));
  AND2_X1   g0542(.A1(KEYINPUT33), .A2(G317), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n207), .A2(new_n396), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n360), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G322), .ZN(new_n749));
  INV_X1    g0549(.A(G283), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n341), .A2(G179), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n739), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n744), .B(new_n749), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n745), .A2(new_n751), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n739), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G303), .A2(new_n755), .B1(new_n758), .B2(G329), .ZN(new_n759));
  INV_X1    g0559(.A(G311), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n739), .A2(new_n746), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n759), .B(new_n324), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n738), .A2(new_n745), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT97), .Z(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT98), .B(G326), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n207), .B1(new_n756), .B2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n764), .A2(new_n765), .B1(G294), .B2(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n753), .B(new_n762), .C1(new_n768), .C2(KEYINPUT99), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n768), .A2(KEYINPUT99), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n766), .A2(new_n559), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(G68), .B2(new_n741), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT96), .Z(new_n773));
  NAND2_X1  g0573(.A1(new_n755), .A2(G87), .ZN(new_n774));
  INV_X1    g0574(.A(G159), .ZN(new_n775));
  OAI21_X1  g0575(.A(KEYINPUT32), .B1(new_n757), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n774), .A2(new_n268), .A3(new_n776), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n747), .A2(new_n295), .B1(new_n752), .B2(new_n387), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n763), .A2(new_n246), .B1(new_n761), .B2(new_n203), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n757), .A2(KEYINPUT32), .A3(new_n775), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n777), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n769), .A2(new_n770), .B1(new_n773), .B2(new_n781), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n737), .B1(new_n724), .B2(new_n782), .C1(new_n665), .C2(new_n728), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT100), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n665), .A2(G330), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n666), .A2(new_n785), .A3(new_n721), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n787), .A2(KEYINPUT101), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(KEYINPUT101), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(G396));
  OR2_X1    g0590(.A1(new_n394), .A2(new_n661), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n397), .A2(new_n385), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n663), .B1(new_n375), .B2(new_n384), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n394), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n712), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n795), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n648), .A2(new_n663), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n721), .B1(new_n799), .B2(new_n697), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n697), .B2(new_n799), .ZN(new_n801));
  INV_X1    g0601(.A(new_n752), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G87), .A2(new_n802), .B1(new_n758), .B2(G311), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n803), .B1(new_n387), .B2(new_n754), .C1(new_n470), .C2(new_n763), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n324), .B1(new_n761), .B2(new_n476), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n750), .A2(new_n740), .B1(new_n747), .B2(new_n531), .ZN(new_n806));
  NOR4_X1   g0606(.A1(new_n804), .A2(new_n771), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(KEYINPUT102), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT102), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n740), .A2(new_n365), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n763), .A2(new_n812), .B1(new_n761), .B2(new_n775), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n811), .B(new_n813), .C1(G143), .C2(new_n748), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n268), .B1(new_n757), .B2(new_n816), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n754), .A2(new_n246), .B1(new_n752), .B2(new_n248), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(G58), .C2(new_n767), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n807), .A2(new_n810), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n723), .B1(new_n809), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n723), .A2(new_n725), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n722), .B1(new_n824), .B2(new_n203), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n823), .B(new_n825), .C1(new_n797), .C2(new_n726), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n801), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G384));
  INV_X1    g0628(.A(KEYINPUT35), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n476), .B1(new_n602), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n227), .B(new_n830), .C1(new_n829), .C2(new_n602), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT36), .Z(new_n832));
  OR3_X1    g0632(.A1(new_n232), .A2(new_n203), .A3(new_n316), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n206), .B(G13), .C1(new_n833), .C2(new_n247), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n419), .A2(new_n663), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n455), .A2(new_n456), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n446), .A2(new_n661), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n795), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n691), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n696), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n329), .A2(new_n320), .ZN(new_n845));
  OR3_X1    g0645(.A1(new_n845), .A2(KEYINPUT103), .A3(KEYINPUT16), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(KEYINPUT103), .B2(KEYINPUT16), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n846), .A2(new_n331), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(new_n310), .A3(new_n307), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n279), .A2(new_n659), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n844), .B1(new_n851), .B2(new_n346), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n332), .B1(new_n311), .B2(new_n314), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n346), .B1(new_n854), .B2(new_n279), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT104), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n854), .B2(new_n659), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n333), .B1(new_n344), .B2(new_n345), .ZN(new_n858));
  INV_X1    g0658(.A(new_n659), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(KEYINPUT104), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n855), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT105), .B1(new_n861), .B2(new_n844), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(new_n857), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n332), .B(new_n342), .C1(new_n311), .C2(new_n314), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n334), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n863), .A2(new_n865), .A3(KEYINPUT105), .A4(new_n844), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n853), .B1(new_n862), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n849), .A2(new_n859), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n337), .B2(new_n347), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT38), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n863), .A2(new_n844), .A3(new_n865), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT105), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n852), .B1(new_n875), .B2(new_n866), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n876), .A2(new_n877), .A3(new_n870), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n843), .B1(new_n872), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(KEYINPUT107), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT107), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n871), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n877), .B1(new_n876), .B2(new_n870), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n842), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n882), .B1(new_n885), .B2(KEYINPUT40), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n348), .A2(new_n863), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n861), .A2(new_n844), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n875), .A2(new_n866), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(KEYINPUT106), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT106), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n875), .A2(new_n891), .A3(new_n866), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n887), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n883), .B1(new_n893), .B2(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n843), .A2(KEYINPUT40), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n881), .A2(new_n886), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n695), .A2(KEYINPUT31), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n693), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n691), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n897), .A2(new_n458), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n881), .A2(new_n886), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n894), .A2(new_n896), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(G330), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(G330), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n899), .B2(new_n691), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n907), .A2(new_n458), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n901), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n711), .A2(new_n458), .A3(new_n714), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n624), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n909), .B(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n621), .A2(new_n659), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n883), .A2(new_n884), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n798), .A2(new_n791), .ZN(new_n916));
  INV_X1    g0716(.A(new_n839), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n446), .A2(new_n450), .A3(new_n836), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n913), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n923), .B(new_n883), .C1(new_n893), .C2(KEYINPUT38), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n914), .A2(KEYINPUT39), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n455), .A2(new_n661), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n922), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n912), .A2(new_n929), .B1(new_n206), .B2(new_n718), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n912), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n835), .B1(new_n930), .B2(new_n931), .ZN(G367));
  NAND4_X1  g0732(.A1(new_n667), .A2(new_n674), .A3(new_n538), .A4(new_n615), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT42), .Z(new_n934));
  NAND2_X1  g0734(.A1(new_n611), .A2(new_n661), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n615), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n639), .B1(new_n936), .B2(new_n537), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT109), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n661), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n938), .B2(new_n937), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n571), .A2(new_n663), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n627), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n635), .B2(new_n941), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT108), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n934), .A2(new_n940), .B1(KEYINPUT43), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n666), .A2(new_n674), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n936), .B1(new_n639), .B2(new_n663), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n948), .B(new_n952), .Z(new_n953));
  INV_X1    g0753(.A(new_n715), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n668), .B(new_n673), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n667), .A2(new_n674), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n669), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n951), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT44), .Z(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(new_n951), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT45), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(new_n949), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n954), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n678), .B(KEYINPUT41), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n719), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n953), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n733), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n968), .A2(new_n241), .B1(new_n219), .B2(new_n378), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n721), .B1(new_n730), .B2(new_n969), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n754), .A2(new_n295), .B1(new_n761), .B2(new_n246), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n324), .B(new_n971), .C1(G150), .C2(new_n748), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n767), .A2(G68), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n764), .A2(G143), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n757), .A2(new_n812), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n752), .A2(new_n203), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n975), .B(new_n976), .C1(G159), .C2(new_n741), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n972), .A2(new_n973), .A3(new_n974), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(KEYINPUT111), .B1(new_n755), .B2(G116), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT46), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n324), .B1(new_n752), .B2(new_n559), .ZN(new_n981));
  INV_X1    g0781(.A(G317), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n747), .A2(new_n470), .B1(new_n757), .B2(new_n982), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n981), .B(new_n983), .C1(G294), .C2(new_n741), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n764), .A2(G311), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n980), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n761), .A2(new_n750), .B1(new_n766), .B2(new_n387), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT110), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n978), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT47), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n724), .B1(new_n989), .B2(new_n990), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n970), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n945), .B2(new_n728), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n967), .A2(new_n994), .ZN(G387));
  INV_X1    g0795(.A(new_n955), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(new_n954), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(new_n679), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n954), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n680), .A2(KEYINPUT112), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n680), .A2(KEYINPUT112), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n460), .B1(new_n248), .B2(new_n203), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT113), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(KEYINPUT113), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n381), .A2(new_n246), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT50), .Z(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n968), .B1(new_n238), .B2(G45), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n219), .A2(new_n268), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(G107), .B2(new_n219), .C1(new_n680), .C2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n722), .B1(new_n1013), .B2(new_n731), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n763), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1015), .A2(G159), .B1(new_n758), .B2(G150), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n741), .A2(new_n298), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n246), .C2(new_n747), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n378), .A2(new_n766), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n268), .B1(new_n752), .B2(new_n559), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n755), .A2(G77), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n248), .B2(new_n761), .ZN(new_n1022));
  NOR4_X1   g0822(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n324), .B1(new_n752), .B2(new_n476), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n761), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G311), .A2(new_n741), .B1(new_n1025), .B2(G303), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n982), .B2(new_n747), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G322), .B2(new_n764), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT48), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n754), .A2(new_n531), .B1(new_n766), .B2(new_n750), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(KEYINPUT49), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1024), .B(new_n1032), .C1(new_n758), .C2(new_n765), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(KEYINPUT49), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1023), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1014), .B1(new_n674), .B2(new_n728), .C1(new_n1035), .C2(new_n724), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n955), .B2(new_n720), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1000), .A2(new_n1038), .ZN(G393));
  AOI21_X1  g0839(.A(new_n679), .B1(new_n997), .B2(new_n962), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n959), .A2(new_n961), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(new_n949), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1040), .B1(new_n997), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n951), .A2(new_n727), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n968), .A2(new_n245), .B1(new_n559), .B2(new_n219), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n721), .B1(new_n730), .B2(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n763), .A2(new_n365), .B1(new_n747), .B2(new_n775), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT51), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G68), .A2(new_n755), .B1(new_n758), .B2(G143), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G50), .A2(new_n741), .B1(new_n1025), .B2(new_n381), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n766), .A2(new_n203), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n324), .B(new_n1051), .C1(G87), .C2(new_n802), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G283), .A2(new_n755), .B1(new_n758), .B2(G322), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1054), .B(new_n324), .C1(new_n387), .C2(new_n752), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT115), .Z(new_n1056));
  OAI22_X1  g0856(.A1(new_n763), .A2(new_n982), .B1(new_n747), .B2(new_n760), .ZN(new_n1057));
  XOR2_X1   g0857(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n767), .A2(G116), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G303), .A2(new_n741), .B1(new_n1025), .B2(G294), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1053), .B1(new_n1056), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1046), .B1(new_n1065), .B2(new_n723), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1042), .A2(new_n720), .B1(new_n1044), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1043), .A2(new_n1067), .ZN(G390));
  AND3_X1   g0868(.A1(new_n907), .A2(KEYINPUT116), .A3(new_n458), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT116), .B1(new_n907), .B2(new_n458), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1071), .A2(new_n910), .A3(new_n624), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n907), .A2(new_n797), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1073), .A2(new_n919), .B1(new_n698), .B2(new_n840), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n706), .A2(new_n663), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(KEYINPUT94), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n708), .A3(new_n791), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n794), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n919), .B1(new_n697), .B2(new_n795), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n907), .A2(new_n840), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n916), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1072), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n927), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n921), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n924), .A2(new_n1087), .A3(new_n925), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1077), .A2(new_n794), .A3(new_n920), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n894), .A2(new_n1089), .A3(new_n1086), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n698), .A2(new_n840), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1081), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1085), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1081), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1071), .A2(new_n910), .A3(new_n624), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1074), .A2(new_n1078), .B1(new_n1082), .B2(new_n916), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1094), .A2(new_n1102), .A3(new_n678), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n824), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT54), .B(G143), .Z(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1106), .A2(new_n761), .B1(new_n812), .B2(new_n740), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G159), .B2(new_n767), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT117), .Z(new_n1109));
  AOI21_X1  g0909(.A(new_n324), .B1(new_n748), .B2(G132), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT119), .Z(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n365), .B2(new_n754), .ZN(new_n1114));
  INV_X1    g0914(.A(G125), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n752), .A2(new_n246), .B1(new_n757), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G128), .B2(new_n1015), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1112), .A2(G150), .A3(new_n755), .ZN(new_n1118));
  AND4_X1   g0918(.A1(new_n1110), .A2(new_n1114), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n774), .A2(new_n324), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT120), .Z(new_n1121));
  OAI22_X1  g0921(.A1(new_n763), .A2(new_n750), .B1(new_n747), .B2(new_n476), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n248), .A2(new_n752), .B1(new_n761), .B2(new_n559), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n740), .A2(new_n387), .B1(new_n757), .B2(new_n531), .ZN(new_n1124));
  NOR4_X1   g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .A4(new_n1051), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1109), .A2(new_n1119), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n721), .B1(new_n298), .B2(new_n1104), .C1(new_n1126), .C2(new_n724), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n926), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n725), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n720), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1103), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT121), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1103), .A2(new_n1131), .A3(KEYINPUT121), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(G378));
  NAND2_X1  g0936(.A1(new_n1102), .A2(new_n1072), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n372), .A2(new_n859), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n618), .A2(new_n623), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1138), .B1(new_n618), .B2(new_n623), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1143), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1140), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT123), .ZN(new_n1148));
  AND4_X1   g0948(.A1(G330), .A2(new_n902), .A3(new_n903), .A4(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1147), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n897), .B2(G330), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n928), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n897), .A2(G330), .A3(new_n1148), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n929), .B(new_n1153), .C1(new_n905), .C2(new_n1150), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1137), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT57), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1137), .A2(new_n1152), .A3(new_n1154), .A4(KEYINPUT57), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n678), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1152), .A2(new_n1154), .A3(new_n720), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n722), .B1(new_n824), .B2(new_n246), .ZN(new_n1161));
  INV_X1    g0961(.A(G128), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1162), .A2(new_n747), .B1(new_n740), .B2(new_n816), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n755), .A2(new_n1105), .B1(new_n1025), .B2(G137), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1115), .B2(new_n763), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(G150), .C2(new_n767), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT59), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n752), .A2(new_n775), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n255), .A2(new_n256), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT122), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G124), .C2(new_n758), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1168), .A2(new_n1169), .A3(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G107), .A2(new_n748), .B1(new_n802), .B2(G58), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n268), .A2(G41), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1175), .A2(new_n973), .A3(new_n1021), .A4(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n763), .A2(new_n476), .B1(new_n757), .B2(new_n750), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n378), .A2(new_n761), .B1(new_n559), .B2(new_n740), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1172), .B(new_n246), .C1(G41), .C2(new_n268), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1183));
  AND4_X1   g0983(.A1(new_n1174), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1161), .B1(new_n724), .B2(new_n1184), .C1(new_n1148), .C2(new_n726), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1160), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1159), .A2(new_n1187), .ZN(G375));
  NAND3_X1  g0988(.A1(new_n1084), .A2(KEYINPUT124), .A3(new_n720), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT124), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1099), .B2(new_n719), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n722), .B1(new_n824), .B2(new_n248), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n763), .A2(new_n531), .B1(new_n761), .B2(new_n387), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(G116), .B2(new_n741), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT125), .Z(new_n1195));
  AOI22_X1  g0995(.A1(G97), .A2(new_n755), .B1(new_n748), .B2(G283), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n470), .B2(new_n757), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1197), .A2(new_n268), .A3(new_n976), .A4(new_n1019), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n1106), .A2(new_n740), .B1(new_n761), .B2(new_n365), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n754), .A2(new_n775), .B1(new_n757), .B2(new_n1162), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n268), .B1(new_n752), .B2(new_n295), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n763), .A2(new_n816), .B1(new_n747), .B2(new_n812), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(G50), .C2(new_n767), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1195), .A2(new_n1198), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1192), .B1(new_n724), .B2(new_n1205), .C1(new_n920), .C2(new_n726), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1189), .A2(new_n1191), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1085), .A2(new_n964), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT126), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(G381));
  AND2_X1   g1012(.A1(new_n1158), .A2(new_n678), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1186), .B1(new_n1213), .B2(new_n1157), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1132), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n967), .A2(new_n994), .A3(new_n1043), .A4(new_n1067), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G393), .A2(G396), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1211), .A2(new_n827), .A3(new_n1218), .ZN(new_n1219));
  OR3_X1    g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1219), .ZN(G407));
  OAI211_X1 g1020(.A(G407), .B(G213), .C1(G343), .C2(new_n1216), .ZN(G409));
  INV_X1    g1021(.A(KEYINPUT61), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n657), .A2(G343), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1159), .A2(G378), .A3(new_n1187), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1155), .A2(new_n965), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1215), .B1(new_n1225), .B2(new_n1186), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1223), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT60), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1208), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1098), .A2(new_n1099), .A3(KEYINPUT60), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n678), .A3(new_n1085), .A4(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1231), .A2(new_n1207), .A3(G384), .ZN(new_n1232));
  AOI21_X1  g1032(.A(G384), .B1(new_n1231), .B2(new_n1207), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1223), .A2(G2897), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1235), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1232), .A2(new_n1233), .A3(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1222), .B1(new_n1227), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1227), .A2(new_n1234), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT63), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G387), .A2(G390), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1217), .ZN(new_n1247));
  INV_X1    g1047(.A(G396), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1000), .B2(new_n1038), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1218), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1246), .B(new_n1217), .C1(new_n1218), .C2(new_n1249), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1227), .A2(KEYINPUT63), .A3(new_n1234), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1242), .A2(new_n1245), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT62), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1227), .A2(new_n1257), .A3(new_n1234), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1257), .B1(new_n1227), .B2(new_n1234), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1258), .A2(new_n1241), .A3(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1256), .B1(new_n1260), .B2(new_n1254), .ZN(G405));
  INV_X1    g1061(.A(KEYINPUT127), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1224), .B(new_n1262), .C1(new_n1214), .C2(new_n1132), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n1253), .A3(new_n1234), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1253), .B1(new_n1263), .B2(new_n1234), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G375), .A2(new_n1215), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1262), .B1(new_n1267), .B2(new_n1224), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1265), .A2(new_n1266), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1263), .A2(new_n1234), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1254), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1268), .B1(new_n1272), .B2(new_n1264), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1270), .A2(new_n1273), .ZN(G402));
endmodule


