

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U560 ( .A1(G651), .A2(G543), .ZN(n653) );
  NOR2_X2 U561 ( .A1(n534), .A2(n640), .ZN(n590) );
  OR2_X1 U562 ( .A1(n775), .A2(n1021), .ZN(n527) );
  AND2_X1 U563 ( .A1(n562), .A2(n561), .ZN(n528) );
  INV_X1 U564 ( .A(n792), .ZN(n775) );
  INV_X1 U565 ( .A(KEYINPUT29), .ZN(n772) );
  XNOR2_X1 U566 ( .A(n772), .B(KEYINPUT99), .ZN(n773) );
  NAND2_X1 U567 ( .A1(n734), .A2(n733), .ZN(n792) );
  NOR2_X2 U568 ( .A1(G2104), .A2(n543), .ZN(n906) );
  NOR2_X1 U569 ( .A1(G651), .A2(n640), .ZN(n658) );
  NOR2_X1 U570 ( .A1(n552), .A2(n551), .ZN(G160) );
  NAND2_X1 U571 ( .A1(n653), .A2(G89), .ZN(n529) );
  XNOR2_X1 U572 ( .A(n529), .B(KEYINPUT4), .ZN(n532) );
  INV_X1 U573 ( .A(G651), .ZN(n534) );
  XOR2_X1 U574 ( .A(G543), .B(KEYINPUT0), .Z(n530) );
  XNOR2_X1 U575 ( .A(KEYINPUT66), .B(n530), .ZN(n640) );
  NAND2_X1 U576 ( .A1(G76), .A2(n590), .ZN(n531) );
  NAND2_X1 U577 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U578 ( .A(n533), .B(KEYINPUT5), .ZN(n540) );
  NOR2_X1 U579 ( .A1(G543), .A2(n534), .ZN(n535) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n535), .Z(n657) );
  NAND2_X1 U581 ( .A1(G63), .A2(n657), .ZN(n537) );
  NAND2_X1 U582 ( .A1(G51), .A2(n658), .ZN(n536) );
  NAND2_X1 U583 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U584 ( .A(KEYINPUT6), .B(n538), .Z(n539) );
  NAND2_X1 U585 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U586 ( .A(n541), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U587 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U588 ( .A(G2105), .ZN(n543) );
  NAND2_X1 U589 ( .A1(G125), .A2(n906), .ZN(n542) );
  XNOR2_X1 U590 ( .A(n542), .B(KEYINPUT64), .ZN(n546) );
  AND2_X1 U591 ( .A1(n543), .A2(G2104), .ZN(n901) );
  NAND2_X1 U592 ( .A1(G101), .A2(n901), .ZN(n544) );
  XOR2_X1 U593 ( .A(KEYINPUT23), .B(n544), .Z(n545) );
  NAND2_X1 U594 ( .A1(n546), .A2(n545), .ZN(n552) );
  AND2_X1 U595 ( .A1(G2104), .A2(G2105), .ZN(n905) );
  NAND2_X1 U596 ( .A1(G113), .A2(n905), .ZN(n550) );
  XNOR2_X1 U597 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n548) );
  NOR2_X1 U598 ( .A1(G2104), .A2(G2105), .ZN(n547) );
  XNOR2_X2 U599 ( .A(n548), .B(n547), .ZN(n902) );
  NAND2_X1 U600 ( .A1(G137), .A2(n902), .ZN(n549) );
  NAND2_X1 U601 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U602 ( .A1(G64), .A2(n657), .ZN(n554) );
  NAND2_X1 U603 ( .A1(G52), .A2(n658), .ZN(n553) );
  NAND2_X1 U604 ( .A1(n554), .A2(n553), .ZN(n560) );
  NAND2_X1 U605 ( .A1(G77), .A2(n590), .ZN(n556) );
  NAND2_X1 U606 ( .A1(G90), .A2(n653), .ZN(n555) );
  NAND2_X1 U607 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U608 ( .A(KEYINPUT68), .B(n557), .Z(n558) );
  XNOR2_X1 U609 ( .A(KEYINPUT9), .B(n558), .ZN(n559) );
  NOR2_X1 U610 ( .A1(n560), .A2(n559), .ZN(G171) );
  AND2_X1 U611 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U612 ( .A(G108), .ZN(G238) );
  INV_X1 U613 ( .A(G120), .ZN(G236) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  NAND2_X1 U615 ( .A1(n902), .A2(G138), .ZN(n565) );
  NAND2_X1 U616 ( .A1(G102), .A2(n901), .ZN(n562) );
  NAND2_X1 U617 ( .A1(G114), .A2(n905), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G126), .A2(n906), .ZN(n563) );
  AND2_X1 U619 ( .A1(n528), .A2(n563), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n565), .A2(n564), .ZN(n567) );
  INV_X1 U621 ( .A(KEYINPUT86), .ZN(n566) );
  XNOR2_X1 U622 ( .A(n567), .B(n566), .ZN(G164) );
  NAND2_X1 U623 ( .A1(G75), .A2(n590), .ZN(n569) );
  NAND2_X1 U624 ( .A1(G62), .A2(n657), .ZN(n568) );
  NAND2_X1 U625 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U626 ( .A1(G88), .A2(n653), .ZN(n570) );
  XNOR2_X1 U627 ( .A(KEYINPUT81), .B(n570), .ZN(n571) );
  NOR2_X1 U628 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U629 ( .A1(n658), .A2(G50), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n574), .A2(n573), .ZN(G303) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U632 ( .A(n575), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U633 ( .A(G567), .ZN(n687) );
  NOR2_X1 U634 ( .A1(G223), .A2(n687), .ZN(n577) );
  XNOR2_X1 U635 ( .A(KEYINPUT70), .B(KEYINPUT11), .ZN(n576) );
  XNOR2_X1 U636 ( .A(n577), .B(n576), .ZN(G234) );
  NAND2_X1 U637 ( .A1(n657), .A2(G56), .ZN(n578) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n578), .Z(n586) );
  NAND2_X1 U639 ( .A1(G68), .A2(n590), .ZN(n582) );
  XOR2_X1 U640 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n580) );
  NAND2_X1 U641 ( .A1(G81), .A2(n653), .ZN(n579) );
  XNOR2_X1 U642 ( .A(n580), .B(n579), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U644 ( .A(n583), .B(KEYINPUT72), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT13), .B(n584), .Z(n585) );
  NOR2_X1 U646 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U647 ( .A1(n658), .A2(G43), .ZN(n587) );
  NAND2_X1 U648 ( .A1(n588), .A2(n587), .ZN(n1020) );
  INV_X1 U649 ( .A(n1020), .ZN(n589) );
  NAND2_X1 U650 ( .A1(n589), .A2(G860), .ZN(G153) );
  INV_X1 U651 ( .A(G171), .ZN(G301) );
  NAND2_X1 U652 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U653 ( .A1(G79), .A2(n590), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G66), .A2(n657), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U656 ( .A1(G92), .A2(n653), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G54), .A2(n658), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U659 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U660 ( .A(KEYINPUT15), .B(n597), .Z(n1018) );
  OR2_X1 U661 ( .A1(n1018), .A2(G868), .ZN(n598) );
  NAND2_X1 U662 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U663 ( .A1(G78), .A2(n590), .ZN(n601) );
  NAND2_X1 U664 ( .A1(G65), .A2(n657), .ZN(n600) );
  NAND2_X1 U665 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U666 ( .A1(G53), .A2(n658), .ZN(n602) );
  XNOR2_X1 U667 ( .A(KEYINPUT69), .B(n602), .ZN(n603) );
  NOR2_X1 U668 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U669 ( .A1(n653), .A2(G91), .ZN(n605) );
  NAND2_X1 U670 ( .A1(n606), .A2(n605), .ZN(G299) );
  INV_X1 U671 ( .A(G868), .ZN(n672) );
  NOR2_X1 U672 ( .A1(G286), .A2(n672), .ZN(n608) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U674 ( .A1(n608), .A2(n607), .ZN(G297) );
  INV_X1 U675 ( .A(G559), .ZN(n609) );
  NOR2_X1 U676 ( .A1(G860), .A2(n609), .ZN(n610) );
  XNOR2_X1 U677 ( .A(KEYINPUT73), .B(n610), .ZN(n611) );
  NAND2_X1 U678 ( .A1(n611), .A2(n1018), .ZN(n612) );
  XNOR2_X1 U679 ( .A(n612), .B(KEYINPUT16), .ZN(n613) );
  XNOR2_X1 U680 ( .A(KEYINPUT74), .B(n613), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n1020), .ZN(n616) );
  NAND2_X1 U682 ( .A1(G868), .A2(n1018), .ZN(n614) );
  NOR2_X1 U683 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U684 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U685 ( .A1(n901), .A2(G99), .ZN(n617) );
  XNOR2_X1 U686 ( .A(KEYINPUT76), .B(n617), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n905), .A2(G111), .ZN(n618) );
  XOR2_X1 U688 ( .A(KEYINPUT75), .B(n618), .Z(n619) );
  NAND2_X1 U689 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U690 ( .A(n621), .B(KEYINPUT77), .ZN(n623) );
  NAND2_X1 U691 ( .A1(G135), .A2(n902), .ZN(n622) );
  NAND2_X1 U692 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U693 ( .A1(n906), .A2(G123), .ZN(n624) );
  XOR2_X1 U694 ( .A(KEYINPUT18), .B(n624), .Z(n625) );
  NOR2_X1 U695 ( .A1(n626), .A2(n625), .ZN(n1001) );
  XNOR2_X1 U696 ( .A(G2096), .B(n1001), .ZN(n628) );
  INV_X1 U697 ( .A(G2100), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n628), .A2(n627), .ZN(G156) );
  NAND2_X1 U699 ( .A1(G80), .A2(n590), .ZN(n630) );
  NAND2_X1 U700 ( .A1(G67), .A2(n657), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U702 ( .A1(G93), .A2(n653), .ZN(n632) );
  NAND2_X1 U703 ( .A1(G55), .A2(n658), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n633) );
  OR2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n671) );
  XNOR2_X1 U706 ( .A(n1020), .B(KEYINPUT78), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n1018), .A2(G559), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(n669) );
  NOR2_X1 U709 ( .A1(n669), .A2(G860), .ZN(n637) );
  XOR2_X1 U710 ( .A(KEYINPUT79), .B(n637), .Z(n638) );
  XOR2_X1 U711 ( .A(n671), .B(n638), .Z(G145) );
  NAND2_X1 U712 ( .A1(G49), .A2(n658), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n639), .B(KEYINPUT80), .ZN(n645) );
  NAND2_X1 U714 ( .A1(G651), .A2(G74), .ZN(n642) );
  NAND2_X1 U715 ( .A1(G87), .A2(n640), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U717 ( .A1(n657), .A2(n643), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n645), .A2(n644), .ZN(G288) );
  NAND2_X1 U719 ( .A1(G86), .A2(n653), .ZN(n647) );
  NAND2_X1 U720 ( .A1(G61), .A2(n657), .ZN(n646) );
  NAND2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n590), .A2(G73), .ZN(n648) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n648), .Z(n649) );
  NOR2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n658), .A2(G48), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n652), .A2(n651), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G72), .A2(n590), .ZN(n655) );
  NAND2_X1 U728 ( .A1(G85), .A2(n653), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U730 ( .A(KEYINPUT67), .B(n656), .ZN(n662) );
  NAND2_X1 U731 ( .A1(G60), .A2(n657), .ZN(n660) );
  NAND2_X1 U732 ( .A1(G47), .A2(n658), .ZN(n659) );
  AND2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U734 ( .A1(n662), .A2(n661), .ZN(G290) );
  INV_X1 U735 ( .A(G303), .ZN(G166) );
  XOR2_X1 U736 ( .A(n671), .B(G288), .Z(n668) );
  XNOR2_X1 U737 ( .A(KEYINPUT82), .B(KEYINPUT19), .ZN(n664) );
  XNOR2_X1 U738 ( .A(G290), .B(G166), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n664), .B(n663), .ZN(n665) );
  XOR2_X1 U740 ( .A(n665), .B(G299), .Z(n666) );
  XNOR2_X1 U741 ( .A(G305), .B(n666), .ZN(n667) );
  XNOR2_X1 U742 ( .A(n668), .B(n667), .ZN(n920) );
  XNOR2_X1 U743 ( .A(n669), .B(n920), .ZN(n670) );
  NAND2_X1 U744 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U745 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U746 ( .A1(n674), .A2(n673), .ZN(G295) );
  INV_X1 U747 ( .A(G2072), .ZN(n760) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XOR2_X1 U751 ( .A(KEYINPUT21), .B(n677), .Z(n678) );
  NOR2_X1 U752 ( .A1(n760), .A2(n678), .ZN(n679) );
  XNOR2_X1 U753 ( .A(KEYINPUT83), .B(n679), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U755 ( .A1(G132), .A2(G82), .ZN(n680) );
  XNOR2_X1 U756 ( .A(n680), .B(KEYINPUT22), .ZN(n681) );
  XNOR2_X1 U757 ( .A(n681), .B(KEYINPUT84), .ZN(n682) );
  NOR2_X1 U758 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U759 ( .A1(G96), .A2(n683), .ZN(n855) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n855), .ZN(n684) );
  XNOR2_X1 U761 ( .A(n684), .B(KEYINPUT85), .ZN(n689) );
  NOR2_X1 U762 ( .A1(G236), .A2(G238), .ZN(n685) );
  NAND2_X1 U763 ( .A1(G69), .A2(n685), .ZN(n686) );
  NOR2_X1 U764 ( .A1(G237), .A2(n686), .ZN(n857) );
  NOR2_X1 U765 ( .A1(n687), .A2(n857), .ZN(n688) );
  NOR2_X1 U766 ( .A1(n689), .A2(n688), .ZN(G319) );
  INV_X1 U767 ( .A(G319), .ZN(n691) );
  NAND2_X1 U768 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U769 ( .A1(n691), .A2(n690), .ZN(n852) );
  NAND2_X1 U770 ( .A1(n852), .A2(G36), .ZN(G176) );
  XOR2_X1 U771 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n716) );
  XOR2_X1 U772 ( .A(KEYINPUT38), .B(KEYINPUT92), .Z(n693) );
  NAND2_X1 U773 ( .A1(G105), .A2(n901), .ZN(n692) );
  XNOR2_X1 U774 ( .A(n693), .B(n692), .ZN(n697) );
  NAND2_X1 U775 ( .A1(G117), .A2(n905), .ZN(n695) );
  NAND2_X1 U776 ( .A1(G141), .A2(n902), .ZN(n694) );
  NAND2_X1 U777 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U778 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U779 ( .A1(n906), .A2(G129), .ZN(n698) );
  NAND2_X1 U780 ( .A1(n699), .A2(n698), .ZN(n897) );
  NOR2_X1 U781 ( .A1(G1996), .A2(n897), .ZN(n992) );
  NAND2_X1 U782 ( .A1(n902), .A2(G131), .ZN(n700) );
  XOR2_X1 U783 ( .A(KEYINPUT89), .B(n700), .Z(n702) );
  NAND2_X1 U784 ( .A1(n901), .A2(G95), .ZN(n701) );
  NAND2_X1 U785 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U786 ( .A(KEYINPUT90), .B(n703), .ZN(n707) );
  NAND2_X1 U787 ( .A1(G107), .A2(n905), .ZN(n705) );
  NAND2_X1 U788 ( .A1(G119), .A2(n906), .ZN(n704) );
  NAND2_X1 U789 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U790 ( .A1(n707), .A2(n706), .ZN(n896) );
  XNOR2_X1 U791 ( .A(KEYINPUT91), .B(G1991), .ZN(n941) );
  NOR2_X1 U792 ( .A1(n896), .A2(n941), .ZN(n709) );
  AND2_X1 U793 ( .A1(n897), .A2(G1996), .ZN(n708) );
  NOR2_X1 U794 ( .A1(n709), .A2(n708), .ZN(n1004) );
  NOR2_X1 U795 ( .A1(G1384), .A2(G164), .ZN(n734) );
  NAND2_X1 U796 ( .A1(G160), .A2(G40), .ZN(n732) );
  NOR2_X1 U797 ( .A1(n734), .A2(n732), .ZN(n710) );
  XNOR2_X1 U798 ( .A(KEYINPUT87), .B(n710), .ZN(n717) );
  NOR2_X1 U799 ( .A1(n1004), .A2(n717), .ZN(n737) );
  NAND2_X1 U800 ( .A1(n896), .A2(n941), .ZN(n711) );
  XOR2_X1 U801 ( .A(KEYINPUT104), .B(n711), .Z(n996) );
  NOR2_X1 U802 ( .A1(G1986), .A2(G290), .ZN(n712) );
  NOR2_X1 U803 ( .A1(n996), .A2(n712), .ZN(n713) );
  NOR2_X1 U804 ( .A1(n737), .A2(n713), .ZN(n714) );
  NOR2_X1 U805 ( .A1(n992), .A2(n714), .ZN(n715) );
  XNOR2_X1 U806 ( .A(n716), .B(n715), .ZN(n728) );
  INV_X1 U807 ( .A(n717), .ZN(n844) );
  NAND2_X1 U808 ( .A1(G104), .A2(n901), .ZN(n719) );
  NAND2_X1 U809 ( .A1(G140), .A2(n902), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U811 ( .A(KEYINPUT34), .B(n720), .ZN(n726) );
  NAND2_X1 U812 ( .A1(n905), .A2(G116), .ZN(n721) );
  XNOR2_X1 U813 ( .A(n721), .B(KEYINPUT88), .ZN(n723) );
  NAND2_X1 U814 ( .A1(G128), .A2(n906), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U816 ( .A(KEYINPUT35), .B(n724), .Z(n725) );
  NOR2_X1 U817 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U818 ( .A(KEYINPUT36), .B(n727), .ZN(n917) );
  XNOR2_X1 U819 ( .A(G2067), .B(KEYINPUT37), .ZN(n729) );
  NOR2_X1 U820 ( .A1(n917), .A2(n729), .ZN(n997) );
  NAND2_X1 U821 ( .A1(n844), .A2(n997), .ZN(n738) );
  NAND2_X1 U822 ( .A1(n728), .A2(n738), .ZN(n730) );
  NAND2_X1 U823 ( .A1(n917), .A2(n729), .ZN(n994) );
  NAND2_X1 U824 ( .A1(n730), .A2(n994), .ZN(n731) );
  NAND2_X1 U825 ( .A1(n731), .A2(n844), .ZN(n843) );
  INV_X1 U826 ( .A(n732), .ZN(n733) );
  NAND2_X1 U827 ( .A1(G8), .A2(n792), .ZN(n828) );
  NOR2_X1 U828 ( .A1(G1981), .A2(G305), .ZN(n735) );
  XOR2_X1 U829 ( .A(n735), .B(KEYINPUT24), .Z(n736) );
  NOR2_X1 U830 ( .A1(n828), .A2(n736), .ZN(n742) );
  OR2_X1 U831 ( .A1(n742), .A2(n828), .ZN(n740) );
  INV_X1 U832 ( .A(n737), .ZN(n739) );
  AND2_X1 U833 ( .A1(n739), .A2(n738), .ZN(n821) );
  AND2_X1 U834 ( .A1(n740), .A2(n821), .ZN(n807) );
  INV_X1 U835 ( .A(n807), .ZN(n746) );
  NOR2_X1 U836 ( .A1(G2090), .A2(G303), .ZN(n741) );
  NAND2_X1 U837 ( .A1(G8), .A2(n741), .ZN(n744) );
  INV_X1 U838 ( .A(n742), .ZN(n743) );
  AND2_X1 U839 ( .A1(n744), .A2(n743), .ZN(n745) );
  OR2_X1 U840 ( .A1(n746), .A2(n745), .ZN(n747) );
  AND2_X1 U841 ( .A1(n843), .A2(n747), .ZN(n810) );
  XOR2_X1 U842 ( .A(G1996), .B(KEYINPUT95), .Z(n951) );
  NAND2_X1 U843 ( .A1(n775), .A2(n951), .ZN(n748) );
  XNOR2_X1 U844 ( .A(n748), .B(KEYINPUT26), .ZN(n749) );
  INV_X1 U845 ( .A(G1341), .ZN(n1021) );
  NAND2_X1 U846 ( .A1(n749), .A2(n527), .ZN(n750) );
  NOR2_X1 U847 ( .A1(n750), .A2(n1020), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n756), .A2(n1018), .ZN(n755) );
  AND2_X1 U849 ( .A1(n775), .A2(G2067), .ZN(n751) );
  XOR2_X1 U850 ( .A(n751), .B(KEYINPUT96), .Z(n753) );
  NAND2_X1 U851 ( .A1(n792), .A2(G1348), .ZN(n752) );
  NAND2_X1 U852 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U853 ( .A1(n755), .A2(n754), .ZN(n758) );
  OR2_X1 U854 ( .A1(n756), .A2(n1018), .ZN(n757) );
  NAND2_X1 U855 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U856 ( .A(n759), .B(KEYINPUT97), .ZN(n766) );
  NOR2_X1 U857 ( .A1(n792), .A2(n760), .ZN(n762) );
  XNOR2_X1 U858 ( .A(KEYINPUT27), .B(KEYINPUT94), .ZN(n761) );
  XNOR2_X1 U859 ( .A(n762), .B(n761), .ZN(n764) );
  NAND2_X1 U860 ( .A1(n792), .A2(G1956), .ZN(n763) );
  NAND2_X1 U861 ( .A1(n764), .A2(n763), .ZN(n768) );
  NOR2_X1 U862 ( .A1(G299), .A2(n768), .ZN(n765) );
  NOR2_X1 U863 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U864 ( .A(KEYINPUT98), .B(n767), .ZN(n771) );
  NAND2_X1 U865 ( .A1(G299), .A2(n768), .ZN(n769) );
  XOR2_X1 U866 ( .A(n769), .B(KEYINPUT28), .Z(n770) );
  NOR2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n774) );
  XNOR2_X1 U868 ( .A(n774), .B(n773), .ZN(n780) );
  XOR2_X1 U869 ( .A(G2078), .B(KEYINPUT25), .Z(n945) );
  NOR2_X1 U870 ( .A1(n945), .A2(n792), .ZN(n777) );
  NOR2_X1 U871 ( .A1(n775), .A2(G1961), .ZN(n776) );
  NOR2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U873 ( .A(KEYINPUT93), .B(n778), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G171), .A2(n784), .ZN(n779) );
  NAND2_X1 U875 ( .A1(n780), .A2(n779), .ZN(n789) );
  NOR2_X1 U876 ( .A1(G1966), .A2(n828), .ZN(n802) );
  NOR2_X1 U877 ( .A1(G2084), .A2(n792), .ZN(n801) );
  NOR2_X1 U878 ( .A1(n802), .A2(n801), .ZN(n781) );
  NAND2_X1 U879 ( .A1(G8), .A2(n781), .ZN(n782) );
  XNOR2_X1 U880 ( .A(KEYINPUT30), .B(n782), .ZN(n783) );
  NOR2_X1 U881 ( .A1(G168), .A2(n783), .ZN(n786) );
  NOR2_X1 U882 ( .A1(G171), .A2(n784), .ZN(n785) );
  NOR2_X1 U883 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U884 ( .A(KEYINPUT31), .B(n787), .Z(n788) );
  NAND2_X1 U885 ( .A1(n789), .A2(n788), .ZN(n806) );
  NAND2_X1 U886 ( .A1(n806), .A2(G286), .ZN(n790) );
  XNOR2_X1 U887 ( .A(n790), .B(KEYINPUT100), .ZN(n797) );
  NOR2_X1 U888 ( .A1(G1971), .A2(n828), .ZN(n791) );
  XNOR2_X1 U889 ( .A(KEYINPUT101), .B(n791), .ZN(n795) );
  NOR2_X1 U890 ( .A1(G2090), .A2(n792), .ZN(n793) );
  NOR2_X1 U891 ( .A1(G166), .A2(n793), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U894 ( .A(n798), .B(KEYINPUT102), .ZN(n799) );
  NAND2_X1 U895 ( .A1(n799), .A2(G8), .ZN(n800) );
  XNOR2_X1 U896 ( .A(KEYINPUT32), .B(n800), .ZN(n824) );
  NAND2_X1 U897 ( .A1(G8), .A2(n801), .ZN(n804) );
  INV_X1 U898 ( .A(n802), .ZN(n803) );
  AND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n811) );
  AND2_X1 U901 ( .A1(n811), .A2(n807), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n824), .A2(n808), .ZN(n809) );
  AND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n842) );
  NAND2_X1 U904 ( .A1(G1976), .A2(G288), .ZN(n1029) );
  AND2_X1 U905 ( .A1(n811), .A2(n1029), .ZN(n813) );
  INV_X1 U906 ( .A(KEYINPUT33), .ZN(n831) );
  AND2_X1 U907 ( .A1(n831), .A2(KEYINPUT103), .ZN(n834) );
  INV_X1 U908 ( .A(n834), .ZN(n812) );
  AND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n820) );
  INV_X1 U910 ( .A(KEYINPUT103), .ZN(n815) );
  NOR2_X1 U911 ( .A1(G1976), .A2(G288), .ZN(n1026) );
  NAND2_X1 U912 ( .A1(n1026), .A2(KEYINPUT33), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n1026), .A2(KEYINPUT103), .ZN(n816) );
  NAND2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U916 ( .A1(n828), .A2(n818), .ZN(n836) );
  INV_X1 U917 ( .A(n836), .ZN(n819) );
  AND2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n822) );
  XOR2_X1 U919 ( .A(G1981), .B(G305), .Z(n1015) );
  AND2_X1 U920 ( .A1(n1015), .A2(n821), .ZN(n825) );
  AND2_X1 U921 ( .A1(n822), .A2(n825), .ZN(n823) );
  NAND2_X1 U922 ( .A1(n824), .A2(n823), .ZN(n840) );
  INV_X1 U923 ( .A(n825), .ZN(n838) );
  INV_X1 U924 ( .A(n1029), .ZN(n830) );
  NOR2_X1 U925 ( .A1(G303), .A2(G1971), .ZN(n826) );
  NOR2_X1 U926 ( .A1(n826), .A2(n1026), .ZN(n827) );
  OR2_X1 U927 ( .A1(n828), .A2(n827), .ZN(n829) );
  OR2_X1 U928 ( .A1(n830), .A2(n829), .ZN(n832) );
  AND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(n833) );
  OR2_X1 U930 ( .A1(n834), .A2(n833), .ZN(n835) );
  OR2_X1 U931 ( .A1(n836), .A2(n835), .ZN(n837) );
  OR2_X1 U932 ( .A1(n838), .A2(n837), .ZN(n839) );
  AND2_X1 U933 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U934 ( .A1(n842), .A2(n841), .ZN(n848) );
  INV_X1 U935 ( .A(n843), .ZN(n846) );
  XNOR2_X1 U936 ( .A(G1986), .B(G290), .ZN(n1032) );
  NAND2_X1 U937 ( .A1(n1032), .A2(n844), .ZN(n845) );
  OR2_X1 U938 ( .A1(n846), .A2(n845), .ZN(n847) );
  AND2_X1 U939 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U940 ( .A(KEYINPUT40), .B(n849), .ZN(G329) );
  INV_X1 U941 ( .A(G223), .ZN(n850) );
  NAND2_X1 U942 ( .A1(G2106), .A2(n850), .ZN(G217) );
  AND2_X1 U943 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U944 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U945 ( .A1(G3), .A2(G1), .ZN(n853) );
  NAND2_X1 U946 ( .A1(n853), .A2(n852), .ZN(n854) );
  XOR2_X1 U947 ( .A(KEYINPUT107), .B(n854), .Z(G188) );
  INV_X1 U949 ( .A(G132), .ZN(G219) );
  INV_X1 U950 ( .A(G82), .ZN(G220) );
  INV_X1 U951 ( .A(n855), .ZN(n856) );
  NAND2_X1 U952 ( .A1(n857), .A2(n856), .ZN(G261) );
  INV_X1 U953 ( .A(G261), .ZN(G325) );
  XOR2_X1 U954 ( .A(G2678), .B(G2096), .Z(n859) );
  XNOR2_X1 U955 ( .A(KEYINPUT108), .B(G2100), .ZN(n858) );
  XNOR2_X1 U956 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U957 ( .A(n860), .B(KEYINPUT109), .Z(n862) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2090), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U960 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n864) );
  XNOR2_X1 U961 ( .A(G2072), .B(KEYINPUT43), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U963 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U964 ( .A(G2078), .B(G2084), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n868), .B(n867), .ZN(G227) );
  XOR2_X1 U966 ( .A(G1976), .B(G1971), .Z(n870) );
  XNOR2_X1 U967 ( .A(G1996), .B(G1986), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U969 ( .A(G1981), .B(G1961), .Z(n872) );
  XNOR2_X1 U970 ( .A(G1966), .B(G1956), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(n874), .B(n873), .Z(n876) );
  XNOR2_X1 U973 ( .A(G2474), .B(KEYINPUT41), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n878) );
  XOR2_X1 U975 ( .A(G1991), .B(KEYINPUT111), .Z(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(G229) );
  NAND2_X1 U977 ( .A1(G124), .A2(n906), .ZN(n879) );
  XNOR2_X1 U978 ( .A(n879), .B(KEYINPUT44), .ZN(n881) );
  NAND2_X1 U979 ( .A1(n901), .A2(G100), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n885) );
  NAND2_X1 U981 ( .A1(G112), .A2(n905), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G136), .A2(n902), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  NOR2_X1 U984 ( .A1(n885), .A2(n884), .ZN(G162) );
  XNOR2_X1 U985 ( .A(G160), .B(G162), .ZN(n894) );
  NAND2_X1 U986 ( .A1(G118), .A2(n905), .ZN(n887) );
  NAND2_X1 U987 ( .A1(G130), .A2(n906), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n892) );
  NAND2_X1 U989 ( .A1(G106), .A2(n901), .ZN(n889) );
  NAND2_X1 U990 ( .A1(G142), .A2(n902), .ZN(n888) );
  NAND2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U992 ( .A(KEYINPUT45), .B(n890), .Z(n891) );
  NOR2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n916) );
  XOR2_X1 U996 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n899) );
  XOR2_X1 U997 ( .A(n897), .B(KEYINPUT112), .Z(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n1001), .B(n900), .ZN(n914) );
  NAND2_X1 U1000 ( .A1(G103), .A2(n901), .ZN(n904) );
  NAND2_X1 U1001 ( .A1(G139), .A2(n902), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(n911) );
  NAND2_X1 U1003 ( .A1(G115), .A2(n905), .ZN(n908) );
  NAND2_X1 U1004 ( .A1(G127), .A2(n906), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1006 ( .A(KEYINPUT47), .B(n909), .Z(n910) );
  NOR2_X1 U1007 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1008 ( .A(KEYINPUT113), .B(n912), .Z(n987) );
  XNOR2_X1 U1009 ( .A(G164), .B(n987), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n918) );
  XOR2_X1 U1012 ( .A(n918), .B(n917), .Z(n919) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n919), .ZN(G395) );
  XNOR2_X1 U1014 ( .A(G171), .B(G286), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(n921), .B(n920), .ZN(n923) );
  XOR2_X1 U1016 ( .A(n1020), .B(n1018), .Z(n922) );
  XNOR2_X1 U1017 ( .A(n923), .B(n922), .ZN(n924) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n924), .ZN(G397) );
  XOR2_X1 U1019 ( .A(G2438), .B(G2435), .Z(n926) );
  XNOR2_X1 U1020 ( .A(G2443), .B(KEYINPUT106), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(n926), .B(n925), .ZN(n927) );
  XOR2_X1 U1022 ( .A(n927), .B(G2454), .Z(n929) );
  XNOR2_X1 U1023 ( .A(G1341), .B(G1348), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(n929), .B(n928), .ZN(n933) );
  XOR2_X1 U1025 ( .A(G2451), .B(G2427), .Z(n931) );
  XNOR2_X1 U1026 ( .A(G2430), .B(G2446), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(n931), .B(n930), .ZN(n932) );
  XOR2_X1 U1028 ( .A(n933), .B(n932), .Z(n934) );
  NAND2_X1 U1029 ( .A1(G14), .A2(n934), .ZN(n940) );
  NAND2_X1 U1030 ( .A1(G319), .A2(n940), .ZN(n937) );
  NOR2_X1 U1031 ( .A1(G227), .A2(G229), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(KEYINPUT49), .B(n935), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(G395), .A2(G397), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(G225) );
  INV_X1 U1036 ( .A(G225), .ZN(G308) );
  INV_X1 U1037 ( .A(G69), .ZN(G235) );
  INV_X1 U1038 ( .A(G96), .ZN(G221) );
  INV_X1 U1039 ( .A(n940), .ZN(G401) );
  XNOR2_X1 U1040 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n1051) );
  XOR2_X1 U1041 ( .A(KEYINPUT55), .B(KEYINPUT117), .Z(n961) );
  XNOR2_X1 U1042 ( .A(G2090), .B(G35), .ZN(n956) );
  XNOR2_X1 U1043 ( .A(G25), .B(n941), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(G33), .B(G2072), .ZN(n942) );
  NOR2_X1 U1046 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1047 ( .A1(G28), .A2(n944), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(G27), .B(n945), .ZN(n946) );
  XNOR2_X1 U1049 ( .A(KEYINPUT116), .B(n946), .ZN(n947) );
  NOR2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(G32), .B(n951), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1054 ( .A(KEYINPUT53), .B(n954), .ZN(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1056 ( .A(G2084), .B(G34), .Z(n957) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n957), .ZN(n958) );
  NAND2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1059 ( .A(n961), .B(n960), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(G29), .A2(n962), .ZN(n1049) );
  XNOR2_X1 U1061 ( .A(G1971), .B(G22), .ZN(n964) );
  XNOR2_X1 U1062 ( .A(G23), .B(G1976), .ZN(n963) );
  NOR2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1064 ( .A(KEYINPUT124), .B(n965), .Z(n967) );
  XNOR2_X1 U1065 ( .A(G1986), .B(G24), .ZN(n966) );
  NOR2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(KEYINPUT58), .B(n968), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G21), .ZN(n970) );
  XNOR2_X1 U1069 ( .A(G5), .B(G1961), .ZN(n969) );
  NOR2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(KEYINPUT59), .B(G1348), .ZN(n973) );
  XNOR2_X1 U1073 ( .A(n973), .B(G4), .ZN(n979) );
  XOR2_X1 U1074 ( .A(G1956), .B(G20), .Z(n975) );
  XNOR2_X1 U1075 ( .A(n1021), .B(G19), .ZN(n974) );
  NAND2_X1 U1076 ( .A1(n975), .A2(n974), .ZN(n977) );
  XNOR2_X1 U1077 ( .A(G6), .B(G1981), .ZN(n976) );
  NOR2_X1 U1078 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1079 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1080 ( .A(KEYINPUT60), .B(n980), .Z(n981) );
  XNOR2_X1 U1081 ( .A(KEYINPUT123), .B(n981), .ZN(n982) );
  NOR2_X1 U1082 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1083 ( .A(KEYINPUT61), .B(n984), .Z(n985) );
  NOR2_X1 U1084 ( .A1(G16), .A2(n985), .ZN(n986) );
  XOR2_X1 U1085 ( .A(KEYINPUT125), .B(n986), .Z(n1046) );
  XOR2_X1 U1086 ( .A(G2072), .B(n987), .Z(n989) );
  XOR2_X1 U1087 ( .A(G164), .B(G2078), .Z(n988) );
  NOR2_X1 U1088 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1089 ( .A(KEYINPUT50), .B(n990), .ZN(n1008) );
  XOR2_X1 U1090 ( .A(G2090), .B(G162), .Z(n991) );
  NOR2_X1 U1091 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1092 ( .A(KEYINPUT51), .B(n993), .Z(n995) );
  NAND2_X1 U1093 ( .A1(n995), .A2(n994), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G160), .B(G2084), .ZN(n999) );
  NOR2_X1 U1095 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1096 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1097 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1098 ( .A(n1002), .B(KEYINPUT114), .ZN(n1003) );
  NAND2_X1 U1099 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1100 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1102 ( .A(n1009), .B(KEYINPUT52), .ZN(n1010) );
  XNOR2_X1 U1103 ( .A(KEYINPUT115), .B(n1010), .ZN(n1012) );
  INV_X1 U1104 ( .A(KEYINPUT55), .ZN(n1011) );
  NAND2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1106 ( .A1(n1013), .A2(G29), .ZN(n1044) );
  XNOR2_X1 U1107 ( .A(G1966), .B(G168), .ZN(n1014) );
  XNOR2_X1 U1108 ( .A(n1014), .B(KEYINPUT118), .ZN(n1016) );
  NAND2_X1 U1109 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1110 ( .A(n1017), .B(KEYINPUT57), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(n1018), .B(G1348), .ZN(n1019) );
  XNOR2_X1 U1112 ( .A(n1019), .B(KEYINPUT119), .ZN(n1023) );
  XOR2_X1 U1113 ( .A(n1021), .B(n1020), .Z(n1022) );
  NOR2_X1 U1114 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1115 ( .A1(n1025), .A2(n1024), .ZN(n1039) );
  XNOR2_X1 U1116 ( .A(G171), .B(G1961), .ZN(n1037) );
  XNOR2_X1 U1117 ( .A(G299), .B(G1956), .ZN(n1028) );
  XNOR2_X1 U1118 ( .A(n1026), .B(KEYINPUT120), .ZN(n1027) );
  NOR2_X1 U1119 ( .A1(n1028), .A2(n1027), .ZN(n1034) );
  XNOR2_X1 U1120 ( .A(G166), .B(G1971), .ZN(n1030) );
  NAND2_X1 U1121 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1122 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1123 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1124 ( .A(KEYINPUT121), .B(n1035), .ZN(n1036) );
  NAND2_X1 U1125 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1126 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XOR2_X1 U1127 ( .A(KEYINPUT122), .B(n1040), .Z(n1042) );
  XNOR2_X1 U1128 ( .A(G16), .B(KEYINPUT56), .ZN(n1041) );
  NAND2_X1 U1129 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NAND2_X1 U1130 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  NOR2_X1 U1131 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  NAND2_X1 U1132 ( .A1(n1047), .A2(G11), .ZN(n1048) );
  NOR2_X1 U1133 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  XNOR2_X1 U1134 ( .A(n1051), .B(n1050), .ZN(n1052) );
  XNOR2_X1 U1135 ( .A(KEYINPUT62), .B(n1052), .ZN(G150) );
  INV_X1 U1136 ( .A(G150), .ZN(G311) );
endmodule

