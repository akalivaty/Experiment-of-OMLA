//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941;
  XOR2_X1   g000(.A(KEYINPUT82), .B(G50gat), .Z(new_n202));
  INV_X1    g001(.A(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G141gat), .B(G148gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(KEYINPUT2), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT76), .B(G162gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G141gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G148gat), .ZN(new_n214));
  INV_X1    g013(.A(G148gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G141gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n204), .B(new_n206), .C1(new_n214), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n209), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT77), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g019(.A(KEYINPUT77), .B(new_n209), .C1(new_n212), .C2(new_n217), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223));
  XNOR2_X1  g022(.A(G197gat), .B(G204gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT22), .ZN(new_n225));
  INV_X1    g024(.A(G211gat), .ZN(new_n226));
  INV_X1    g025(.A(G218gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G211gat), .B(G218gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n230), .B1(new_n228), .B2(new_n224), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n223), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n222), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G228gat), .ZN(new_n238));
  INV_X1    g037(.A(G233gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n232), .A2(new_n233), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n235), .B(new_n209), .C1(new_n212), .C2(new_n217), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n241), .B1(new_n243), .B2(KEYINPUT29), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n237), .A2(new_n240), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT81), .ZN(new_n246));
  INV_X1    g045(.A(new_n240), .ZN(new_n247));
  INV_X1    g046(.A(new_n244), .ZN(new_n248));
  INV_X1    g047(.A(new_n218), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n249), .B1(new_n235), .B2(new_n234), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n247), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT81), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n237), .A2(new_n252), .A3(new_n240), .A4(new_n244), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n246), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G22gat), .ZN(new_n255));
  INV_X1    g054(.A(G22gat), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n246), .A2(new_n251), .A3(new_n256), .A4(new_n253), .ZN(new_n257));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n258), .B1(new_n255), .B2(new_n257), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n202), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n255), .A2(new_n257), .ZN(new_n263));
  INV_X1    g062(.A(new_n258), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n202), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n259), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n262), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n268), .B1(new_n262), .B2(new_n267), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n273));
  INV_X1    g072(.A(G134gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G127gat), .ZN(new_n275));
  INV_X1    g074(.A(G127gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G134gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(G113gat), .B(G120gat), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n279), .B(new_n280), .C1(KEYINPUT1), .C2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n283));
  XNOR2_X1  g082(.A(G127gat), .B(G134gat), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G113gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT70), .B1(new_n285), .B2(G120gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n283), .B(new_n284), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n282), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n292), .B1(new_n282), .B2(new_n291), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n273), .B1(new_n295), .B2(new_n218), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n282), .A2(new_n291), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(new_n218), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT4), .ZN(new_n299));
  INV_X1    g098(.A(new_n221), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n207), .A2(new_n208), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n203), .A2(KEYINPUT76), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT76), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G162gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n304), .A3(G155gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT77), .B1(new_n307), .B2(new_n209), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT3), .B1(new_n300), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n242), .B1(new_n309), .B2(KEYINPUT78), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n235), .B1(new_n220), .B2(new_n221), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT78), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n297), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n296), .B(new_n299), .C1(new_n310), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(KEYINPUT5), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n249), .B(KEYINPUT4), .C1(new_n293), .C2(new_n294), .ZN(new_n319));
  OAI22_X1  g118(.A1(new_n297), .A2(new_n218), .B1(new_n273), .B2(new_n316), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n282), .A2(new_n291), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n322), .B1(new_n309), .B2(KEYINPUT78), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n243), .B1(new_n311), .B2(new_n312), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n322), .B1(new_n220), .B2(new_n221), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(new_n298), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT5), .B1(new_n327), .B2(new_n315), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n314), .A2(new_n318), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT0), .B(G57gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G85gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G1gat), .B(G29gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n331), .B(new_n332), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT6), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n321), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n310), .B2(new_n313), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT5), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n326), .A2(new_n298), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(new_n316), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n324), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n344), .A2(new_n317), .A3(new_n296), .A4(new_n299), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n345), .A3(new_n333), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n346), .A2(new_n336), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n329), .A2(KEYINPUT84), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT84), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n334), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n337), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT87), .B(KEYINPUT35), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n272), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n356));
  AND2_X1   g155(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n357));
  AND2_X1   g156(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n359));
  OAI22_X1  g158(.A1(new_n356), .A2(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT28), .ZN(new_n361));
  NAND2_X1  g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT66), .B(G190gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT27), .B(G183gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n361), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT68), .ZN(new_n368));
  NAND2_X1  g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT26), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(KEYINPUT26), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n367), .A2(new_n368), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n361), .A2(new_n374), .A3(new_n362), .A4(new_n366), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT68), .B1(new_n376), .B2(new_n372), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT67), .ZN(new_n379));
  INV_X1    g178(.A(G183gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n357), .B2(new_n356), .ZN(new_n381));
  NAND3_X1  g180(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT24), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT23), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n370), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n385), .A2(KEYINPUT25), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391));
  AND2_X1   g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(KEYINPUT24), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n384), .A2(KEYINPUT65), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT65), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT25), .B1(new_n398), .B2(new_n389), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n379), .B1(new_n390), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT25), .A3(new_n389), .ZN(new_n401));
  INV_X1    g200(.A(new_n388), .ZN(new_n402));
  NOR3_X1   g201(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n369), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n395), .B(KEYINPUT65), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n404), .B1(new_n405), .B2(new_n393), .ZN(new_n406));
  OAI211_X1 g205(.A(KEYINPUT67), .B(new_n401), .C1(new_n406), .C2(KEYINPUT25), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n378), .A2(new_n408), .A3(new_n295), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n295), .B1(new_n378), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT64), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n409), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT72), .B1(new_n414), .B2(KEYINPUT33), .ZN(new_n415));
  XNOR2_X1  g214(.A(G15gat), .B(G43gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(G71gat), .ZN(new_n417));
  INV_X1    g216(.A(G99gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n378), .A2(new_n408), .ZN(new_n420));
  INV_X1    g219(.A(new_n295), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n377), .A2(new_n375), .B1(new_n400), .B2(new_n407), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n295), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n424), .A3(new_n412), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT32), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT72), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n415), .A2(new_n419), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n419), .A2(KEYINPUT33), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n425), .A2(KEYINPUT32), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n422), .A2(new_n424), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT34), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n413), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n433), .B2(new_n413), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n430), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n430), .B2(new_n432), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n444), .B(KEYINPUT74), .Z(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n376), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT25), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n392), .A2(KEYINPUT65), .A3(KEYINPUT24), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n382), .B1(G183gat), .B2(G190gat), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n396), .B1(new_n362), .B2(new_n383), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n448), .B1(new_n452), .B2(new_n404), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n447), .A2(new_n373), .B1(new_n453), .B2(new_n401), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n446), .B1(new_n454), .B2(KEYINPUT29), .ZN(new_n455));
  INV_X1    g254(.A(new_n241), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n455), .B(new_n456), .C1(new_n423), .C2(new_n446), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n445), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n446), .A2(new_n223), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n241), .B(new_n458), .C1(new_n423), .C2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n460), .A3(KEYINPUT75), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n420), .A2(new_n223), .A3(new_n446), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT75), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n462), .A2(new_n463), .A3(new_n241), .A4(new_n458), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(G8gat), .B(G36gat), .Z(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(G64gat), .ZN(new_n467));
  INV_X1    g266(.A(G92gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n461), .A2(new_n464), .A3(new_n469), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(KEYINPUT30), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT30), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n465), .A2(new_n474), .A3(new_n470), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n443), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n335), .A2(KEYINPUT79), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT79), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n329), .A2(new_n480), .A3(new_n334), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n347), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n337), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n272), .A2(new_n484), .A3(new_n476), .A4(new_n442), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n355), .A2(new_n478), .B1(new_n485), .B2(KEYINPUT35), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n430), .A2(new_n432), .ZN(new_n487));
  INV_X1    g286(.A(new_n438), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT73), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n489), .B(new_n439), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  OAI22_X1  g293(.A1(new_n440), .A2(new_n441), .B1(new_n490), .B2(new_n491), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n268), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n260), .A2(new_n261), .A3(new_n202), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n266), .B1(new_n265), .B2(new_n259), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n501), .A2(new_n269), .B1(new_n484), .B2(new_n476), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n497), .A2(KEYINPUT83), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n504));
  INV_X1    g303(.A(new_n484), .ZN(new_n505));
  OAI22_X1  g304(.A1(new_n270), .A2(new_n271), .B1(new_n505), .B2(new_n477), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n506), .B2(new_n496), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n455), .B(new_n241), .C1(new_n423), .C2(new_n446), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n456), .B(new_n458), .C1(new_n423), .C2(new_n459), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT37), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT85), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT37), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n470), .B1(new_n465), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT38), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n351), .A2(new_n347), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n483), .A4(new_n471), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT86), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n514), .B1(new_n513), .B2(new_n465), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT38), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT86), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n352), .A2(new_n522), .A3(new_n471), .A4(new_n516), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n314), .A2(new_n316), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n327), .A2(new_n315), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n525), .A2(KEYINPUT39), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT39), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n314), .A2(new_n528), .A3(new_n316), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n333), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT40), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n525), .A2(KEYINPUT39), .A3(new_n526), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT40), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n333), .A4(new_n529), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n535), .A2(new_n475), .A3(new_n473), .A4(new_n351), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n536), .A2(new_n501), .A3(new_n269), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n524), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n486), .B1(new_n508), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT10), .ZN(new_n540));
  OR2_X1    g339(.A1(G57gat), .A2(G64gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(G57gat), .A2(G64gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(G71gat), .A2(G78gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n544), .A2(KEYINPUT9), .ZN(new_n545));
  NOR2_X1   g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  OAI22_X1  g345(.A1(new_n543), .A2(new_n545), .B1(KEYINPUT96), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n544), .A2(new_n546), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552));
  INV_X1    g351(.A(G85gat), .ZN(new_n553));
  AOI22_X1  g352(.A1(KEYINPUT8), .A2(new_n552), .B1(new_n553), .B2(new_n468), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n549), .B1(KEYINPUT99), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G99gat), .B(G106gat), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n555), .B(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT100), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n540), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n557), .A2(new_n559), .ZN(new_n563));
  INV_X1    g362(.A(new_n549), .ZN(new_n564));
  OAI211_X1 g363(.A(KEYINPUT100), .B(KEYINPUT10), .C1(new_n564), .C2(new_n559), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n563), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n569), .B2(new_n560), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G120gat), .B(G148gat), .Z(new_n572));
  XNOR2_X1  g371(.A(G176gat), .B(G204gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n568), .A2(new_n570), .A3(new_n576), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G15gat), .B(G22gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT91), .ZN(new_n583));
  INV_X1    g382(.A(G1gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n586));
  AOI21_X1  g385(.A(G8gat), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n584), .A2(KEYINPUT16), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n585), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n587), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G43gat), .B(G50gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT15), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT89), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n591), .A2(KEYINPUT15), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G29gat), .A2(G36gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT88), .ZN(new_n597));
  OR3_X1    g396(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n598), .A2(KEYINPUT90), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(KEYINPUT90), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n597), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n597), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n598), .A2(new_n600), .ZN(new_n605));
  OAI211_X1 g404(.A(KEYINPUT15), .B(new_n591), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n590), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT17), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n607), .B(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n608), .B1(new_n610), .B2(new_n590), .ZN(new_n611));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT93), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT18), .B1(new_n614), .B2(KEYINPUT94), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(KEYINPUT94), .B2(new_n614), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n590), .B(new_n607), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n613), .B(KEYINPUT13), .Z(new_n618));
  AOI22_X1  g417(.A1(new_n614), .A2(KEYINPUT18), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT11), .B(G169gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G197gat), .ZN(new_n622));
  XOR2_X1   g421(.A(G113gat), .B(G141gat), .Z(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  INV_X1    g424(.A(KEYINPUT95), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n619), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n620), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n620), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT21), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n590), .B1(new_n632), .B2(new_n564), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n380), .ZN(new_n634));
  XOR2_X1   g433(.A(G127gat), .B(G155gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT97), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT98), .B(G211gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n636), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n564), .A2(new_n632), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n641), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n610), .A2(new_n559), .ZN(new_n647));
  NAND3_X1  g446(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n647), .B(new_n648), .C1(new_n559), .C2(new_n607), .ZN(new_n649));
  XOR2_X1   g448(.A(G134gat), .B(G162gat), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G190gat), .B(G218gat), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n651), .B(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n646), .A2(new_n656), .ZN(new_n657));
  NOR4_X1   g456(.A1(new_n539), .A2(new_n581), .A3(new_n631), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n505), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n477), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT16), .B(G8gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT42), .Z(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(G8gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(G1325gat));
  AOI21_X1  g466(.A(G15gat), .B1(new_n658), .B2(new_n442), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT104), .Z(new_n669));
  NOR2_X1   g468(.A1(new_n492), .A2(new_n493), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n440), .A2(new_n441), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n492), .B1(new_n489), .B2(new_n439), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT105), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n494), .A2(new_n495), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n677), .A2(G15gat), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n669), .B1(new_n658), .B2(new_n678), .ZN(G1326gat));
  INV_X1    g478(.A(new_n272), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n658), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  INV_X1    g482(.A(new_n539), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n631), .A2(new_n581), .A3(new_n646), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n684), .A2(new_n655), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(G29gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n686), .A2(new_n687), .A3(new_n505), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT45), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT44), .B1(new_n539), .B2(new_n656), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n355), .A2(new_n478), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694));
  AND4_X1   g493(.A1(new_n694), .A2(new_n676), .A3(new_n538), .A4(new_n506), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n502), .B1(new_n673), .B2(new_n675), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n694), .B1(new_n696), .B2(new_n538), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n693), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n699), .A3(new_n655), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n690), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n685), .ZN(new_n702));
  OAI21_X1  g501(.A(G29gat), .B1(new_n702), .B2(new_n484), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n689), .A2(new_n703), .ZN(G1328gat));
  INV_X1    g503(.A(G36gat), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n686), .A2(new_n705), .A3(new_n477), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT46), .Z(new_n707));
  OAI21_X1  g506(.A(G36gat), .B1(new_n702), .B2(new_n476), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1329gat));
  INV_X1    g508(.A(G43gat), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n686), .A2(new_n710), .A3(new_n442), .ZN(new_n711));
  INV_X1    g510(.A(new_n702), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n713), .A3(new_n677), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G43gat), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n712), .B2(new_n677), .ZN(new_n716));
  OAI211_X1 g515(.A(KEYINPUT47), .B(new_n711), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n711), .B(KEYINPUT107), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n710), .B1(new_n712), .B2(new_n677), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n717), .B1(KEYINPUT47), .B2(new_n720), .ZN(G1330gat));
  OAI21_X1  g520(.A(G50gat), .B1(new_n702), .B2(new_n272), .ZN(new_n722));
  INV_X1    g521(.A(G50gat), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n686), .A2(new_n723), .A3(new_n680), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT48), .Z(G1331gat));
  NOR2_X1   g525(.A1(new_n657), .A2(new_n630), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n698), .A2(new_n581), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n505), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(new_n477), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n732), .B(new_n733), .Z(G1333gat));
  NAND3_X1  g533(.A1(new_n728), .A2(G71gat), .A3(new_n677), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n728), .A2(new_n442), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(G71gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n728), .A2(new_n680), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT109), .B(G78gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n630), .A2(new_n646), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n581), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n701), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n484), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n698), .A2(new_n655), .A3(new_n742), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n698), .A2(KEYINPUT51), .A3(new_n655), .A4(new_n742), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(KEYINPUT110), .A3(new_n750), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n747), .A2(KEYINPUT110), .A3(new_n748), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n580), .A2(new_n484), .A3(G85gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT111), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n746), .A2(new_n755), .ZN(G1336gat));
  NAND3_X1  g555(.A1(new_n749), .A2(KEYINPUT113), .A3(new_n750), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n580), .A2(new_n476), .A3(G92gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n747), .A2(new_n759), .A3(new_n748), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n757), .A2(KEYINPUT114), .A3(new_n758), .A4(new_n760), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765));
  AOI211_X1 g564(.A(new_n476), .B(new_n743), .C1(new_n690), .C2(new_n700), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(new_n468), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n701), .A2(new_n477), .A3(new_n744), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(KEYINPUT112), .A3(G92gat), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n763), .A2(new_n764), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT52), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n476), .A2(G92gat), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n751), .A2(new_n752), .A3(new_n581), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n768), .A2(G92gat), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n777), .A2(KEYINPUT52), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(KEYINPUT52), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n775), .A2(new_n776), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n770), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n773), .A2(new_n780), .A3(new_n781), .ZN(G1337gat));
  NOR3_X1   g581(.A1(new_n745), .A2(new_n418), .A3(new_n676), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n751), .A2(new_n752), .A3(new_n581), .A4(new_n442), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n418), .B2(new_n784), .ZN(G1338gat));
  NOR2_X1   g584(.A1(new_n272), .A2(G106gat), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n751), .A2(new_n752), .A3(new_n581), .A4(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G106gat), .B1(new_n745), .B2(new_n272), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n757), .A2(new_n581), .A3(new_n760), .A4(new_n786), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n788), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n792), .A2(KEYINPUT117), .A3(KEYINPUT53), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT117), .B1(new_n792), .B2(KEYINPUT53), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n790), .B1(new_n793), .B2(new_n794), .ZN(G1339gat));
  NAND2_X1  g594(.A1(new_n727), .A2(new_n580), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n616), .A2(new_n619), .A3(new_n625), .ZN(new_n798));
  INV_X1    g597(.A(new_n624), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n611), .A2(new_n613), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n617), .A2(new_n618), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(KEYINPUT118), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n566), .A2(new_n567), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n568), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n807), .B(new_n577), .C1(KEYINPUT54), .C2(new_n568), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n810), .A2(new_n579), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n655), .B(new_n812), .C1(new_n803), .C2(new_n813), .ZN(new_n814));
  OR3_X1    g613(.A1(new_n805), .A2(new_n814), .A3(KEYINPUT119), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT119), .B1(new_n805), .B2(new_n814), .ZN(new_n816));
  INV_X1    g615(.A(new_n812), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n628), .B2(new_n629), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n580), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n656), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n646), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n797), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n823), .A2(new_n443), .A3(new_n680), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n505), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(new_n476), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n630), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G113gat), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n285), .A3(new_n630), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1340gat));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n581), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(G120gat), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n826), .A2(new_n287), .A3(new_n581), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1341gat));
  NAND3_X1  g633(.A1(new_n825), .A2(new_n646), .A3(new_n476), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g635(.A1(new_n656), .A2(new_n477), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT120), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n825), .A2(new_n274), .A3(new_n838), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n825), .A2(new_n837), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n840), .B(new_n841), .C1(new_n274), .C2(new_n842), .ZN(G1343gat));
  NOR2_X1   g642(.A1(new_n823), .A2(new_n272), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n628), .A2(new_n629), .B1(new_n812), .B2(KEYINPUT121), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n812), .A2(KEYINPUT121), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n819), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n815), .B(new_n816), .C1(new_n849), .C2(new_n655), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n797), .B1(new_n850), .B2(new_n822), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT57), .B1(new_n851), .B2(new_n272), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n677), .A2(new_n484), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n476), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n846), .A2(new_n852), .A3(new_n630), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G141gat), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n823), .A2(new_n272), .A3(new_n854), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n213), .A3(new_n630), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT58), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n857), .A2(new_n862), .A3(new_n859), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(G1344gat));
  NAND3_X1  g663(.A1(new_n858), .A2(new_n215), .A3(new_n581), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n849), .A2(new_n655), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n805), .A2(new_n814), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n646), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n796), .A2(KEYINPUT122), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n727), .A2(new_n871), .A3(new_n580), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n845), .B(new_n680), .C1(new_n869), .C2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT57), .B1(new_n823), .B2(new_n272), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n874), .A2(new_n875), .A3(new_n581), .A4(new_n855), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n215), .B1(new_n876), .B2(KEYINPUT123), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n878), .A2(new_n879), .A3(new_n581), .A4(new_n855), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n866), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n846), .A2(new_n852), .A3(new_n581), .A4(new_n855), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n882), .A2(new_n866), .A3(G148gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n865), .B1(new_n881), .B2(new_n883), .ZN(G1345gat));
  AOI21_X1  g683(.A(G155gat), .B1(new_n858), .B2(new_n646), .ZN(new_n885));
  AND4_X1   g684(.A1(new_n646), .A2(new_n846), .A3(new_n852), .A4(new_n855), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(G155gat), .ZN(G1346gat));
  NAND4_X1  g686(.A1(new_n846), .A2(new_n852), .A3(new_n655), .A4(new_n855), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n211), .A3(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n211), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n844), .A2(new_n893), .A3(new_n838), .A4(new_n853), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n505), .A2(new_n476), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n824), .A2(new_n896), .ZN(new_n897));
  OR3_X1    g696(.A1(new_n897), .A2(G169gat), .A3(new_n631), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n896), .B(KEYINPUT125), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n824), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n631), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n901), .ZN(G1348gat));
  INV_X1    g701(.A(new_n897), .ZN(new_n903));
  AOI21_X1  g702(.A(G176gat), .B1(new_n903), .B2(new_n581), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n900), .A2(new_n580), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(G176gat), .B2(new_n905), .ZN(G1349gat));
  OAI21_X1  g705(.A(G183gat), .B1(new_n900), .B2(new_n822), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n646), .A2(new_n364), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n897), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT60), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n907), .B(new_n911), .C1(new_n897), .C2(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1350gat));
  NAND3_X1  g712(.A1(new_n903), .A2(new_n655), .A3(new_n363), .ZN(new_n914));
  OAI21_X1  g713(.A(G190gat), .B1(new_n900), .B2(new_n656), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n915), .A2(KEYINPUT61), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(KEYINPUT61), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G1351gat));
  AND3_X1   g717(.A1(new_n844), .A2(new_n676), .A3(new_n896), .ZN(new_n919));
  INV_X1    g718(.A(G197gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n920), .A3(new_n630), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n874), .A2(new_n875), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n874), .A2(new_n875), .A3(KEYINPUT126), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n899), .A2(new_n676), .ZN(new_n926));
  AND4_X1   g725(.A1(new_n630), .A2(new_n924), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n921), .B1(new_n927), .B2(new_n920), .ZN(G1352gat));
  INV_X1    g727(.A(G204gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n919), .A2(new_n929), .A3(new_n581), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n932));
  AND4_X1   g731(.A1(new_n581), .A2(new_n924), .A3(new_n925), .A4(new_n926), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n931), .B(new_n932), .C1(new_n933), .C2(new_n929), .ZN(G1353gat));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n226), .A3(new_n646), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n878), .A2(new_n646), .A3(new_n926), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  NAND3_X1  g738(.A1(new_n919), .A2(new_n227), .A3(new_n655), .ZN(new_n940));
  AND4_X1   g739(.A1(new_n655), .A2(new_n924), .A3(new_n925), .A4(new_n926), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n227), .ZN(G1355gat));
endmodule


