

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n387, n388, n389, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784;

  INV_X1 U372 ( .A(n639), .ZN(n351) );
  AND2_X1 U373 ( .A1(n450), .A2(n391), .ZN(n697) );
  AND2_X1 U374 ( .A1(n415), .A2(n417), .ZN(n365) );
  AND2_X1 U375 ( .A1(n409), .A2(n416), .ZN(n411) );
  AND2_X1 U376 ( .A1(n570), .A2(n569), .ZN(n703) );
  XNOR2_X1 U377 ( .A(n467), .B(n364), .ZN(n406) );
  XNOR2_X1 U378 ( .A(n402), .B(n766), .ZN(n530) );
  XNOR2_X1 U379 ( .A(n400), .B(n551), .ZN(n765) );
  XNOR2_X1 U380 ( .A(n453), .B(G101), .ZN(n552) );
  INV_X1 U381 ( .A(KEYINPUT69), .ZN(n453) );
  NOR2_X1 U382 ( .A1(n776), .A2(n351), .ZN(n360) );
  XNOR2_X2 U383 ( .A(n442), .B(n533), .ZN(n685) );
  NAND2_X1 U384 ( .A1(n566), .A2(n523), .ZN(n384) );
  XNOR2_X1 U385 ( .A(n493), .B(n492), .ZN(n566) );
  XNOR2_X2 U386 ( .A(n442), .B(n362), .ZN(n651) );
  NAND2_X1 U387 ( .A1(n427), .A2(n354), .ZN(n641) );
  NAND2_X1 U388 ( .A1(n357), .A2(n358), .ZN(n427) );
  XNOR2_X2 U389 ( .A(n420), .B(KEYINPUT83), .ZN(n658) );
  NAND2_X2 U390 ( .A1(n630), .A2(n629), .ZN(n420) );
  XNOR2_X2 U391 ( .A(n352), .B(n369), .ZN(n776) );
  NAND2_X1 U392 ( .A1(n575), .A2(n421), .ZN(n352) );
  INV_X1 U393 ( .A(KEYINPUT89), .ZN(n394) );
  XNOR2_X2 U394 ( .A(n361), .B(n640), .ZN(n676) );
  INV_X2 U395 ( .A(G122), .ZN(n472) );
  NOR2_X2 U396 ( .A1(n567), .A2(n746), .ZN(n395) );
  NAND2_X2 U397 ( .A1(n413), .A2(n412), .ZN(n564) );
  XNOR2_X2 U398 ( .A(n553), .B(n368), .ZN(n601) );
  NOR2_X2 U399 ( .A1(n784), .A2(n657), .ZN(n424) );
  XNOR2_X2 U400 ( .A(n586), .B(n585), .ZN(n784) );
  XNOR2_X2 U401 ( .A(n589), .B(KEYINPUT106), .ZN(n608) );
  XNOR2_X1 U402 ( .A(n371), .B(n465), .ZN(n464) );
  OR2_X1 U403 ( .A1(n622), .A2(n385), .ZN(n604) );
  NOR2_X1 U404 ( .A1(n583), .A2(n483), .ZN(n484) );
  XNOR2_X1 U405 ( .A(n530), .B(n765), .ZN(n377) );
  XNOR2_X1 U406 ( .A(n399), .B(G119), .ZN(n551) );
  INV_X1 U407 ( .A(KEYINPUT80), .ZN(n392) );
  INV_X1 U408 ( .A(G131), .ZN(n463) );
  NAND2_X1 U409 ( .A1(n419), .A2(KEYINPUT2), .ZN(n631) );
  AND2_X1 U410 ( .A1(n571), .A2(n609), .ZN(n375) );
  AND2_X1 U411 ( .A1(n444), .A2(n703), .ZN(n443) );
  NAND2_X1 U412 ( .A1(n437), .A2(n436), .ZN(n722) );
  NAND2_X1 U413 ( .A1(n448), .A2(n584), .ZN(n444) );
  NOR2_X1 U414 ( .A1(n726), .A2(n728), .ZN(n593) );
  NOR2_X1 U415 ( .A1(n607), .A2(n491), .ZN(n493) );
  XNOR2_X1 U416 ( .A(n588), .B(n470), .ZN(n735) );
  XNOR2_X1 U417 ( .A(n506), .B(n505), .ZN(n570) );
  AND2_X1 U418 ( .A1(n406), .A2(n598), .ZN(n382) );
  NAND2_X1 U419 ( .A1(n433), .A2(n429), .ZN(n383) );
  AND2_X1 U420 ( .A1(n435), .A2(n434), .ZN(n433) );
  NOR2_X1 U421 ( .A1(n651), .A2(G902), .ZN(n467) );
  XNOR2_X1 U422 ( .A(n377), .B(n477), .ZN(n644) );
  XNOR2_X1 U423 ( .A(n405), .B(n403), .ZN(n477) );
  XNOR2_X1 U424 ( .A(n511), .B(n510), .ZN(n536) );
  XNOR2_X1 U425 ( .A(n539), .B(n454), .ZN(n540) );
  XNOR2_X1 U426 ( .A(n463), .B(KEYINPUT70), .ZN(n531) );
  XNOR2_X1 U427 ( .A(n394), .B(G110), .ZN(n401) );
  XNOR2_X1 U428 ( .A(G113), .B(G143), .ZN(n499) );
  INV_X1 U429 ( .A(KEYINPUT16), .ZN(n473) );
  XNOR2_X1 U430 ( .A(G137), .B(KEYINPUT4), .ZN(n449) );
  XNOR2_X1 U431 ( .A(G104), .B(G107), .ZN(n471) );
  INV_X1 U432 ( .A(KEYINPUT64), .ZN(n474) );
  INV_X1 U433 ( .A(KEYINPUT118), .ZN(n353) );
  XNOR2_X1 U434 ( .A(n353), .B(n764), .ZN(G75) );
  XNOR2_X1 U435 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U436 ( .A(n512), .B(n473), .ZN(n400) );
  XNOR2_X1 U437 ( .A(n484), .B(KEYINPUT19), .ZN(n607) );
  XNOR2_X1 U438 ( .A(n393), .B(n392), .ZN(n354) );
  XNOR2_X1 U439 ( .A(n393), .B(n392), .ZN(n720) );
  BUF_X1 U440 ( .A(n722), .Z(n355) );
  BUF_X1 U441 ( .A(n776), .Z(n356) );
  NAND2_X1 U442 ( .A1(n387), .A2(n360), .ZN(n357) );
  OR2_X1 U443 ( .A1(n359), .A2(n637), .ZN(n358) );
  INV_X1 U444 ( .A(n639), .ZN(n359) );
  NAND2_X1 U445 ( .A1(n427), .A2(n720), .ZN(n361) );
  NAND2_X1 U446 ( .A1(n433), .A2(n429), .ZN(n588) );
  NOR2_X1 U447 ( .A1(n587), .A2(n737), .ZN(n597) );
  XNOR2_X1 U448 ( .A(n426), .B(n425), .ZN(n582) );
  INV_X1 U449 ( .A(KEYINPUT30), .ZN(n425) );
  NOR2_X1 U450 ( .A1(G902), .A2(G237), .ZN(n478) );
  NAND2_X1 U451 ( .A1(G469), .A2(G902), .ZN(n434) );
  NAND2_X1 U452 ( .A1(n432), .A2(n431), .ZN(n430) );
  INV_X1 U453 ( .A(G469), .ZN(n432) );
  INV_X1 U454 ( .A(G902), .ZN(n431) );
  XNOR2_X1 U455 ( .A(n550), .B(KEYINPUT78), .ZN(n469) );
  XNOR2_X1 U456 ( .A(n459), .B(n531), .ZN(n458) );
  XNOR2_X1 U457 ( .A(n449), .B(KEYINPUT72), .ZN(n459) );
  NOR2_X1 U458 ( .A1(n690), .A2(n375), .ZN(n374) );
  XNOR2_X1 U459 ( .A(KEYINPUT15), .B(G902), .ZN(n638) );
  XNOR2_X1 U460 ( .A(G113), .B(KEYINPUT3), .ZN(n399) );
  XNOR2_X1 U461 ( .A(G146), .B(G125), .ZN(n496) );
  XNOR2_X1 U462 ( .A(KEYINPUT88), .B(KEYINPUT0), .ZN(n492) );
  XNOR2_X1 U463 ( .A(n545), .B(n544), .ZN(n546) );
  INV_X1 U464 ( .A(KEYINPUT25), .ZN(n544) );
  AND2_X1 U465 ( .A1(n398), .A2(n447), .ZN(n445) );
  NAND2_X1 U466 ( .A1(n396), .A2(n741), .ZN(n746) );
  NAND2_X1 U467 ( .A1(n381), .A2(n582), .ZN(n448) );
  INV_X1 U468 ( .A(KEYINPUT102), .ZN(n451) );
  BUF_X1 U469 ( .A(n738), .Z(n389) );
  XNOR2_X1 U470 ( .A(KEYINPUT85), .B(KEYINPUT48), .ZN(n620) );
  XOR2_X1 U471 ( .A(G122), .B(G104), .Z(n500) );
  NAND2_X1 U472 ( .A1(G234), .A2(G237), .ZN(n485) );
  NOR2_X1 U473 ( .A1(G953), .A2(G237), .ZN(n548) );
  XNOR2_X1 U474 ( .A(G140), .B(KEYINPUT97), .ZN(n494) );
  XOR2_X1 U475 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n495) );
  INV_X1 U476 ( .A(KEYINPUT79), .ZN(n388) );
  XNOR2_X1 U477 ( .A(G140), .B(KEYINPUT71), .ZN(n534) );
  INV_X1 U478 ( .A(n601), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n457), .B(KEYINPUT103), .ZN(n439) );
  OR2_X2 U480 ( .A1(n644), .A2(n633), .ZN(n481) );
  XNOR2_X1 U481 ( .A(n551), .B(n469), .ZN(n468) );
  XNOR2_X1 U482 ( .A(n538), .B(n455), .ZN(n454) );
  XNOR2_X1 U483 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n455) );
  INV_X1 U484 ( .A(G134), .ZN(n508) );
  INV_X1 U485 ( .A(KEYINPUT8), .ZN(n510) );
  XNOR2_X1 U486 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n475) );
  XNOR2_X1 U487 ( .A(n552), .B(KEYINPUT73), .ZN(n402) );
  XNOR2_X1 U488 ( .A(n404), .B(n496), .ZN(n403) );
  INV_X1 U489 ( .A(KEYINPUT28), .ZN(n456) );
  INV_X1 U490 ( .A(KEYINPUT94), .ZN(n465) );
  NAND2_X1 U491 ( .A1(n383), .A2(n734), .ZN(n371) );
  INV_X1 U492 ( .A(G953), .ZN(n760) );
  XNOR2_X1 U493 ( .A(n395), .B(n568), .ZN(n710) );
  INV_X1 U494 ( .A(n448), .ZN(n466) );
  NOR2_X1 U495 ( .A1(n741), .A2(n587), .ZN(n391) );
  AND2_X1 U496 ( .A1(n574), .A2(n376), .ZN(n690) );
  NOR2_X1 U497 ( .A1(n422), .A2(n389), .ZN(n376) );
  XNOR2_X1 U498 ( .A(n378), .B(n370), .ZN(n689) );
  XOR2_X1 U499 ( .A(n468), .B(n366), .Z(n362) );
  XOR2_X1 U500 ( .A(n495), .B(n494), .Z(n363) );
  XNOR2_X1 U501 ( .A(G472), .B(KEYINPUT75), .ZN(n364) );
  XOR2_X1 U502 ( .A(n552), .B(n549), .Z(n366) );
  XOR2_X1 U503 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n367) );
  XOR2_X1 U504 ( .A(KEYINPUT6), .B(KEYINPUT100), .Z(n368) );
  XOR2_X1 U505 ( .A(KEYINPUT84), .B(KEYINPUT45), .Z(n369) );
  XOR2_X1 U506 ( .A(n687), .B(n686), .Z(n370) );
  NOR2_X2 U507 ( .A1(n738), .A2(n737), .ZN(n734) );
  XNOR2_X1 U508 ( .A(n372), .B(KEYINPUT87), .ZN(n421) );
  NAND2_X1 U509 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U510 ( .A1(n564), .A2(KEYINPUT44), .ZN(n373) );
  NAND2_X1 U511 ( .A1(n684), .A2(G469), .ZN(n378) );
  XNOR2_X2 U512 ( .A(n641), .B(n640), .ZN(n684) );
  XNOR2_X1 U513 ( .A(n651), .B(KEYINPUT62), .ZN(n652) );
  INV_X1 U514 ( .A(n567), .ZN(n379) );
  XNOR2_X2 U515 ( .A(n384), .B(n525), .ZN(n554) );
  BUF_X1 U516 ( .A(n660), .Z(n380) );
  AND2_X1 U517 ( .A1(n464), .A2(n598), .ZN(n381) );
  NOR2_X2 U518 ( .A1(n669), .A2(G902), .ZN(n547) );
  INV_X1 U519 ( .A(n566), .ZN(n567) );
  XNOR2_X1 U520 ( .A(n428), .B(n498), .ZN(n677) );
  BUF_X1 U521 ( .A(n607), .Z(n423) );
  XNOR2_X1 U522 ( .A(n503), .B(n363), .ZN(n428) );
  XNOR2_X1 U523 ( .A(n583), .B(KEYINPUT38), .ZN(n724) );
  BUF_X1 U524 ( .A(n583), .Z(n385) );
  BUF_X1 U525 ( .A(n658), .Z(n717) );
  XNOR2_X2 U526 ( .A(n401), .B(n471), .ZN(n766) );
  NOR2_X2 U527 ( .A1(n783), .A2(n697), .ZN(n561) );
  NAND2_X1 U528 ( .A1(n443), .A2(n445), .ZN(n586) );
  XNOR2_X1 U529 ( .A(n658), .B(n388), .ZN(n387) );
  NAND2_X1 U530 ( .A1(n735), .A2(n734), .ZN(n457) );
  NOR2_X2 U531 ( .A1(n776), .A2(n631), .ZN(n393) );
  NAND2_X1 U532 ( .A1(n567), .A2(KEYINPUT34), .ZN(n462) );
  XNOR2_X1 U533 ( .A(n408), .B(n456), .ZN(n407) );
  NAND2_X1 U534 ( .A1(n554), .A2(n601), .ZN(n573) );
  INV_X1 U535 ( .A(n457), .ZN(n396) );
  NAND2_X1 U536 ( .A1(n397), .A2(n381), .ZN(n398) );
  AND2_X1 U537 ( .A1(n446), .A2(n582), .ZN(n397) );
  XNOR2_X2 U538 ( .A(n472), .B(G116), .ZN(n512) );
  NAND2_X1 U539 ( .A1(n526), .A2(G224), .ZN(n404) );
  XNOR2_X1 U540 ( .A(n509), .B(n476), .ZN(n405) );
  INV_X1 U541 ( .A(n406), .ZN(n553) );
  NAND2_X1 U542 ( .A1(n406), .A2(n723), .ZN(n426) );
  NAND2_X1 U543 ( .A1(n407), .A2(n383), .ZN(n589) );
  NAND2_X1 U544 ( .A1(n382), .A2(n597), .ZN(n408) );
  NAND2_X1 U545 ( .A1(n722), .A2(KEYINPUT34), .ZN(n416) );
  INV_X1 U546 ( .A(n461), .ZN(n409) );
  NAND2_X1 U547 ( .A1(n440), .A2(n410), .ZN(n417) );
  INV_X1 U548 ( .A(n722), .ZN(n410) );
  NOR2_X1 U549 ( .A1(n461), .A2(KEYINPUT35), .ZN(n415) );
  NAND2_X1 U550 ( .A1(n411), .A2(n417), .ZN(n414) );
  NAND2_X1 U551 ( .A1(n365), .A2(n416), .ZN(n412) );
  NAND2_X1 U552 ( .A1(n414), .A2(KEYINPUT35), .ZN(n413) );
  NAND2_X1 U553 ( .A1(n439), .A2(n418), .ZN(n438) );
  INV_X1 U554 ( .A(n420), .ZN(n419) );
  NAND2_X1 U555 ( .A1(n462), .A2(n612), .ZN(n461) );
  BUF_X1 U556 ( .A(n735), .Z(n422) );
  XNOR2_X1 U557 ( .A(n452), .B(n451), .ZN(n450) );
  XNOR2_X1 U558 ( .A(n424), .B(KEYINPUT46), .ZN(n619) );
  NOR2_X2 U559 ( .A1(n606), .A2(n605), .ZN(n713) );
  NAND2_X1 U560 ( .A1(n685), .A2(G469), .ZN(n435) );
  OR2_X1 U561 ( .A1(n685), .A2(n430), .ZN(n429) );
  NAND2_X1 U562 ( .A1(n441), .A2(n439), .ZN(n436) );
  NAND2_X1 U563 ( .A1(n438), .A2(n367), .ZN(n437) );
  NOR2_X1 U564 ( .A1(n567), .A2(KEYINPUT34), .ZN(n440) );
  NOR2_X1 U565 ( .A1(n601), .A2(n367), .ZN(n441) );
  XNOR2_X2 U566 ( .A(n660), .B(G146), .ZN(n442) );
  NAND2_X1 U567 ( .A1(n445), .A2(n444), .ZN(n627) );
  AND2_X1 U568 ( .A1(n724), .A2(KEYINPUT39), .ZN(n446) );
  OR2_X1 U569 ( .A1(n724), .A2(KEYINPUT39), .ZN(n447) );
  NAND2_X1 U570 ( .A1(n554), .A2(n605), .ZN(n452) );
  XNOR2_X2 U571 ( .A(n532), .B(n458), .ZN(n660) );
  XNOR2_X2 U572 ( .A(n509), .B(n508), .ZN(n532) );
  XNOR2_X2 U573 ( .A(n460), .B(G143), .ZN(n509) );
  XNOR2_X2 U574 ( .A(G128), .B(KEYINPUT65), .ZN(n460) );
  AND2_X1 U575 ( .A1(n464), .A2(n553), .ZN(n565) );
  NAND2_X1 U576 ( .A1(n466), .A2(n613), .ZN(n614) );
  NOR2_X2 U577 ( .A1(n608), .A2(n423), .ZN(n704) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(KEYINPUT67), .Z(n470) );
  INV_X1 U579 ( .A(KEYINPUT44), .ZN(n559) );
  INV_X1 U580 ( .A(KEYINPUT22), .ZN(n524) );
  XNOR2_X1 U581 ( .A(n524), .B(KEYINPUT76), .ZN(n525) );
  INV_X1 U582 ( .A(n422), .ZN(n605) );
  NOR2_X1 U583 ( .A1(n573), .A2(n556), .ZN(n558) );
  INV_X1 U584 ( .A(n553), .ZN(n741) );
  INV_X1 U585 ( .A(KEYINPUT63), .ZN(n655) );
  XNOR2_X2 U586 ( .A(n474), .B(G953), .ZN(n526) );
  XNOR2_X1 U587 ( .A(n475), .B(KEYINPUT4), .ZN(n476) );
  INV_X1 U588 ( .A(n638), .ZN(n633) );
  XNOR2_X1 U589 ( .A(n478), .B(KEYINPUT77), .ZN(n482) );
  NAND2_X1 U590 ( .A1(n482), .A2(G210), .ZN(n479) );
  XNOR2_X1 U591 ( .A(n479), .B(KEYINPUT90), .ZN(n480) );
  XNOR2_X2 U592 ( .A(n481), .B(n480), .ZN(n583) );
  NAND2_X1 U593 ( .A1(n482), .A2(G214), .ZN(n723) );
  INV_X1 U594 ( .A(n723), .ZN(n483) );
  XNOR2_X1 U595 ( .A(KEYINPUT91), .B(G898), .ZN(n774) );
  NAND2_X1 U596 ( .A1(G953), .A2(n774), .ZN(n770) );
  XNOR2_X1 U597 ( .A(n485), .B(KEYINPUT14), .ZN(n488) );
  NAND2_X1 U598 ( .A1(G902), .A2(n488), .ZN(n486) );
  NOR2_X1 U599 ( .A1(n770), .A2(n486), .ZN(n487) );
  XNOR2_X1 U600 ( .A(n487), .B(KEYINPUT92), .ZN(n490) );
  NAND2_X1 U601 ( .A1(G952), .A2(n760), .ZN(n576) );
  INV_X1 U602 ( .A(n488), .ZN(n753) );
  NOR2_X1 U603 ( .A1(n576), .A2(n753), .ZN(n489) );
  NOR2_X1 U604 ( .A1(n490), .A2(n489), .ZN(n491) );
  NAND2_X1 U605 ( .A1(G214), .A2(n548), .ZN(n497) );
  XNOR2_X1 U606 ( .A(KEYINPUT10), .B(n496), .ZN(n535) );
  XNOR2_X1 U607 ( .A(n497), .B(n535), .ZN(n498) );
  XNOR2_X1 U608 ( .A(n531), .B(KEYINPUT96), .ZN(n502) );
  XNOR2_X1 U609 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U610 ( .A(n502), .B(n501), .ZN(n503) );
  NOR2_X1 U611 ( .A1(G902), .A2(n677), .ZN(n504) );
  XOR2_X1 U612 ( .A(G475), .B(n504), .Z(n506) );
  INV_X1 U613 ( .A(KEYINPUT13), .ZN(n505) );
  INV_X1 U614 ( .A(n570), .ZN(n520) );
  XOR2_X1 U615 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n507) );
  XNOR2_X1 U616 ( .A(G478), .B(n507), .ZN(n519) );
  NAND2_X1 U617 ( .A1(n526), .A2(G234), .ZN(n511) );
  NAND2_X1 U618 ( .A1(n536), .A2(G217), .ZN(n516) );
  XOR2_X1 U619 ( .A(KEYINPUT7), .B(n512), .Z(n514) );
  XNOR2_X1 U620 ( .A(G107), .B(KEYINPUT9), .ZN(n513) );
  XNOR2_X1 U621 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U622 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U623 ( .A(n532), .B(n517), .ZN(n673) );
  NOR2_X1 U624 ( .A1(G902), .A2(n673), .ZN(n518) );
  XNOR2_X1 U625 ( .A(n519), .B(n518), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n520), .A2(n569), .ZN(n726) );
  NAND2_X1 U627 ( .A1(n638), .A2(G234), .ZN(n521) );
  XNOR2_X1 U628 ( .A(n521), .B(KEYINPUT20), .ZN(n543) );
  NAND2_X1 U629 ( .A1(G221), .A2(n543), .ZN(n522) );
  XNOR2_X1 U630 ( .A(KEYINPUT21), .B(n522), .ZN(n737) );
  NOR2_X1 U631 ( .A1(n726), .A2(n737), .ZN(n523) );
  INV_X1 U632 ( .A(n534), .ZN(n528) );
  NAND2_X1 U633 ( .A1(n526), .A2(G227), .ZN(n527) );
  XOR2_X1 U634 ( .A(n528), .B(n527), .Z(n529) );
  XNOR2_X1 U635 ( .A(n530), .B(n529), .ZN(n533) );
  XNOR2_X1 U636 ( .A(n535), .B(n534), .ZN(n659) );
  NAND2_X1 U637 ( .A1(n536), .A2(G221), .ZN(n541) );
  XNOR2_X1 U638 ( .A(G128), .B(G110), .ZN(n537) );
  XNOR2_X1 U639 ( .A(n537), .B(KEYINPUT23), .ZN(n539) );
  XNOR2_X1 U640 ( .A(G119), .B(G137), .ZN(n538) );
  XNOR2_X1 U641 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U642 ( .A(n542), .B(n659), .ZN(n669) );
  NAND2_X1 U643 ( .A1(n543), .A2(G217), .ZN(n545) );
  XNOR2_X2 U644 ( .A(n547), .B(n546), .ZN(n738) );
  NAND2_X1 U645 ( .A1(n548), .A2(G210), .ZN(n550) );
  XOR2_X1 U646 ( .A(G116), .B(KEYINPUT5), .Z(n549) );
  INV_X1 U647 ( .A(n738), .ZN(n587) );
  NOR2_X1 U648 ( .A1(n605), .A2(n587), .ZN(n555) );
  XNOR2_X1 U649 ( .A(n555), .B(KEYINPUT101), .ZN(n556) );
  XOR2_X1 U650 ( .A(KEYINPUT81), .B(KEYINPUT32), .Z(n557) );
  XNOR2_X1 U651 ( .A(n558), .B(n557), .ZN(n783) );
  XNOR2_X1 U652 ( .A(n561), .B(n559), .ZN(n563) );
  INV_X1 U653 ( .A(n569), .ZN(n560) );
  AND2_X1 U654 ( .A1(n570), .A2(n560), .ZN(n612) );
  NAND2_X1 U655 ( .A1(n561), .A2(n564), .ZN(n562) );
  NAND2_X1 U656 ( .A1(n563), .A2(n562), .ZN(n575) );
  NAND2_X1 U657 ( .A1(n379), .A2(n565), .ZN(n694) );
  XOR2_X1 U658 ( .A(KEYINPUT95), .B(KEYINPUT31), .Z(n568) );
  NAND2_X1 U659 ( .A1(n694), .A2(n710), .ZN(n571) );
  NOR2_X1 U660 ( .A1(n570), .A2(n569), .ZN(n700) );
  NOR2_X1 U661 ( .A1(n700), .A2(n703), .ZN(n729) );
  INV_X1 U662 ( .A(n729), .ZN(n609) );
  INV_X1 U663 ( .A(KEYINPUT86), .ZN(n572) );
  XNOR2_X1 U664 ( .A(n573), .B(n572), .ZN(n574) );
  INV_X1 U665 ( .A(n576), .ZN(n580) );
  INV_X1 U666 ( .A(G900), .ZN(n577) );
  NAND2_X1 U667 ( .A1(n577), .A2(G902), .ZN(n578) );
  NOR2_X1 U668 ( .A1(n526), .A2(n578), .ZN(n579) );
  NOR2_X1 U669 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U670 ( .A1(n581), .A2(n753), .ZN(n598) );
  INV_X1 U671 ( .A(KEYINPUT39), .ZN(n584) );
  INV_X1 U672 ( .A(KEYINPUT40), .ZN(n585) );
  NAND2_X1 U673 ( .A1(n724), .A2(n723), .ZN(n728) );
  XNOR2_X1 U674 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n591) );
  INV_X1 U675 ( .A(KEYINPUT107), .ZN(n590) );
  XNOR2_X1 U676 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U677 ( .A(n593), .B(n592), .ZN(n757) );
  NOR2_X1 U678 ( .A1(n608), .A2(n757), .ZN(n596) );
  INV_X1 U679 ( .A(KEYINPUT109), .ZN(n594) );
  XNOR2_X1 U680 ( .A(n594), .B(KEYINPUT42), .ZN(n595) );
  XNOR2_X1 U681 ( .A(n596), .B(n595), .ZN(n657) );
  INV_X1 U682 ( .A(n597), .ZN(n600) );
  NAND2_X1 U683 ( .A1(n598), .A2(n723), .ZN(n599) );
  NOR2_X1 U684 ( .A1(n600), .A2(n599), .ZN(n603) );
  INV_X1 U685 ( .A(n703), .ZN(n706) );
  NOR2_X1 U686 ( .A1(n601), .A2(n706), .ZN(n602) );
  NAND2_X1 U687 ( .A1(n603), .A2(n602), .ZN(n622) );
  XNOR2_X1 U688 ( .A(n604), .B(KEYINPUT36), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n609), .A2(n704), .ZN(n611) );
  INV_X1 U690 ( .A(KEYINPUT47), .ZN(n610) );
  XNOR2_X1 U691 ( .A(n611), .B(n610), .ZN(n616) );
  INV_X1 U692 ( .A(n385), .ZN(n624) );
  AND2_X1 U693 ( .A1(n612), .A2(n624), .ZN(n613) );
  XNOR2_X1 U694 ( .A(n614), .B(KEYINPUT105), .ZN(n781) );
  INV_X1 U695 ( .A(n781), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n713), .A2(n617), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n621), .B(n620), .ZN(n630) );
  NOR2_X1 U700 ( .A1(n422), .A2(n622), .ZN(n623) );
  XNOR2_X1 U701 ( .A(n623), .B(KEYINPUT43), .ZN(n625) );
  NOR2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U703 ( .A(n626), .B(KEYINPUT104), .ZN(n782) );
  INV_X1 U704 ( .A(n700), .ZN(n709) );
  OR2_X1 U705 ( .A1(n627), .A2(n709), .ZN(n715) );
  INV_X1 U706 ( .A(n715), .ZN(n628) );
  NOR2_X1 U707 ( .A1(n782), .A2(n628), .ZN(n629) );
  INV_X1 U708 ( .A(KEYINPUT2), .ZN(n634) );
  NOR2_X1 U709 ( .A1(n634), .A2(KEYINPUT68), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n634), .A2(KEYINPUT68), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(KEYINPUT68), .ZN(n639) );
  INV_X1 U714 ( .A(KEYINPUT66), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n676), .A2(G210), .ZN(n646) );
  XNOR2_X1 U716 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n642) );
  XOR2_X1 U717 ( .A(n642), .B(KEYINPUT120), .Z(n643) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(n649) );
  INV_X1 U719 ( .A(n526), .ZN(n648) );
  INV_X1 U720 ( .A(G952), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n648), .A2(n647), .ZN(n680) );
  INV_X1 U722 ( .A(n680), .ZN(n688) );
  NOR2_X2 U723 ( .A1(n649), .A2(n688), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n650), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U725 ( .A1(n676), .A2(G472), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X2 U727 ( .A1(n654), .A2(n688), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n656), .B(n655), .ZN(G57) );
  XOR2_X1 U729 ( .A(n657), .B(G137), .Z(G39) );
  XNOR2_X1 U730 ( .A(n380), .B(n659), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n717), .B(n662), .ZN(n661) );
  NAND2_X1 U732 ( .A1(n661), .A2(n526), .ZN(n668) );
  XOR2_X1 U733 ( .A(n662), .B(G227), .Z(n663) );
  XNOR2_X1 U734 ( .A(n663), .B(KEYINPUT126), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n664), .A2(G900), .ZN(n665) );
  NAND2_X1 U736 ( .A1(G953), .A2(n665), .ZN(n666) );
  XOR2_X1 U737 ( .A(KEYINPUT127), .B(n666), .Z(n667) );
  NAND2_X1 U738 ( .A1(n668), .A2(n667), .ZN(G72) );
  NAND2_X1 U739 ( .A1(n684), .A2(G217), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n669), .B(KEYINPUT122), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U742 ( .A1(n672), .A2(n688), .ZN(G66) );
  NAND2_X1 U743 ( .A1(n684), .A2(G478), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U745 ( .A1(n675), .A2(n688), .ZN(G63) );
  NAND2_X1 U746 ( .A1(n684), .A2(G475), .ZN(n679) );
  XNOR2_X1 U747 ( .A(n677), .B(KEYINPUT59), .ZN(n678) );
  XNOR2_X1 U748 ( .A(n679), .B(n678), .ZN(n681) );
  NAND2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n683) );
  INV_X1 U750 ( .A(KEYINPUT60), .ZN(n682) );
  XNOR2_X1 U751 ( .A(n683), .B(n682), .ZN(G60) );
  XOR2_X1 U752 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n687) );
  XNOR2_X1 U753 ( .A(n685), .B(KEYINPUT121), .ZN(n686) );
  NOR2_X1 U754 ( .A1(n689), .A2(n688), .ZN(G54) );
  XOR2_X1 U755 ( .A(n690), .B(G101), .Z(G3) );
  NOR2_X1 U756 ( .A1(n706), .A2(n694), .ZN(n691) );
  XOR2_X1 U757 ( .A(G104), .B(n691), .Z(G6) );
  XOR2_X1 U758 ( .A(KEYINPUT110), .B(KEYINPUT26), .Z(n693) );
  XNOR2_X1 U759 ( .A(G107), .B(KEYINPUT27), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n693), .B(n692), .ZN(n696) );
  NOR2_X1 U761 ( .A1(n709), .A2(n694), .ZN(n695) );
  XOR2_X1 U762 ( .A(n696), .B(n695), .Z(G9) );
  XOR2_X1 U763 ( .A(n697), .B(G110), .Z(G12) );
  XOR2_X1 U764 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n699) );
  XNOR2_X1 U765 ( .A(G128), .B(KEYINPUT29), .ZN(n698) );
  XNOR2_X1 U766 ( .A(n699), .B(n698), .ZN(n702) );
  NAND2_X1 U767 ( .A1(n704), .A2(n700), .ZN(n701) );
  XOR2_X1 U768 ( .A(n702), .B(n701), .Z(G30) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U770 ( .A(n705), .B(G146), .ZN(G48) );
  NOR2_X1 U771 ( .A1(n706), .A2(n710), .ZN(n708) );
  XNOR2_X1 U772 ( .A(G113), .B(KEYINPUT113), .ZN(n707) );
  XNOR2_X1 U773 ( .A(n708), .B(n707), .ZN(G15) );
  NOR2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U775 ( .A(KEYINPUT114), .B(n711), .Z(n712) );
  XNOR2_X1 U776 ( .A(G116), .B(n712), .ZN(G18) );
  XNOR2_X1 U777 ( .A(G125), .B(n713), .ZN(n714) );
  XNOR2_X1 U778 ( .A(n714), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U779 ( .A(G134), .B(n715), .ZN(G36) );
  XOR2_X1 U780 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n763) );
  NAND2_X1 U781 ( .A1(n776), .A2(n634), .ZN(n716) );
  XOR2_X1 U782 ( .A(KEYINPUT82), .B(n716), .Z(n719) );
  NOR2_X1 U783 ( .A1(n717), .A2(KEYINPUT2), .ZN(n718) );
  NOR2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n721) );
  NAND2_X1 U785 ( .A1(n721), .A2(n720), .ZN(n756) );
  NOR2_X1 U786 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U787 ( .A(n725), .B(KEYINPUT116), .ZN(n727) );
  NOR2_X1 U788 ( .A1(n727), .A2(n726), .ZN(n731) );
  NOR2_X1 U789 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U790 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U791 ( .A(KEYINPUT117), .B(n732), .Z(n733) );
  NOR2_X1 U792 ( .A1(n355), .A2(n733), .ZN(n750) );
  OR2_X1 U793 ( .A1(n422), .A2(n734), .ZN(n736) );
  XNOR2_X1 U794 ( .A(KEYINPUT50), .B(n736), .ZN(n744) );
  XOR2_X1 U795 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n740) );
  NAND2_X1 U796 ( .A1(n389), .A2(n737), .ZN(n739) );
  XNOR2_X1 U797 ( .A(n740), .B(n739), .ZN(n742) );
  NOR2_X1 U798 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U799 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U800 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U801 ( .A(KEYINPUT51), .B(n747), .ZN(n748) );
  NOR2_X1 U802 ( .A1(n748), .A2(n757), .ZN(n749) );
  NOR2_X1 U803 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U804 ( .A(n751), .B(KEYINPUT52), .ZN(n752) );
  NOR2_X1 U805 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U806 ( .A1(n754), .A2(G952), .ZN(n755) );
  NAND2_X1 U807 ( .A1(n756), .A2(n755), .ZN(n759) );
  NOR2_X1 U808 ( .A1(n355), .A2(n757), .ZN(n758) );
  NOR2_X1 U809 ( .A1(n759), .A2(n758), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U811 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U812 ( .A(n765), .B(KEYINPUT125), .ZN(n768) );
  XNOR2_X1 U813 ( .A(G101), .B(n766), .ZN(n767) );
  XNOR2_X1 U814 ( .A(n768), .B(n767), .ZN(n769) );
  NAND2_X1 U815 ( .A1(n770), .A2(n769), .ZN(n780) );
  NAND2_X1 U816 ( .A1(G224), .A2(G953), .ZN(n771) );
  XNOR2_X1 U817 ( .A(n771), .B(KEYINPUT123), .ZN(n772) );
  XNOR2_X1 U818 ( .A(n772), .B(KEYINPUT61), .ZN(n773) );
  NOR2_X1 U819 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U820 ( .A(n775), .B(KEYINPUT124), .ZN(n778) );
  NOR2_X1 U821 ( .A1(G953), .A2(n356), .ZN(n777) );
  NOR2_X1 U822 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U823 ( .A(n780), .B(n779), .ZN(G69) );
  XOR2_X1 U824 ( .A(G143), .B(n781), .Z(G45) );
  XOR2_X1 U825 ( .A(n564), .B(G122), .Z(G24) );
  XOR2_X1 U826 ( .A(G140), .B(n782), .Z(G42) );
  XOR2_X1 U827 ( .A(n783), .B(G119), .Z(G21) );
  XOR2_X1 U828 ( .A(n784), .B(G131), .Z(G33) );
endmodule

